module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  input  [31:0] I_2,
  input  [31:0] I_3,
  output [31:0] O_0,
  output [31:0] O_1,
  output [31:0] O_2,
  output [31:0] O_3
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x342_TREADY(dontcare), // @[:@1298.4]
    .io_in_x342_TDATA({I_0,I_1}), // @[:@1298.4]
    .io_in_x342_TID(8'h0),
    .io_in_x342_TDEST(8'h0),
    .io_in_x343_TVALID(valid_down), // @[:@1298.4]
    .io_in_x343_TDATA({O_0,O_1}), // @[:@1298.4]
    .io_in_x343_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x350_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(reset), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh57); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh57); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x344_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x740_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x671_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x345_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x346_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh4); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh4); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x350_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x372_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x720_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x356_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x372_inr_Foreach_kernelx372_inr_Foreach_concrete1( // @[:@5178.2]
  input         clock, // @[:@5179.4]
  input         reset, // @[:@5180.4]
  output        io_in_x346_fifoinpacked_0_wPort_0_en_0, // @[:@5181.4]
  input         io_in_x346_fifoinpacked_0_full, // @[:@5181.4]
  output        io_in_x346_fifoinpacked_0_active_0_in, // @[:@5181.4]
  input         io_in_x346_fifoinpacked_0_active_0_out, // @[:@5181.4]
  input         io_sigsIn_backpressure, // @[:@5181.4]
  input         io_sigsIn_datapathEn, // @[:@5181.4]
  input         io_sigsIn_break, // @[:@5181.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@5181.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@5181.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@5181.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@5181.4]
  input         io_rr // @[:@5181.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@5215.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@5215.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@5227.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@5227.4]
  wire  x720_sub_1_clock; // @[Math.scala 191:24:@5254.4]
  wire  x720_sub_1_reset; // @[Math.scala 191:24:@5254.4]
  wire [31:0] x720_sub_1_io_a; // @[Math.scala 191:24:@5254.4]
  wire [31:0] x720_sub_1_io_b; // @[Math.scala 191:24:@5254.4]
  wire  x720_sub_1_io_flow; // @[Math.scala 191:24:@5254.4]
  wire [31:0] x720_sub_1_io_result; // @[Math.scala 191:24:@5254.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5264.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5264.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5264.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5264.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5264.4]
  wire  x356_sum_1_clock; // @[Math.scala 150:24:@5273.4]
  wire  x356_sum_1_reset; // @[Math.scala 150:24:@5273.4]
  wire [31:0] x356_sum_1_io_a; // @[Math.scala 150:24:@5273.4]
  wire [31:0] x356_sum_1_io_b; // @[Math.scala 150:24:@5273.4]
  wire  x356_sum_1_io_flow; // @[Math.scala 150:24:@5273.4]
  wire [31:0] x356_sum_1_io_result; // @[Math.scala 150:24:@5273.4]
  wire  x357_sum_1_clock; // @[Math.scala 150:24:@5285.4]
  wire  x357_sum_1_reset; // @[Math.scala 150:24:@5285.4]
  wire [31:0] x357_sum_1_io_a; // @[Math.scala 150:24:@5285.4]
  wire [31:0] x357_sum_1_io_b; // @[Math.scala 150:24:@5285.4]
  wire  x357_sum_1_io_flow; // @[Math.scala 150:24:@5285.4]
  wire [31:0] x357_sum_1_io_result; // @[Math.scala 150:24:@5285.4]
  wire [31:0] x359_1_io_b; // @[Math.scala 720:24:@5306.4]
  wire [31:0] x359_1_io_result; // @[Math.scala 720:24:@5306.4]
  wire  x360_sum_1_clock; // @[Math.scala 150:24:@5317.4]
  wire  x360_sum_1_reset; // @[Math.scala 150:24:@5317.4]
  wire [31:0] x360_sum_1_io_a; // @[Math.scala 150:24:@5317.4]
  wire [31:0] x360_sum_1_io_b; // @[Math.scala 150:24:@5317.4]
  wire  x360_sum_1_io_flow; // @[Math.scala 150:24:@5317.4]
  wire [31:0] x360_sum_1_io_result; // @[Math.scala 150:24:@5317.4]
  wire [31:0] x362_1_io_b; // @[Math.scala 720:24:@5338.4]
  wire [31:0] x362_1_io_result; // @[Math.scala 720:24:@5338.4]
  wire  x363_sum_1_clock; // @[Math.scala 150:24:@5349.4]
  wire  x363_sum_1_reset; // @[Math.scala 150:24:@5349.4]
  wire [31:0] x363_sum_1_io_a; // @[Math.scala 150:24:@5349.4]
  wire [31:0] x363_sum_1_io_b; // @[Math.scala 150:24:@5349.4]
  wire  x363_sum_1_io_flow; // @[Math.scala 150:24:@5349.4]
  wire [31:0] x363_sum_1_io_result; // @[Math.scala 150:24:@5349.4]
  wire [31:0] x365_1_io_b; // @[Math.scala 720:24:@5370.4]
  wire [31:0] x365_1_io_result; // @[Math.scala 720:24:@5370.4]
  wire  x366_sum_1_clock; // @[Math.scala 150:24:@5381.4]
  wire  x366_sum_1_reset; // @[Math.scala 150:24:@5381.4]
  wire [31:0] x366_sum_1_io_a; // @[Math.scala 150:24:@5381.4]
  wire [31:0] x366_sum_1_io_b; // @[Math.scala 150:24:@5381.4]
  wire  x366_sum_1_io_flow; // @[Math.scala 150:24:@5381.4]
  wire [31:0] x366_sum_1_io_result; // @[Math.scala 150:24:@5381.4]
  wire [31:0] x368_1_io_b; // @[Math.scala 720:24:@5402.4]
  wire [31:0] x368_1_io_result; // @[Math.scala 720:24:@5402.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5421.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5421.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5421.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5421.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5421.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5430.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5430.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5430.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5430.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5430.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5441.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5441.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5441.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5441.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5441.4]
  wire  _T_327; // @[sm_x372_inr_Foreach.scala 62:18:@5240.4]
  wire  _T_328; // @[sm_x372_inr_Foreach.scala 62:55:@5241.4]
  wire [31:0] b351_number; // @[Math.scala 723:22:@5220.4 Math.scala 724:14:@5221.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@5245.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@5245.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@5250.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@5250.4]
  wire [31:0] x357_sum_number; // @[Math.scala 154:22:@5291.4 Math.scala 155:14:@5292.4]
  wire [31:0] _T_358; // @[Math.scala 406:49:@5298.4]
  wire [31:0] _T_360; // @[Math.scala 406:56:@5300.4]
  wire [31:0] _T_361; // @[Math.scala 406:56:@5301.4]
  wire [31:0] x360_sum_number; // @[Math.scala 154:22:@5323.4 Math.scala 155:14:@5324.4]
  wire [31:0] _T_380; // @[Math.scala 406:49:@5330.4]
  wire [31:0] _T_382; // @[Math.scala 406:56:@5332.4]
  wire [31:0] _T_383; // @[Math.scala 406:56:@5333.4]
  wire [31:0] x363_sum_number; // @[Math.scala 154:22:@5355.4 Math.scala 155:14:@5356.4]
  wire [31:0] _T_402; // @[Math.scala 406:49:@5362.4]
  wire [31:0] _T_404; // @[Math.scala 406:56:@5364.4]
  wire [31:0] _T_405; // @[Math.scala 406:56:@5365.4]
  wire [31:0] x366_sum_number; // @[Math.scala 154:22:@5387.4 Math.scala 155:14:@5388.4]
  wire [31:0] _T_424; // @[Math.scala 406:49:@5394.4]
  wire [31:0] _T_426; // @[Math.scala 406:56:@5396.4]
  wire [31:0] _T_427; // @[Math.scala 406:56:@5397.4]
  wire  _T_451; // @[sm_x372_inr_Foreach.scala 107:131:@5438.4]
  wire  _T_455; // @[package.scala 96:25:@5446.4 package.scala 96:25:@5447.4]
  wire  _T_457; // @[implicits.scala 55:10:@5448.4]
  wire  _T_458; // @[sm_x372_inr_Foreach.scala 107:148:@5449.4]
  wire  _T_460; // @[sm_x372_inr_Foreach.scala 107:236:@5451.4]
  wire  _T_461; // @[sm_x372_inr_Foreach.scala 107:255:@5452.4]
  wire  x744_b353_D3; // @[package.scala 96:25:@5435.4 package.scala 96:25:@5436.4]
  wire  _T_464; // @[sm_x372_inr_Foreach.scala 107:291:@5454.4]
  wire  x743_b354_D3; // @[package.scala 96:25:@5426.4 package.scala 96:25:@5427.4]
  _ _ ( // @[Math.scala 720:24:@5215.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@5227.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x720_sub x720_sub_1 ( // @[Math.scala 191:24:@5254.4]
    .clock(x720_sub_1_clock),
    .reset(x720_sub_1_reset),
    .io_a(x720_sub_1_io_a),
    .io_b(x720_sub_1_io_b),
    .io_flow(x720_sub_1_io_flow),
    .io_result(x720_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@5264.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x356_sum x356_sum_1 ( // @[Math.scala 150:24:@5273.4]
    .clock(x356_sum_1_clock),
    .reset(x356_sum_1_reset),
    .io_a(x356_sum_1_io_a),
    .io_b(x356_sum_1_io_b),
    .io_flow(x356_sum_1_io_flow),
    .io_result(x356_sum_1_io_result)
  );
  x356_sum x357_sum_1 ( // @[Math.scala 150:24:@5285.4]
    .clock(x357_sum_1_clock),
    .reset(x357_sum_1_reset),
    .io_a(x357_sum_1_io_a),
    .io_b(x357_sum_1_io_b),
    .io_flow(x357_sum_1_io_flow),
    .io_result(x357_sum_1_io_result)
  );
  _ x359_1 ( // @[Math.scala 720:24:@5306.4]
    .io_b(x359_1_io_b),
    .io_result(x359_1_io_result)
  );
  x356_sum x360_sum_1 ( // @[Math.scala 150:24:@5317.4]
    .clock(x360_sum_1_clock),
    .reset(x360_sum_1_reset),
    .io_a(x360_sum_1_io_a),
    .io_b(x360_sum_1_io_b),
    .io_flow(x360_sum_1_io_flow),
    .io_result(x360_sum_1_io_result)
  );
  _ x362_1 ( // @[Math.scala 720:24:@5338.4]
    .io_b(x362_1_io_b),
    .io_result(x362_1_io_result)
  );
  x356_sum x363_sum_1 ( // @[Math.scala 150:24:@5349.4]
    .clock(x363_sum_1_clock),
    .reset(x363_sum_1_reset),
    .io_a(x363_sum_1_io_a),
    .io_b(x363_sum_1_io_b),
    .io_flow(x363_sum_1_io_flow),
    .io_result(x363_sum_1_io_result)
  );
  _ x365_1 ( // @[Math.scala 720:24:@5370.4]
    .io_b(x365_1_io_b),
    .io_result(x365_1_io_result)
  );
  x356_sum x366_sum_1 ( // @[Math.scala 150:24:@5381.4]
    .clock(x366_sum_1_clock),
    .reset(x366_sum_1_reset),
    .io_a(x366_sum_1_io_a),
    .io_b(x366_sum_1_io_b),
    .io_flow(x366_sum_1_io_flow),
    .io_result(x366_sum_1_io_result)
  );
  _ x368_1 ( // @[Math.scala 720:24:@5402.4]
    .io_b(x368_1_io_b),
    .io_result(x368_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@5421.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@5430.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@5441.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x346_fifoinpacked_0_full; // @[sm_x372_inr_Foreach.scala 62:18:@5240.4]
  assign _T_328 = ~ io_in_x346_fifoinpacked_0_active_0_out; // @[sm_x372_inr_Foreach.scala 62:55:@5241.4]
  assign b351_number = __io_result; // @[Math.scala 723:22:@5220.4 Math.scala 724:14:@5221.4]
  assign _GEN_0 = {{11'd0}, b351_number}; // @[Math.scala 461:32:@5245.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@5245.4]
  assign _GEN_1 = {{7'd0}, b351_number}; // @[Math.scala 461:32:@5250.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@5250.4]
  assign x357_sum_number = x357_sum_1_io_result; // @[Math.scala 154:22:@5291.4 Math.scala 155:14:@5292.4]
  assign _T_358 = $signed(x357_sum_number); // @[Math.scala 406:49:@5298.4]
  assign _T_360 = $signed(_T_358) & $signed(32'shff); // @[Math.scala 406:56:@5300.4]
  assign _T_361 = $signed(_T_360); // @[Math.scala 406:56:@5301.4]
  assign x360_sum_number = x360_sum_1_io_result; // @[Math.scala 154:22:@5323.4 Math.scala 155:14:@5324.4]
  assign _T_380 = $signed(x360_sum_number); // @[Math.scala 406:49:@5330.4]
  assign _T_382 = $signed(_T_380) & $signed(32'shff); // @[Math.scala 406:56:@5332.4]
  assign _T_383 = $signed(_T_382); // @[Math.scala 406:56:@5333.4]
  assign x363_sum_number = x363_sum_1_io_result; // @[Math.scala 154:22:@5355.4 Math.scala 155:14:@5356.4]
  assign _T_402 = $signed(x363_sum_number); // @[Math.scala 406:49:@5362.4]
  assign _T_404 = $signed(_T_402) & $signed(32'shff); // @[Math.scala 406:56:@5364.4]
  assign _T_405 = $signed(_T_404); // @[Math.scala 406:56:@5365.4]
  assign x366_sum_number = x366_sum_1_io_result; // @[Math.scala 154:22:@5387.4 Math.scala 155:14:@5388.4]
  assign _T_424 = $signed(x366_sum_number); // @[Math.scala 406:49:@5394.4]
  assign _T_426 = $signed(_T_424) & $signed(32'shff); // @[Math.scala 406:56:@5396.4]
  assign _T_427 = $signed(_T_426); // @[Math.scala 406:56:@5397.4]
  assign _T_451 = ~ io_sigsIn_break; // @[sm_x372_inr_Foreach.scala 107:131:@5438.4]
  assign _T_455 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@5446.4 package.scala 96:25:@5447.4]
  assign _T_457 = io_rr ? _T_455 : 1'h0; // @[implicits.scala 55:10:@5448.4]
  assign _T_458 = _T_451 & _T_457; // @[sm_x372_inr_Foreach.scala 107:148:@5449.4]
  assign _T_460 = _T_458 & _T_451; // @[sm_x372_inr_Foreach.scala 107:236:@5451.4]
  assign _T_461 = _T_460 & io_sigsIn_backpressure; // @[sm_x372_inr_Foreach.scala 107:255:@5452.4]
  assign x744_b353_D3 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@5435.4 package.scala 96:25:@5436.4]
  assign _T_464 = _T_461 & x744_b353_D3; // @[sm_x372_inr_Foreach.scala 107:291:@5454.4]
  assign x743_b354_D3 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5426.4 package.scala 96:25:@5427.4]
  assign io_in_x346_fifoinpacked_0_wPort_0_en_0 = _T_464 & x743_b354_D3; // @[MemInterfaceType.scala 93:57:@5458.4]
  assign io_in_x346_fifoinpacked_0_active_0_in = x744_b353_D3 & x743_b354_D3; // @[MemInterfaceType.scala 147:18:@5461.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@5218.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@5230.4]
  assign x720_sub_1_clock = clock; // @[:@5255.4]
  assign x720_sub_1_reset = reset; // @[:@5256.4]
  assign x720_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@5257.4]
  assign x720_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@5258.4]
  assign x720_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@5259.4]
  assign RetimeWrapper_clock = clock; // @[:@5265.4]
  assign RetimeWrapper_reset = reset; // @[:@5266.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5268.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@5267.4]
  assign x356_sum_1_clock = clock; // @[:@5274.4]
  assign x356_sum_1_reset = reset; // @[:@5275.4]
  assign x356_sum_1_io_a = x720_sub_1_io_result; // @[Math.scala 151:17:@5276.4]
  assign x356_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@5277.4]
  assign x356_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5278.4]
  assign x357_sum_1_clock = clock; // @[:@5286.4]
  assign x357_sum_1_reset = reset; // @[:@5287.4]
  assign x357_sum_1_io_a = x356_sum_1_io_result; // @[Math.scala 151:17:@5288.4]
  assign x357_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@5289.4]
  assign x357_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5290.4]
  assign x359_1_io_b = $unsigned(_T_361); // @[Math.scala 721:17:@5309.4]
  assign x360_sum_1_clock = clock; // @[:@5318.4]
  assign x360_sum_1_reset = reset; // @[:@5319.4]
  assign x360_sum_1_io_a = x356_sum_1_io_result; // @[Math.scala 151:17:@5320.4]
  assign x360_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@5321.4]
  assign x360_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5322.4]
  assign x362_1_io_b = $unsigned(_T_383); // @[Math.scala 721:17:@5341.4]
  assign x363_sum_1_clock = clock; // @[:@5350.4]
  assign x363_sum_1_reset = reset; // @[:@5351.4]
  assign x363_sum_1_io_a = x356_sum_1_io_result; // @[Math.scala 151:17:@5352.4]
  assign x363_sum_1_io_b = 32'h3; // @[Math.scala 152:17:@5353.4]
  assign x363_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5354.4]
  assign x365_1_io_b = $unsigned(_T_405); // @[Math.scala 721:17:@5373.4]
  assign x366_sum_1_clock = clock; // @[:@5382.4]
  assign x366_sum_1_reset = reset; // @[:@5383.4]
  assign x366_sum_1_io_a = x356_sum_1_io_result; // @[Math.scala 151:17:@5384.4]
  assign x366_sum_1_io_b = 32'h4; // @[Math.scala 152:17:@5385.4]
  assign x366_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5386.4]
  assign x368_1_io_b = $unsigned(_T_427); // @[Math.scala 721:17:@5405.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5422.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5423.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5425.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@5424.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5431.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5432.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5434.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@5433.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5442.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5443.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5445.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5444.4]
endmodule
module RetimeWrapper_44( // @[:@6579.2]
  input   clock, // @[:@6580.4]
  input   reset, // @[:@6581.4]
  input   io_flow, // @[:@6582.4]
  input   io_in, // @[:@6582.4]
  output  io_out // @[:@6582.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6584.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6584.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6584.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6584.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6584.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6584.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(175)) sr ( // @[RetimeShiftRegister.scala 15:20:@6584.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6597.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6596.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6595.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6594.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6593.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6591.4]
endmodule
module RetimeWrapper_48( // @[:@6707.2]
  input   clock, // @[:@6708.4]
  input   reset, // @[:@6709.4]
  input   io_flow, // @[:@6710.4]
  input   io_in, // @[:@6710.4]
  output  io_out // @[:@6710.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6712.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6712.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6712.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6712.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6712.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6712.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(174)) sr ( // @[RetimeShiftRegister.scala 15:20:@6712.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6725.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6724.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6723.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6722.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6721.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6719.4]
endmodule
module x669_inr_Foreach_SAMPLER_BOX_sm( // @[:@6727.2]
  input   clock, // @[:@6728.4]
  input   reset, // @[:@6729.4]
  input   io_enable, // @[:@6730.4]
  output  io_done, // @[:@6730.4]
  output  io_doneLatch, // @[:@6730.4]
  input   io_ctrDone, // @[:@6730.4]
  output  io_datapathEn, // @[:@6730.4]
  output  io_ctrInc, // @[:@6730.4]
  output  io_ctrRst, // @[:@6730.4]
  input   io_parentAck, // @[:@6730.4]
  input   io_backpressure, // @[:@6730.4]
  input   io_break // @[:@6730.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6732.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6732.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6732.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6732.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6732.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6732.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6735.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6735.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6735.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6735.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6735.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6735.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6769.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6769.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6769.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6769.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6769.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6791.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6791.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6791.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6791.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6791.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6803.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6803.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6803.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6803.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6803.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6811.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6811.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6811.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6811.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6811.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6827.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6827.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6827.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6827.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6827.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6740.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6741.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6742.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6743.4]
  wire  _T_100; // @[package.scala 100:49:@6760.4]
  reg  _T_103; // @[package.scala 48:56:@6761.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6774.4 package.scala 96:25:@6775.4]
  wire  _T_110; // @[package.scala 100:49:@6776.4]
  reg  _T_113; // @[package.scala 48:56:@6777.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6779.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6784.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6785.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6788.4]
  wire  _T_124; // @[package.scala 96:25:@6796.4 package.scala 96:25:@6797.4]
  wire  _T_126; // @[package.scala 100:49:@6798.4]
  reg  _T_129; // @[package.scala 48:56:@6799.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6821.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6823.4]
  reg  _T_153; // @[package.scala 48:56:@6824.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6832.4 package.scala 96:25:@6833.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6834.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6835.4]
  SRFF active ( // @[Controllers.scala 261:22:@6732.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6735.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_44 RetimeWrapper ( // @[package.scala 93:22:@6769.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_1 ( // @[package.scala 93:22:@6791.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6803.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6811.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_4 ( // @[package.scala 93:22:@6827.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6740.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6741.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6742.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6743.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6760.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6774.4 package.scala 96:25:@6775.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6776.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6779.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6784.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6785.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6788.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6796.4 package.scala 96:25:@6797.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6798.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6823.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6832.4 package.scala 96:25:@6833.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6834.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6835.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6802.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6837.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6787.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6790.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6782.4]
  assign active_clock = clock; // @[:@6733.4]
  assign active_reset = reset; // @[:@6734.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6745.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6749.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6750.4]
  assign done_clock = clock; // @[:@6736.4]
  assign done_reset = reset; // @[:@6737.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6765.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6758.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6759.4]
  assign RetimeWrapper_clock = clock; // @[:@6770.4]
  assign RetimeWrapper_reset = reset; // @[:@6771.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6773.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6772.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6792.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6793.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6795.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6794.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6804.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6805.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6807.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6806.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6812.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6813.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6815.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6814.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6828.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6829.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6831.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6830.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_52( // @[:@7028.2]
  input          clock, // @[:@7029.4]
  input          reset, // @[:@7030.4]
  input          io_flow, // @[:@7031.4]
  input  [127:0] io_in, // @[:@7031.4]
  output [127:0] io_out // @[:@7031.4]
);
  wire [127:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7033.4]
  wire [127:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7033.4]
  wire [127:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7033.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7033.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7033.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7033.4]
  RetimeShiftRegister #(.WIDTH(128), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7033.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7046.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7045.4]
  assign sr_init = 128'h0; // @[RetimeShiftRegister.scala 19:16:@7044.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7043.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7042.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7040.4]
endmodule
module SRAM_1( // @[:@7064.2]
  input         clock, // @[:@7065.4]
  input         reset, // @[:@7066.4]
  input  [8:0]  io_raddr, // @[:@7067.4]
  input         io_wen, // @[:@7067.4]
  input  [8:0]  io_waddr, // @[:@7067.4]
  input  [31:0] io_wdata, // @[:@7067.4]
  output [31:0] io_rdata, // @[:@7067.4]
  input         io_backpressure // @[:@7067.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@7069.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@7069.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@7069.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@7069.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@7069.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@7069.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@7069.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@7069.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@7069.4]
  wire  _T_19; // @[SRAM.scala 182:49:@7087.4]
  wire  _T_20; // @[SRAM.scala 182:37:@7088.4]
  reg  _T_23; // @[SRAM.scala 182:29:@7089.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@7091.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(320), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@7069.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@7087.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@7088.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@7096.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@7083.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@7084.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@7081.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@7086.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@7085.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@7082.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@7080.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@7079.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_53( // @[:@7110.2]
  input        clock, // @[:@7111.4]
  input        reset, // @[:@7112.4]
  input        io_flow, // @[:@7113.4]
  input  [8:0] io_in, // @[:@7113.4]
  output [8:0] io_out // @[:@7113.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7115.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7115.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7115.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7115.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7115.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7115.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7115.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7128.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7127.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@7126.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7125.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7124.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7122.4]
endmodule
module Mem1D_5( // @[:@7130.2]
  input         clock, // @[:@7131.4]
  input         reset, // @[:@7132.4]
  input  [8:0]  io_r_ofs_0, // @[:@7133.4]
  input         io_r_backpressure, // @[:@7133.4]
  input  [8:0]  io_w_ofs_0, // @[:@7133.4]
  input  [31:0] io_w_data_0, // @[:@7133.4]
  input         io_w_en_0, // @[:@7133.4]
  output [31:0] io_output // @[:@7133.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@7137.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@7137.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@7137.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@7137.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@7137.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@7137.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@7137.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@7137.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7140.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7140.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7140.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7140.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7140.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@7135.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@7137.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_53 RetimeWrapper ( // @[package.scala 93:22:@7140.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h140; // @[MemPrimitives.scala 702:32:@7135.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@7153.4]
  assign SRAM_clock = clock; // @[:@7138.4]
  assign SRAM_reset = reset; // @[:@7139.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@7147.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@7150.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@7148.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@7151.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@7152.4]
  assign RetimeWrapper_clock = clock; // @[:@7141.4]
  assign RetimeWrapper_reset = reset; // @[:@7142.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@7144.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@7143.4]
endmodule
module StickySelects_1( // @[:@9616.2]
  input   clock, // @[:@9617.4]
  input   reset, // @[:@9618.4]
  input   io_ins_0, // @[:@9619.4]
  input   io_ins_1, // @[:@9619.4]
  input   io_ins_2, // @[:@9619.4]
  input   io_ins_3, // @[:@9619.4]
  input   io_ins_4, // @[:@9619.4]
  input   io_ins_5, // @[:@9619.4]
  input   io_ins_6, // @[:@9619.4]
  input   io_ins_7, // @[:@9619.4]
  input   io_ins_8, // @[:@9619.4]
  output  io_outs_0, // @[:@9619.4]
  output  io_outs_1, // @[:@9619.4]
  output  io_outs_2, // @[:@9619.4]
  output  io_outs_3, // @[:@9619.4]
  output  io_outs_4, // @[:@9619.4]
  output  io_outs_5, // @[:@9619.4]
  output  io_outs_6, // @[:@9619.4]
  output  io_outs_7, // @[:@9619.4]
  output  io_outs_8 // @[:@9619.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@9621.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@9622.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@9623.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@9624.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@9625.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@9626.4]
  reg [31:0] _RAND_5;
  reg  _T_37; // @[StickySelects.scala 37:46:@9627.4]
  reg [31:0] _RAND_6;
  reg  _T_40; // @[StickySelects.scala 37:46:@9628.4]
  reg [31:0] _RAND_7;
  reg  _T_43; // @[StickySelects.scala 37:46:@9629.4]
  reg [31:0] _RAND_8;
  wire  _T_44; // @[StickySelects.scala 47:46:@9630.4]
  wire  _T_45; // @[StickySelects.scala 47:46:@9631.4]
  wire  _T_46; // @[StickySelects.scala 47:46:@9632.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@9633.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@9634.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@9635.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@9636.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@9637.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@9638.4]
  wire  _T_53; // @[StickySelects.scala 47:46:@9640.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@9641.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@9642.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@9643.4]
  wire  _T_57; // @[StickySelects.scala 47:46:@9644.4]
  wire  _T_58; // @[StickySelects.scala 47:46:@9645.4]
  wire  _T_59; // @[StickySelects.scala 47:46:@9646.4]
  wire  _T_60; // @[StickySelects.scala 49:53:@9647.4]
  wire  _T_61; // @[StickySelects.scala 49:21:@9648.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@9650.4]
  wire  _T_63; // @[StickySelects.scala 47:46:@9651.4]
  wire  _T_64; // @[StickySelects.scala 47:46:@9652.4]
  wire  _T_65; // @[StickySelects.scala 47:46:@9653.4]
  wire  _T_66; // @[StickySelects.scala 47:46:@9654.4]
  wire  _T_67; // @[StickySelects.scala 47:46:@9655.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@9656.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@9657.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@9658.4]
  wire  _T_72; // @[StickySelects.scala 47:46:@9661.4]
  wire  _T_73; // @[StickySelects.scala 47:46:@9662.4]
  wire  _T_74; // @[StickySelects.scala 47:46:@9663.4]
  wire  _T_75; // @[StickySelects.scala 47:46:@9664.4]
  wire  _T_76; // @[StickySelects.scala 47:46:@9665.4]
  wire  _T_77; // @[StickySelects.scala 47:46:@9666.4]
  wire  _T_78; // @[StickySelects.scala 49:53:@9667.4]
  wire  _T_79; // @[StickySelects.scala 49:21:@9668.4]
  wire  _T_82; // @[StickySelects.scala 47:46:@9672.4]
  wire  _T_83; // @[StickySelects.scala 47:46:@9673.4]
  wire  _T_84; // @[StickySelects.scala 47:46:@9674.4]
  wire  _T_85; // @[StickySelects.scala 47:46:@9675.4]
  wire  _T_86; // @[StickySelects.scala 47:46:@9676.4]
  wire  _T_87; // @[StickySelects.scala 49:53:@9677.4]
  wire  _T_88; // @[StickySelects.scala 49:21:@9678.4]
  wire  _T_92; // @[StickySelects.scala 47:46:@9683.4]
  wire  _T_93; // @[StickySelects.scala 47:46:@9684.4]
  wire  _T_94; // @[StickySelects.scala 47:46:@9685.4]
  wire  _T_95; // @[StickySelects.scala 47:46:@9686.4]
  wire  _T_96; // @[StickySelects.scala 49:53:@9687.4]
  wire  _T_97; // @[StickySelects.scala 49:21:@9688.4]
  wire  _T_102; // @[StickySelects.scala 47:46:@9694.4]
  wire  _T_103; // @[StickySelects.scala 47:46:@9695.4]
  wire  _T_104; // @[StickySelects.scala 47:46:@9696.4]
  wire  _T_105; // @[StickySelects.scala 49:53:@9697.4]
  wire  _T_106; // @[StickySelects.scala 49:21:@9698.4]
  wire  _T_112; // @[StickySelects.scala 47:46:@9705.4]
  wire  _T_113; // @[StickySelects.scala 47:46:@9706.4]
  wire  _T_114; // @[StickySelects.scala 49:53:@9707.4]
  wire  _T_115; // @[StickySelects.scala 49:21:@9708.4]
  wire  _T_122; // @[StickySelects.scala 47:46:@9716.4]
  wire  _T_123; // @[StickySelects.scala 49:53:@9717.4]
  wire  _T_124; // @[StickySelects.scala 49:21:@9718.4]
  assign _T_44 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@9630.4]
  assign _T_45 = _T_44 | io_ins_3; // @[StickySelects.scala 47:46:@9631.4]
  assign _T_46 = _T_45 | io_ins_4; // @[StickySelects.scala 47:46:@9632.4]
  assign _T_47 = _T_46 | io_ins_5; // @[StickySelects.scala 47:46:@9633.4]
  assign _T_48 = _T_47 | io_ins_6; // @[StickySelects.scala 47:46:@9634.4]
  assign _T_49 = _T_48 | io_ins_7; // @[StickySelects.scala 47:46:@9635.4]
  assign _T_50 = _T_49 | io_ins_8; // @[StickySelects.scala 47:46:@9636.4]
  assign _T_51 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@9637.4]
  assign _T_52 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 49:21:@9638.4]
  assign _T_53 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@9640.4]
  assign _T_54 = _T_53 | io_ins_3; // @[StickySelects.scala 47:46:@9641.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@9642.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@9643.4]
  assign _T_57 = _T_56 | io_ins_6; // @[StickySelects.scala 47:46:@9644.4]
  assign _T_58 = _T_57 | io_ins_7; // @[StickySelects.scala 47:46:@9645.4]
  assign _T_59 = _T_58 | io_ins_8; // @[StickySelects.scala 47:46:@9646.4]
  assign _T_60 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@9647.4]
  assign _T_61 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 49:21:@9648.4]
  assign _T_62 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@9650.4]
  assign _T_63 = _T_62 | io_ins_3; // @[StickySelects.scala 47:46:@9651.4]
  assign _T_64 = _T_63 | io_ins_4; // @[StickySelects.scala 47:46:@9652.4]
  assign _T_65 = _T_64 | io_ins_5; // @[StickySelects.scala 47:46:@9653.4]
  assign _T_66 = _T_65 | io_ins_6; // @[StickySelects.scala 47:46:@9654.4]
  assign _T_67 = _T_66 | io_ins_7; // @[StickySelects.scala 47:46:@9655.4]
  assign _T_68 = _T_67 | io_ins_8; // @[StickySelects.scala 47:46:@9656.4]
  assign _T_69 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@9657.4]
  assign _T_70 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 49:21:@9658.4]
  assign _T_72 = _T_62 | io_ins_2; // @[StickySelects.scala 47:46:@9661.4]
  assign _T_73 = _T_72 | io_ins_4; // @[StickySelects.scala 47:46:@9662.4]
  assign _T_74 = _T_73 | io_ins_5; // @[StickySelects.scala 47:46:@9663.4]
  assign _T_75 = _T_74 | io_ins_6; // @[StickySelects.scala 47:46:@9664.4]
  assign _T_76 = _T_75 | io_ins_7; // @[StickySelects.scala 47:46:@9665.4]
  assign _T_77 = _T_76 | io_ins_8; // @[StickySelects.scala 47:46:@9666.4]
  assign _T_78 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@9667.4]
  assign _T_79 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 49:21:@9668.4]
  assign _T_82 = _T_72 | io_ins_3; // @[StickySelects.scala 47:46:@9672.4]
  assign _T_83 = _T_82 | io_ins_5; // @[StickySelects.scala 47:46:@9673.4]
  assign _T_84 = _T_83 | io_ins_6; // @[StickySelects.scala 47:46:@9674.4]
  assign _T_85 = _T_84 | io_ins_7; // @[StickySelects.scala 47:46:@9675.4]
  assign _T_86 = _T_85 | io_ins_8; // @[StickySelects.scala 47:46:@9676.4]
  assign _T_87 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@9677.4]
  assign _T_88 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 49:21:@9678.4]
  assign _T_92 = _T_82 | io_ins_4; // @[StickySelects.scala 47:46:@9683.4]
  assign _T_93 = _T_92 | io_ins_6; // @[StickySelects.scala 47:46:@9684.4]
  assign _T_94 = _T_93 | io_ins_7; // @[StickySelects.scala 47:46:@9685.4]
  assign _T_95 = _T_94 | io_ins_8; // @[StickySelects.scala 47:46:@9686.4]
  assign _T_96 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@9687.4]
  assign _T_97 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 49:21:@9688.4]
  assign _T_102 = _T_92 | io_ins_5; // @[StickySelects.scala 47:46:@9694.4]
  assign _T_103 = _T_102 | io_ins_7; // @[StickySelects.scala 47:46:@9695.4]
  assign _T_104 = _T_103 | io_ins_8; // @[StickySelects.scala 47:46:@9696.4]
  assign _T_105 = io_ins_6 | _T_37; // @[StickySelects.scala 49:53:@9697.4]
  assign _T_106 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 49:21:@9698.4]
  assign _T_112 = _T_102 | io_ins_6; // @[StickySelects.scala 47:46:@9705.4]
  assign _T_113 = _T_112 | io_ins_8; // @[StickySelects.scala 47:46:@9706.4]
  assign _T_114 = io_ins_7 | _T_40; // @[StickySelects.scala 49:53:@9707.4]
  assign _T_115 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 49:21:@9708.4]
  assign _T_122 = _T_112 | io_ins_7; // @[StickySelects.scala 47:46:@9716.4]
  assign _T_123 = io_ins_8 | _T_43; // @[StickySelects.scala 49:53:@9717.4]
  assign _T_124 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 49:21:@9718.4]
  assign io_outs_0 = _T_50 ? io_ins_0 : _T_51; // @[StickySelects.scala 53:57:@9720.4]
  assign io_outs_1 = _T_59 ? io_ins_1 : _T_60; // @[StickySelects.scala 53:57:@9721.4]
  assign io_outs_2 = _T_68 ? io_ins_2 : _T_69; // @[StickySelects.scala 53:57:@9722.4]
  assign io_outs_3 = _T_77 ? io_ins_3 : _T_78; // @[StickySelects.scala 53:57:@9723.4]
  assign io_outs_4 = _T_86 ? io_ins_4 : _T_87; // @[StickySelects.scala 53:57:@9724.4]
  assign io_outs_5 = _T_95 ? io_ins_5 : _T_96; // @[StickySelects.scala 53:57:@9725.4]
  assign io_outs_6 = _T_104 ? io_ins_6 : _T_105; // @[StickySelects.scala 53:57:@9726.4]
  assign io_outs_7 = _T_113 ? io_ins_7 : _T_114; // @[StickySelects.scala 53:57:@9727.4]
  assign io_outs_8 = _T_122 ? io_ins_8 : _T_123; // @[StickySelects.scala 53:57:@9728.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_37 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_40 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_43 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_51;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_59) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_60;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_69;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_77) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_78;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_86) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_87;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_95) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_96;
      end
    end
    if (reset) begin
      _T_37 <= 1'h0;
    end else begin
      if (_T_104) begin
        _T_37 <= io_ins_6;
      end else begin
        _T_37 <= _T_105;
      end
    end
    if (reset) begin
      _T_40 <= 1'h0;
    end else begin
      if (_T_113) begin
        _T_40 <= io_ins_7;
      end else begin
        _T_40 <= _T_114;
      end
    end
    if (reset) begin
      _T_43 <= 1'h0;
    end else begin
      if (_T_122) begin
        _T_43 <= io_ins_8;
      end else begin
        _T_43 <= _T_123;
      end
    end
  end
endmodule
module x383_lb_0( // @[:@19264.2]
  input         clock, // @[:@19265.4]
  input         reset, // @[:@19266.4]
  input  [2:0]  io_rPort_17_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_17_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_17_ofs_0, // @[:@19267.4]
  input         io_rPort_17_en_0, // @[:@19267.4]
  input         io_rPort_17_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_17_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_16_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_16_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_16_ofs_0, // @[:@19267.4]
  input         io_rPort_16_en_0, // @[:@19267.4]
  input         io_rPort_16_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_16_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_15_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_15_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_15_ofs_0, // @[:@19267.4]
  input         io_rPort_15_en_0, // @[:@19267.4]
  input         io_rPort_15_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_15_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_14_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_14_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_14_ofs_0, // @[:@19267.4]
  input         io_rPort_14_en_0, // @[:@19267.4]
  input         io_rPort_14_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_14_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_13_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_13_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_13_ofs_0, // @[:@19267.4]
  input         io_rPort_13_en_0, // @[:@19267.4]
  input         io_rPort_13_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_13_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_12_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_12_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_12_ofs_0, // @[:@19267.4]
  input         io_rPort_12_en_0, // @[:@19267.4]
  input         io_rPort_12_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_12_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_11_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_11_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_11_ofs_0, // @[:@19267.4]
  input         io_rPort_11_en_0, // @[:@19267.4]
  input         io_rPort_11_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_11_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_10_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_10_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_10_ofs_0, // @[:@19267.4]
  input         io_rPort_10_en_0, // @[:@19267.4]
  input         io_rPort_10_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_10_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@19267.4]
  input         io_rPort_9_en_0, // @[:@19267.4]
  input         io_rPort_9_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_9_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@19267.4]
  input         io_rPort_8_en_0, // @[:@19267.4]
  input         io_rPort_8_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_8_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@19267.4]
  input         io_rPort_7_en_0, // @[:@19267.4]
  input         io_rPort_7_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_7_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@19267.4]
  input         io_rPort_6_en_0, // @[:@19267.4]
  input         io_rPort_6_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_6_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@19267.4]
  input         io_rPort_5_en_0, // @[:@19267.4]
  input         io_rPort_5_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_5_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@19267.4]
  input         io_rPort_4_en_0, // @[:@19267.4]
  input         io_rPort_4_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_4_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@19267.4]
  input         io_rPort_3_en_0, // @[:@19267.4]
  input         io_rPort_3_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_3_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@19267.4]
  input         io_rPort_2_en_0, // @[:@19267.4]
  input         io_rPort_2_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_2_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@19267.4]
  input         io_rPort_1_en_0, // @[:@19267.4]
  input         io_rPort_1_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_1_output_0, // @[:@19267.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@19267.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@19267.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@19267.4]
  input         io_rPort_0_en_0, // @[:@19267.4]
  input         io_rPort_0_backpressure, // @[:@19267.4]
  output [31:0] io_rPort_0_output_0, // @[:@19267.4]
  input  [2:0]  io_wPort_3_banks_1, // @[:@19267.4]
  input  [2:0]  io_wPort_3_banks_0, // @[:@19267.4]
  input  [8:0]  io_wPort_3_ofs_0, // @[:@19267.4]
  input  [31:0] io_wPort_3_data_0, // @[:@19267.4]
  input         io_wPort_3_en_0, // @[:@19267.4]
  input  [2:0]  io_wPort_2_banks_1, // @[:@19267.4]
  input  [2:0]  io_wPort_2_banks_0, // @[:@19267.4]
  input  [8:0]  io_wPort_2_ofs_0, // @[:@19267.4]
  input  [31:0] io_wPort_2_data_0, // @[:@19267.4]
  input         io_wPort_2_en_0, // @[:@19267.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@19267.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@19267.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@19267.4]
  input  [31:0] io_wPort_1_data_0, // @[:@19267.4]
  input         io_wPort_1_en_0, // @[:@19267.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@19267.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@19267.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@19267.4]
  input  [31:0] io_wPort_0_data_0, // @[:@19267.4]
  input         io_wPort_0_en_0 // @[:@19267.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@19410.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@19410.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19410.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19410.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19410.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@19410.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@19410.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@19410.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@19426.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@19426.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19426.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19426.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19426.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@19426.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@19426.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@19426.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@19442.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@19442.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19442.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19442.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19442.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@19442.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@19442.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@19442.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@19458.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@19458.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19458.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19458.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19458.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@19458.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@19458.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@19458.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@19474.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@19474.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19474.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19474.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19474.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@19474.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@19474.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@19474.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@19490.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@19490.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19490.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19490.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19490.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@19490.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@19490.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@19490.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@19506.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@19506.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19506.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19506.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19506.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@19506.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@19506.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@19506.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@19522.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@19522.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19522.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19522.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19522.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@19522.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@19522.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@19522.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@19538.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@19538.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19538.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19538.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19538.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@19538.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@19538.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@19538.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@19554.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@19554.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19554.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19554.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19554.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@19554.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@19554.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@19554.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@19570.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@19570.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19570.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19570.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19570.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@19570.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@19570.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@19570.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@19586.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@19586.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19586.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19586.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19586.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@19586.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@19586.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@19586.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@19602.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@19602.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19602.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19602.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19602.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@19602.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@19602.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@19602.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@19618.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@19618.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19618.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19618.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19618.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@19618.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@19618.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@19618.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@19634.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@19634.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19634.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19634.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19634.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@19634.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@19634.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@19634.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@19650.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@19650.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19650.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19650.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19650.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@19650.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@19650.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@19650.4]
  wire  Mem1D_16_clock; // @[MemPrimitives.scala 64:21:@19666.4]
  wire  Mem1D_16_reset; // @[MemPrimitives.scala 64:21:@19666.4]
  wire [8:0] Mem1D_16_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19666.4]
  wire  Mem1D_16_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19666.4]
  wire [8:0] Mem1D_16_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19666.4]
  wire [31:0] Mem1D_16_io_w_data_0; // @[MemPrimitives.scala 64:21:@19666.4]
  wire  Mem1D_16_io_w_en_0; // @[MemPrimitives.scala 64:21:@19666.4]
  wire [31:0] Mem1D_16_io_output; // @[MemPrimitives.scala 64:21:@19666.4]
  wire  Mem1D_17_clock; // @[MemPrimitives.scala 64:21:@19682.4]
  wire  Mem1D_17_reset; // @[MemPrimitives.scala 64:21:@19682.4]
  wire [8:0] Mem1D_17_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19682.4]
  wire  Mem1D_17_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19682.4]
  wire [8:0] Mem1D_17_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19682.4]
  wire [31:0] Mem1D_17_io_w_data_0; // @[MemPrimitives.scala 64:21:@19682.4]
  wire  Mem1D_17_io_w_en_0; // @[MemPrimitives.scala 64:21:@19682.4]
  wire [31:0] Mem1D_17_io_output; // @[MemPrimitives.scala 64:21:@19682.4]
  wire  Mem1D_18_clock; // @[MemPrimitives.scala 64:21:@19698.4]
  wire  Mem1D_18_reset; // @[MemPrimitives.scala 64:21:@19698.4]
  wire [8:0] Mem1D_18_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19698.4]
  wire  Mem1D_18_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19698.4]
  wire [8:0] Mem1D_18_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19698.4]
  wire [31:0] Mem1D_18_io_w_data_0; // @[MemPrimitives.scala 64:21:@19698.4]
  wire  Mem1D_18_io_w_en_0; // @[MemPrimitives.scala 64:21:@19698.4]
  wire [31:0] Mem1D_18_io_output; // @[MemPrimitives.scala 64:21:@19698.4]
  wire  Mem1D_19_clock; // @[MemPrimitives.scala 64:21:@19714.4]
  wire  Mem1D_19_reset; // @[MemPrimitives.scala 64:21:@19714.4]
  wire [8:0] Mem1D_19_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19714.4]
  wire  Mem1D_19_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19714.4]
  wire [8:0] Mem1D_19_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19714.4]
  wire [31:0] Mem1D_19_io_w_data_0; // @[MemPrimitives.scala 64:21:@19714.4]
  wire  Mem1D_19_io_w_en_0; // @[MemPrimitives.scala 64:21:@19714.4]
  wire [31:0] Mem1D_19_io_output; // @[MemPrimitives.scala 64:21:@19714.4]
  wire  Mem1D_20_clock; // @[MemPrimitives.scala 64:21:@19730.4]
  wire  Mem1D_20_reset; // @[MemPrimitives.scala 64:21:@19730.4]
  wire [8:0] Mem1D_20_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19730.4]
  wire  Mem1D_20_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19730.4]
  wire [8:0] Mem1D_20_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19730.4]
  wire [31:0] Mem1D_20_io_w_data_0; // @[MemPrimitives.scala 64:21:@19730.4]
  wire  Mem1D_20_io_w_en_0; // @[MemPrimitives.scala 64:21:@19730.4]
  wire [31:0] Mem1D_20_io_output; // @[MemPrimitives.scala 64:21:@19730.4]
  wire  Mem1D_21_clock; // @[MemPrimitives.scala 64:21:@19746.4]
  wire  Mem1D_21_reset; // @[MemPrimitives.scala 64:21:@19746.4]
  wire [8:0] Mem1D_21_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19746.4]
  wire  Mem1D_21_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19746.4]
  wire [8:0] Mem1D_21_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19746.4]
  wire [31:0] Mem1D_21_io_w_data_0; // @[MemPrimitives.scala 64:21:@19746.4]
  wire  Mem1D_21_io_w_en_0; // @[MemPrimitives.scala 64:21:@19746.4]
  wire [31:0] Mem1D_21_io_output; // @[MemPrimitives.scala 64:21:@19746.4]
  wire  Mem1D_22_clock; // @[MemPrimitives.scala 64:21:@19762.4]
  wire  Mem1D_22_reset; // @[MemPrimitives.scala 64:21:@19762.4]
  wire [8:0] Mem1D_22_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19762.4]
  wire  Mem1D_22_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19762.4]
  wire [8:0] Mem1D_22_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19762.4]
  wire [31:0] Mem1D_22_io_w_data_0; // @[MemPrimitives.scala 64:21:@19762.4]
  wire  Mem1D_22_io_w_en_0; // @[MemPrimitives.scala 64:21:@19762.4]
  wire [31:0] Mem1D_22_io_output; // @[MemPrimitives.scala 64:21:@19762.4]
  wire  Mem1D_23_clock; // @[MemPrimitives.scala 64:21:@19778.4]
  wire  Mem1D_23_reset; // @[MemPrimitives.scala 64:21:@19778.4]
  wire [8:0] Mem1D_23_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@19778.4]
  wire  Mem1D_23_io_r_backpressure; // @[MemPrimitives.scala 64:21:@19778.4]
  wire [8:0] Mem1D_23_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@19778.4]
  wire [31:0] Mem1D_23_io_w_data_0; // @[MemPrimitives.scala 64:21:@19778.4]
  wire  Mem1D_23_io_w_en_0; // @[MemPrimitives.scala 64:21:@19778.4]
  wire [31:0] Mem1D_23_io_output; // @[MemPrimitives.scala 64:21:@19778.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_6; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_7; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_ins_8; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_6; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_7; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_io_outs_8; // @[MemPrimitives.scala 124:33:@20286.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_6; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_7; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_ins_8; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_6; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_7; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_1_io_outs_8; // @[MemPrimitives.scala 124:33:@20375.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_6; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_7; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_ins_8; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_6; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_7; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_2_io_outs_8; // @[MemPrimitives.scala 124:33:@20464.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_6; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_7; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_ins_8; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_6; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_7; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_3_io_outs_8; // @[MemPrimitives.scala 124:33:@20553.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_6; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_7; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_ins_8; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_6; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_7; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_4_io_outs_8; // @[MemPrimitives.scala 124:33:@20642.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_6; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_7; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_ins_8; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_6; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_7; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_5_io_outs_8; // @[MemPrimitives.scala 124:33:@20731.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_6; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_7; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_ins_8; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_6; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_7; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_6_io_outs_8; // @[MemPrimitives.scala 124:33:@20820.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_6; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_7; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_ins_8; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_6; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_7; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_7_io_outs_8; // @[MemPrimitives.scala 124:33:@20909.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_6; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_7; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_ins_8; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_6; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_7; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_8_io_outs_8; // @[MemPrimitives.scala 124:33:@20998.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_6; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_7; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_ins_8; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_6; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_7; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_9_io_outs_8; // @[MemPrimitives.scala 124:33:@21087.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_6; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_7; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_ins_8; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_6; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_7; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_10_io_outs_8; // @[MemPrimitives.scala 124:33:@21176.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_6; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_7; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_ins_8; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_6; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_7; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_11_io_outs_8; // @[MemPrimitives.scala 124:33:@21265.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_6; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_7; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_ins_8; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_6; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_7; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_12_io_outs_8; // @[MemPrimitives.scala 124:33:@21354.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_6; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_7; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_ins_8; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_6; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_7; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_13_io_outs_8; // @[MemPrimitives.scala 124:33:@21443.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_6; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_7; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_ins_8; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_6; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_7; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_14_io_outs_8; // @[MemPrimitives.scala 124:33:@21532.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_6; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_7; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_ins_8; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_6; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_7; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_15_io_outs_8; // @[MemPrimitives.scala 124:33:@21621.4]
  wire  StickySelects_16_clock; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_reset; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_0; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_1; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_2; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_3; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_4; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_5; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_6; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_7; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_ins_8; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_0; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_1; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_2; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_3; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_4; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_5; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_6; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_7; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_16_io_outs_8; // @[MemPrimitives.scala 124:33:@21710.4]
  wire  StickySelects_17_clock; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_reset; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_0; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_1; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_2; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_3; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_4; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_5; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_6; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_7; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_ins_8; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_0; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_1; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_2; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_3; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_4; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_5; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_6; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_7; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_17_io_outs_8; // @[MemPrimitives.scala 124:33:@21799.4]
  wire  StickySelects_18_clock; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_reset; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_0; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_1; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_2; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_3; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_4; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_5; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_6; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_7; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_ins_8; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_0; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_1; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_2; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_3; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_4; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_5; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_6; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_7; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_18_io_outs_8; // @[MemPrimitives.scala 124:33:@21888.4]
  wire  StickySelects_19_clock; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_reset; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_0; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_1; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_2; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_3; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_4; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_5; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_6; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_7; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_ins_8; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_0; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_1; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_2; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_3; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_4; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_5; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_6; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_7; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_19_io_outs_8; // @[MemPrimitives.scala 124:33:@21977.4]
  wire  StickySelects_20_clock; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_reset; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_0; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_1; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_2; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_3; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_4; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_5; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_6; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_7; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_ins_8; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_0; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_1; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_2; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_3; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_4; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_5; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_6; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_7; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_20_io_outs_8; // @[MemPrimitives.scala 124:33:@22066.4]
  wire  StickySelects_21_clock; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_reset; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_0; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_1; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_2; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_3; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_4; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_5; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_6; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_7; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_ins_8; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_0; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_1; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_2; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_3; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_4; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_5; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_6; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_7; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_21_io_outs_8; // @[MemPrimitives.scala 124:33:@22155.4]
  wire  StickySelects_22_clock; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_reset; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_0; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_1; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_2; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_3; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_4; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_5; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_6; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_7; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_ins_8; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_0; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_1; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_2; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_3; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_4; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_5; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_6; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_7; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_22_io_outs_8; // @[MemPrimitives.scala 124:33:@22244.4]
  wire  StickySelects_23_clock; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_reset; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_0; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_1; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_2; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_3; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_4; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_5; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_6; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_7; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_ins_8; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_0; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_1; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_2; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_3; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_4; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_5; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_6; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_7; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  StickySelects_23_io_outs_8; // @[MemPrimitives.scala 124:33:@22333.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@22423.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@22423.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@22423.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@22423.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@22423.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@22431.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@22431.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@22431.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@22431.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@22431.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@22439.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@22447.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@22447.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@22447.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@22447.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@22447.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@22455.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@22455.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@22455.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@22455.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@22455.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@22463.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@22463.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@22463.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@22463.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@22463.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@22471.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@22471.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@22471.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@22471.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@22471.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@22479.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@22479.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@22479.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@22479.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@22479.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@22487.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@22487.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@22487.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@22487.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@22487.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@22495.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@22495.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@22495.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@22495.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@22495.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@22503.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@22503.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@22503.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@22503.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@22503.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@22511.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@22511.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@22511.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@22511.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@22511.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@22567.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@22567.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@22567.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@22567.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@22567.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@22575.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@22575.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@22575.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@22575.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@22575.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@22583.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@22583.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@22583.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@22583.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@22583.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@22591.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@22591.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@22591.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@22591.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@22591.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@22599.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@22599.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@22599.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@22599.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@22599.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@22607.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@22607.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@22607.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@22607.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@22607.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@22615.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@22615.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@22615.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@22615.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@22615.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@22623.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@22623.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@22623.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@22623.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@22623.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@22631.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@22631.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@22631.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@22631.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@22631.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@22639.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@22639.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@22639.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@22639.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@22639.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@22647.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@22647.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@22647.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@22647.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@22647.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@22655.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@22655.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@22655.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@22655.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@22655.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@22711.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@22711.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@22711.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@22711.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@22711.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@22719.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@22719.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@22719.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@22719.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@22719.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@22727.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@22727.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@22727.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@22727.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@22727.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@22735.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@22735.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@22735.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@22735.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@22735.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@22743.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@22743.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@22743.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@22743.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@22743.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@22751.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@22751.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@22751.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@22751.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@22751.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@22759.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@22759.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@22759.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@22759.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@22759.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@22767.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@22767.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@22767.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@22767.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@22767.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@22775.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@22775.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@22775.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@22775.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@22775.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@22783.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@22783.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@22783.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@22783.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@22783.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@22791.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@22791.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@22791.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@22791.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@22791.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@22799.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@22799.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@22799.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@22799.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@22799.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@22855.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@22855.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@22855.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@22855.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@22855.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@22863.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@22863.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@22863.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@22863.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@22863.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@22871.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@22871.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@22871.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@22871.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@22871.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@22879.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@22879.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@22879.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@22879.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@22879.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@22887.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@22887.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@22887.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@22887.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@22887.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@22895.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@22895.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@22895.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@22895.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@22895.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@22903.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@22903.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@22903.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@22903.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@22903.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@22911.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@22911.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@22911.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@22911.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@22911.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@22919.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@22919.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@22919.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@22919.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@22919.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@22927.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@22927.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@22927.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@22927.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@22927.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@22935.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@22935.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@22935.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@22935.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@22935.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@22943.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@22943.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@22943.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@22943.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@22943.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@22999.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@22999.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@22999.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@22999.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@22999.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@23007.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@23007.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@23007.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@23007.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@23007.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@23015.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@23015.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@23015.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@23015.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@23015.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@23023.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@23023.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@23023.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@23023.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@23023.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@23031.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@23031.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@23031.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@23031.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@23031.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@23039.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@23039.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@23039.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@23039.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@23039.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@23047.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@23047.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@23047.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@23047.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@23047.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@23055.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@23055.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@23055.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@23055.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@23055.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@23063.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@23063.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@23063.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@23063.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@23063.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@23071.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@23071.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@23071.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@23071.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@23071.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@23079.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@23079.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@23079.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@23079.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@23079.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@23087.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@23087.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@23087.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@23087.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@23087.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@23143.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@23143.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@23143.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@23143.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@23143.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@23151.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@23151.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@23151.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@23151.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@23151.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@23159.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@23159.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@23159.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@23159.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@23159.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@23167.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@23167.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@23167.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@23167.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@23167.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@23175.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@23175.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@23175.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@23175.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@23175.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@23183.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@23183.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@23183.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@23183.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@23183.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@23191.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@23191.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@23191.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@23191.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@23191.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@23199.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@23207.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@23215.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@23223.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@23231.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@23287.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@23295.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@23295.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@23295.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@23295.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@23295.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@23303.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@23303.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@23303.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@23303.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@23303.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@23311.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@23311.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@23311.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@23311.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@23311.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@23319.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@23319.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@23319.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@23319.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@23319.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@23327.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@23327.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@23327.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@23327.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@23327.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@23335.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@23335.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@23335.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@23335.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@23335.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@23343.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@23351.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@23359.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@23367.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@23375.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@23431.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@23439.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@23439.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@23439.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@23439.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@23439.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@23447.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@23447.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@23447.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@23447.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@23447.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@23455.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@23455.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@23455.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@23455.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@23455.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@23463.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@23463.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@23463.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@23463.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@23463.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@23471.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@23471.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@23471.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@23471.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@23471.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@23479.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@23479.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@23479.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@23479.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@23479.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@23487.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@23495.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@23503.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@23511.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@23519.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@23575.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@23583.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@23583.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@23583.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@23583.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@23583.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@23591.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@23591.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@23591.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@23591.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@23591.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@23599.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@23599.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@23599.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@23599.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@23599.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@23607.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@23607.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@23607.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@23607.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@23607.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@23615.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@23615.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@23615.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@23615.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@23615.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@23623.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@23623.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@23623.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@23623.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@23623.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@23631.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@23639.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@23647.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@23655.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@23663.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@23719.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@23727.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@23727.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@23727.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@23727.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@23727.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@23735.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@23735.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@23735.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@23735.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@23735.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@23743.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@23743.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@23743.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@23743.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@23743.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@23751.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@23751.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@23751.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@23751.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@23751.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@23759.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@23759.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@23759.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@23759.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@23759.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@23767.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@23767.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@23767.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@23767.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@23767.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@23775.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@23783.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@23791.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@23799.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@23807.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_120_io_in; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_120_io_out; // @[package.scala 93:22:@23863.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@23871.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@23871.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@23871.4]
  wire  RetimeWrapper_121_io_in; // @[package.scala 93:22:@23871.4]
  wire  RetimeWrapper_121_io_out; // @[package.scala 93:22:@23871.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@23879.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@23879.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@23879.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@23879.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@23879.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@23887.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@23887.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@23887.4]
  wire  RetimeWrapper_123_io_in; // @[package.scala 93:22:@23887.4]
  wire  RetimeWrapper_123_io_out; // @[package.scala 93:22:@23887.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@23895.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@23895.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@23895.4]
  wire  RetimeWrapper_124_io_in; // @[package.scala 93:22:@23895.4]
  wire  RetimeWrapper_124_io_out; // @[package.scala 93:22:@23895.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@23903.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@23903.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@23903.4]
  wire  RetimeWrapper_125_io_in; // @[package.scala 93:22:@23903.4]
  wire  RetimeWrapper_125_io_out; // @[package.scala 93:22:@23903.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@23911.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@23911.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@23911.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@23911.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@23911.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@23919.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@23927.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_129_io_in; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_129_io_out; // @[package.scala 93:22:@23935.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@23943.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_131_io_in; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_131_io_out; // @[package.scala 93:22:@23951.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_132_io_in; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_132_io_out; // @[package.scala 93:22:@24007.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@24015.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@24015.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@24015.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@24015.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@24015.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@24023.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@24023.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@24023.4]
  wire  RetimeWrapper_134_io_in; // @[package.scala 93:22:@24023.4]
  wire  RetimeWrapper_134_io_out; // @[package.scala 93:22:@24023.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@24031.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@24031.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@24031.4]
  wire  RetimeWrapper_135_io_in; // @[package.scala 93:22:@24031.4]
  wire  RetimeWrapper_135_io_out; // @[package.scala 93:22:@24031.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@24039.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@24039.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@24039.4]
  wire  RetimeWrapper_136_io_in; // @[package.scala 93:22:@24039.4]
  wire  RetimeWrapper_136_io_out; // @[package.scala 93:22:@24039.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@24047.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@24055.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@24055.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@24055.4]
  wire  RetimeWrapper_138_io_in; // @[package.scala 93:22:@24055.4]
  wire  RetimeWrapper_138_io_out; // @[package.scala 93:22:@24055.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_139_io_in; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_139_io_out; // @[package.scala 93:22:@24063.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@24071.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@24079.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_142_io_in; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_142_io_out; // @[package.scala 93:22:@24087.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_143_io_in; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_143_io_out; // @[package.scala 93:22:@24095.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@24151.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@24159.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@24159.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@24159.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@24159.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@24159.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@24167.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@24167.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@24167.4]
  wire  RetimeWrapper_146_io_in; // @[package.scala 93:22:@24167.4]
  wire  RetimeWrapper_146_io_out; // @[package.scala 93:22:@24167.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@24175.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@24175.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@24175.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@24175.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@24175.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@24183.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@24183.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@24183.4]
  wire  RetimeWrapper_148_io_in; // @[package.scala 93:22:@24183.4]
  wire  RetimeWrapper_148_io_out; // @[package.scala 93:22:@24183.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@24191.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@24191.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@24191.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@24191.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@24191.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@24199.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@24199.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@24199.4]
  wire  RetimeWrapper_150_io_in; // @[package.scala 93:22:@24199.4]
  wire  RetimeWrapper_150_io_out; // @[package.scala 93:22:@24199.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@24207.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_152_io_in; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_152_io_out; // @[package.scala 93:22:@24215.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@24223.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_154_io_in; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_154_io_out; // @[package.scala 93:22:@24231.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@24239.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_156_io_in; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_156_io_out; // @[package.scala 93:22:@24295.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@24303.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@24303.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@24303.4]
  wire  RetimeWrapper_157_io_in; // @[package.scala 93:22:@24303.4]
  wire  RetimeWrapper_157_io_out; // @[package.scala 93:22:@24303.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@24311.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@24311.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@24311.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@24311.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@24311.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@24319.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@24319.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@24319.4]
  wire  RetimeWrapper_159_io_in; // @[package.scala 93:22:@24319.4]
  wire  RetimeWrapper_159_io_out; // @[package.scala 93:22:@24319.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@24327.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@24327.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@24327.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@24327.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@24327.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@24335.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@24335.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@24335.4]
  wire  RetimeWrapper_161_io_in; // @[package.scala 93:22:@24335.4]
  wire  RetimeWrapper_161_io_out; // @[package.scala 93:22:@24335.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@24343.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@24343.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@24343.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@24343.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@24343.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_163_io_in; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_163_io_out; // @[package.scala 93:22:@24351.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_164_io_in; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_164_io_out; // @[package.scala 93:22:@24359.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_165_io_in; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_165_io_out; // @[package.scala 93:22:@24367.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_166_io_in; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_166_io_out; // @[package.scala 93:22:@24375.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_167_io_in; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_167_io_out; // @[package.scala 93:22:@24383.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_168_io_in; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_168_io_out; // @[package.scala 93:22:@24439.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@24447.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@24447.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@24447.4]
  wire  RetimeWrapper_169_io_in; // @[package.scala 93:22:@24447.4]
  wire  RetimeWrapper_169_io_out; // @[package.scala 93:22:@24447.4]
  wire  RetimeWrapper_170_clock; // @[package.scala 93:22:@24455.4]
  wire  RetimeWrapper_170_reset; // @[package.scala 93:22:@24455.4]
  wire  RetimeWrapper_170_io_flow; // @[package.scala 93:22:@24455.4]
  wire  RetimeWrapper_170_io_in; // @[package.scala 93:22:@24455.4]
  wire  RetimeWrapper_170_io_out; // @[package.scala 93:22:@24455.4]
  wire  RetimeWrapper_171_clock; // @[package.scala 93:22:@24463.4]
  wire  RetimeWrapper_171_reset; // @[package.scala 93:22:@24463.4]
  wire  RetimeWrapper_171_io_flow; // @[package.scala 93:22:@24463.4]
  wire  RetimeWrapper_171_io_in; // @[package.scala 93:22:@24463.4]
  wire  RetimeWrapper_171_io_out; // @[package.scala 93:22:@24463.4]
  wire  RetimeWrapper_172_clock; // @[package.scala 93:22:@24471.4]
  wire  RetimeWrapper_172_reset; // @[package.scala 93:22:@24471.4]
  wire  RetimeWrapper_172_io_flow; // @[package.scala 93:22:@24471.4]
  wire  RetimeWrapper_172_io_in; // @[package.scala 93:22:@24471.4]
  wire  RetimeWrapper_172_io_out; // @[package.scala 93:22:@24471.4]
  wire  RetimeWrapper_173_clock; // @[package.scala 93:22:@24479.4]
  wire  RetimeWrapper_173_reset; // @[package.scala 93:22:@24479.4]
  wire  RetimeWrapper_173_io_flow; // @[package.scala 93:22:@24479.4]
  wire  RetimeWrapper_173_io_in; // @[package.scala 93:22:@24479.4]
  wire  RetimeWrapper_173_io_out; // @[package.scala 93:22:@24479.4]
  wire  RetimeWrapper_174_clock; // @[package.scala 93:22:@24487.4]
  wire  RetimeWrapper_174_reset; // @[package.scala 93:22:@24487.4]
  wire  RetimeWrapper_174_io_flow; // @[package.scala 93:22:@24487.4]
  wire  RetimeWrapper_174_io_in; // @[package.scala 93:22:@24487.4]
  wire  RetimeWrapper_174_io_out; // @[package.scala 93:22:@24487.4]
  wire  RetimeWrapper_175_clock; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_175_reset; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_175_io_flow; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_175_io_in; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_175_io_out; // @[package.scala 93:22:@24495.4]
  wire  RetimeWrapper_176_clock; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_176_reset; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_176_io_flow; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_176_io_in; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_176_io_out; // @[package.scala 93:22:@24503.4]
  wire  RetimeWrapper_177_clock; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_177_reset; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_177_io_flow; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_177_io_in; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_177_io_out; // @[package.scala 93:22:@24511.4]
  wire  RetimeWrapper_178_clock; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_178_reset; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_178_io_flow; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_178_io_in; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_178_io_out; // @[package.scala 93:22:@24519.4]
  wire  RetimeWrapper_179_clock; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_179_reset; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_179_io_flow; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_179_io_in; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_179_io_out; // @[package.scala 93:22:@24527.4]
  wire  RetimeWrapper_180_clock; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_180_reset; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_180_io_flow; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_180_io_in; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_180_io_out; // @[package.scala 93:22:@24583.4]
  wire  RetimeWrapper_181_clock; // @[package.scala 93:22:@24591.4]
  wire  RetimeWrapper_181_reset; // @[package.scala 93:22:@24591.4]
  wire  RetimeWrapper_181_io_flow; // @[package.scala 93:22:@24591.4]
  wire  RetimeWrapper_181_io_in; // @[package.scala 93:22:@24591.4]
  wire  RetimeWrapper_181_io_out; // @[package.scala 93:22:@24591.4]
  wire  RetimeWrapper_182_clock; // @[package.scala 93:22:@24599.4]
  wire  RetimeWrapper_182_reset; // @[package.scala 93:22:@24599.4]
  wire  RetimeWrapper_182_io_flow; // @[package.scala 93:22:@24599.4]
  wire  RetimeWrapper_182_io_in; // @[package.scala 93:22:@24599.4]
  wire  RetimeWrapper_182_io_out; // @[package.scala 93:22:@24599.4]
  wire  RetimeWrapper_183_clock; // @[package.scala 93:22:@24607.4]
  wire  RetimeWrapper_183_reset; // @[package.scala 93:22:@24607.4]
  wire  RetimeWrapper_183_io_flow; // @[package.scala 93:22:@24607.4]
  wire  RetimeWrapper_183_io_in; // @[package.scala 93:22:@24607.4]
  wire  RetimeWrapper_183_io_out; // @[package.scala 93:22:@24607.4]
  wire  RetimeWrapper_184_clock; // @[package.scala 93:22:@24615.4]
  wire  RetimeWrapper_184_reset; // @[package.scala 93:22:@24615.4]
  wire  RetimeWrapper_184_io_flow; // @[package.scala 93:22:@24615.4]
  wire  RetimeWrapper_184_io_in; // @[package.scala 93:22:@24615.4]
  wire  RetimeWrapper_184_io_out; // @[package.scala 93:22:@24615.4]
  wire  RetimeWrapper_185_clock; // @[package.scala 93:22:@24623.4]
  wire  RetimeWrapper_185_reset; // @[package.scala 93:22:@24623.4]
  wire  RetimeWrapper_185_io_flow; // @[package.scala 93:22:@24623.4]
  wire  RetimeWrapper_185_io_in; // @[package.scala 93:22:@24623.4]
  wire  RetimeWrapper_185_io_out; // @[package.scala 93:22:@24623.4]
  wire  RetimeWrapper_186_clock; // @[package.scala 93:22:@24631.4]
  wire  RetimeWrapper_186_reset; // @[package.scala 93:22:@24631.4]
  wire  RetimeWrapper_186_io_flow; // @[package.scala 93:22:@24631.4]
  wire  RetimeWrapper_186_io_in; // @[package.scala 93:22:@24631.4]
  wire  RetimeWrapper_186_io_out; // @[package.scala 93:22:@24631.4]
  wire  RetimeWrapper_187_clock; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_187_reset; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_187_io_flow; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_187_io_in; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_187_io_out; // @[package.scala 93:22:@24639.4]
  wire  RetimeWrapper_188_clock; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_188_reset; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_188_io_flow; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_188_io_in; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_188_io_out; // @[package.scala 93:22:@24647.4]
  wire  RetimeWrapper_189_clock; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_189_reset; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_189_io_flow; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_189_io_in; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_189_io_out; // @[package.scala 93:22:@24655.4]
  wire  RetimeWrapper_190_clock; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_190_reset; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_190_io_flow; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_190_io_in; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_190_io_out; // @[package.scala 93:22:@24663.4]
  wire  RetimeWrapper_191_clock; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_191_reset; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_191_io_flow; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_191_io_in; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_191_io_out; // @[package.scala 93:22:@24671.4]
  wire  RetimeWrapper_192_clock; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_192_reset; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_192_io_flow; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_192_io_in; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_192_io_out; // @[package.scala 93:22:@24727.4]
  wire  RetimeWrapper_193_clock; // @[package.scala 93:22:@24735.4]
  wire  RetimeWrapper_193_reset; // @[package.scala 93:22:@24735.4]
  wire  RetimeWrapper_193_io_flow; // @[package.scala 93:22:@24735.4]
  wire  RetimeWrapper_193_io_in; // @[package.scala 93:22:@24735.4]
  wire  RetimeWrapper_193_io_out; // @[package.scala 93:22:@24735.4]
  wire  RetimeWrapper_194_clock; // @[package.scala 93:22:@24743.4]
  wire  RetimeWrapper_194_reset; // @[package.scala 93:22:@24743.4]
  wire  RetimeWrapper_194_io_flow; // @[package.scala 93:22:@24743.4]
  wire  RetimeWrapper_194_io_in; // @[package.scala 93:22:@24743.4]
  wire  RetimeWrapper_194_io_out; // @[package.scala 93:22:@24743.4]
  wire  RetimeWrapper_195_clock; // @[package.scala 93:22:@24751.4]
  wire  RetimeWrapper_195_reset; // @[package.scala 93:22:@24751.4]
  wire  RetimeWrapper_195_io_flow; // @[package.scala 93:22:@24751.4]
  wire  RetimeWrapper_195_io_in; // @[package.scala 93:22:@24751.4]
  wire  RetimeWrapper_195_io_out; // @[package.scala 93:22:@24751.4]
  wire  RetimeWrapper_196_clock; // @[package.scala 93:22:@24759.4]
  wire  RetimeWrapper_196_reset; // @[package.scala 93:22:@24759.4]
  wire  RetimeWrapper_196_io_flow; // @[package.scala 93:22:@24759.4]
  wire  RetimeWrapper_196_io_in; // @[package.scala 93:22:@24759.4]
  wire  RetimeWrapper_196_io_out; // @[package.scala 93:22:@24759.4]
  wire  RetimeWrapper_197_clock; // @[package.scala 93:22:@24767.4]
  wire  RetimeWrapper_197_reset; // @[package.scala 93:22:@24767.4]
  wire  RetimeWrapper_197_io_flow; // @[package.scala 93:22:@24767.4]
  wire  RetimeWrapper_197_io_in; // @[package.scala 93:22:@24767.4]
  wire  RetimeWrapper_197_io_out; // @[package.scala 93:22:@24767.4]
  wire  RetimeWrapper_198_clock; // @[package.scala 93:22:@24775.4]
  wire  RetimeWrapper_198_reset; // @[package.scala 93:22:@24775.4]
  wire  RetimeWrapper_198_io_flow; // @[package.scala 93:22:@24775.4]
  wire  RetimeWrapper_198_io_in; // @[package.scala 93:22:@24775.4]
  wire  RetimeWrapper_198_io_out; // @[package.scala 93:22:@24775.4]
  wire  RetimeWrapper_199_clock; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_199_reset; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_199_io_flow; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_199_io_in; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_199_io_out; // @[package.scala 93:22:@24783.4]
  wire  RetimeWrapper_200_clock; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_200_reset; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_200_io_flow; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_200_io_in; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_200_io_out; // @[package.scala 93:22:@24791.4]
  wire  RetimeWrapper_201_clock; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_201_reset; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_201_io_flow; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_201_io_in; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_201_io_out; // @[package.scala 93:22:@24799.4]
  wire  RetimeWrapper_202_clock; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_202_reset; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_202_io_flow; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_202_io_in; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_202_io_out; // @[package.scala 93:22:@24807.4]
  wire  RetimeWrapper_203_clock; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_203_reset; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_203_io_flow; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_203_io_in; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_203_io_out; // @[package.scala 93:22:@24815.4]
  wire  RetimeWrapper_204_clock; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_204_reset; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_204_io_flow; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_204_io_in; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_204_io_out; // @[package.scala 93:22:@24871.4]
  wire  RetimeWrapper_205_clock; // @[package.scala 93:22:@24879.4]
  wire  RetimeWrapper_205_reset; // @[package.scala 93:22:@24879.4]
  wire  RetimeWrapper_205_io_flow; // @[package.scala 93:22:@24879.4]
  wire  RetimeWrapper_205_io_in; // @[package.scala 93:22:@24879.4]
  wire  RetimeWrapper_205_io_out; // @[package.scala 93:22:@24879.4]
  wire  RetimeWrapper_206_clock; // @[package.scala 93:22:@24887.4]
  wire  RetimeWrapper_206_reset; // @[package.scala 93:22:@24887.4]
  wire  RetimeWrapper_206_io_flow; // @[package.scala 93:22:@24887.4]
  wire  RetimeWrapper_206_io_in; // @[package.scala 93:22:@24887.4]
  wire  RetimeWrapper_206_io_out; // @[package.scala 93:22:@24887.4]
  wire  RetimeWrapper_207_clock; // @[package.scala 93:22:@24895.4]
  wire  RetimeWrapper_207_reset; // @[package.scala 93:22:@24895.4]
  wire  RetimeWrapper_207_io_flow; // @[package.scala 93:22:@24895.4]
  wire  RetimeWrapper_207_io_in; // @[package.scala 93:22:@24895.4]
  wire  RetimeWrapper_207_io_out; // @[package.scala 93:22:@24895.4]
  wire  RetimeWrapper_208_clock; // @[package.scala 93:22:@24903.4]
  wire  RetimeWrapper_208_reset; // @[package.scala 93:22:@24903.4]
  wire  RetimeWrapper_208_io_flow; // @[package.scala 93:22:@24903.4]
  wire  RetimeWrapper_208_io_in; // @[package.scala 93:22:@24903.4]
  wire  RetimeWrapper_208_io_out; // @[package.scala 93:22:@24903.4]
  wire  RetimeWrapper_209_clock; // @[package.scala 93:22:@24911.4]
  wire  RetimeWrapper_209_reset; // @[package.scala 93:22:@24911.4]
  wire  RetimeWrapper_209_io_flow; // @[package.scala 93:22:@24911.4]
  wire  RetimeWrapper_209_io_in; // @[package.scala 93:22:@24911.4]
  wire  RetimeWrapper_209_io_out; // @[package.scala 93:22:@24911.4]
  wire  RetimeWrapper_210_clock; // @[package.scala 93:22:@24919.4]
  wire  RetimeWrapper_210_reset; // @[package.scala 93:22:@24919.4]
  wire  RetimeWrapper_210_io_flow; // @[package.scala 93:22:@24919.4]
  wire  RetimeWrapper_210_io_in; // @[package.scala 93:22:@24919.4]
  wire  RetimeWrapper_210_io_out; // @[package.scala 93:22:@24919.4]
  wire  RetimeWrapper_211_clock; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_211_reset; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_211_io_flow; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_211_io_in; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_211_io_out; // @[package.scala 93:22:@24927.4]
  wire  RetimeWrapper_212_clock; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_212_reset; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_212_io_flow; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_212_io_in; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_212_io_out; // @[package.scala 93:22:@24935.4]
  wire  RetimeWrapper_213_clock; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_213_reset; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_213_io_flow; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_213_io_in; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_213_io_out; // @[package.scala 93:22:@24943.4]
  wire  RetimeWrapper_214_clock; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_214_reset; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_214_io_flow; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_214_io_in; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_214_io_out; // @[package.scala 93:22:@24951.4]
  wire  RetimeWrapper_215_clock; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_215_reset; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_215_io_flow; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_215_io_in; // @[package.scala 93:22:@24959.4]
  wire  RetimeWrapper_215_io_out; // @[package.scala 93:22:@24959.4]
  wire  _T_700; // @[MemPrimitives.scala 82:210:@19794.4]
  wire  _T_702; // @[MemPrimitives.scala 82:210:@19795.4]
  wire  _T_703; // @[MemPrimitives.scala 82:228:@19796.4]
  wire  _T_704; // @[MemPrimitives.scala 83:102:@19797.4]
  wire  _T_706; // @[MemPrimitives.scala 82:210:@19798.4]
  wire  _T_708; // @[MemPrimitives.scala 82:210:@19799.4]
  wire  _T_709; // @[MemPrimitives.scala 82:228:@19800.4]
  wire  _T_710; // @[MemPrimitives.scala 83:102:@19801.4]
  wire [41:0] _T_712; // @[Cat.scala 30:58:@19803.4]
  wire [41:0] _T_714; // @[Cat.scala 30:58:@19805.4]
  wire [41:0] _T_715; // @[Mux.scala 31:69:@19806.4]
  wire  _T_720; // @[MemPrimitives.scala 82:210:@19813.4]
  wire  _T_722; // @[MemPrimitives.scala 82:210:@19814.4]
  wire  _T_723; // @[MemPrimitives.scala 82:228:@19815.4]
  wire  _T_724; // @[MemPrimitives.scala 83:102:@19816.4]
  wire  _T_726; // @[MemPrimitives.scala 82:210:@19817.4]
  wire  _T_728; // @[MemPrimitives.scala 82:210:@19818.4]
  wire  _T_729; // @[MemPrimitives.scala 82:228:@19819.4]
  wire  _T_730; // @[MemPrimitives.scala 83:102:@19820.4]
  wire [41:0] _T_732; // @[Cat.scala 30:58:@19822.4]
  wire [41:0] _T_734; // @[Cat.scala 30:58:@19824.4]
  wire [41:0] _T_735; // @[Mux.scala 31:69:@19825.4]
  wire  _T_742; // @[MemPrimitives.scala 82:210:@19833.4]
  wire  _T_743; // @[MemPrimitives.scala 82:228:@19834.4]
  wire  _T_744; // @[MemPrimitives.scala 83:102:@19835.4]
  wire  _T_748; // @[MemPrimitives.scala 82:210:@19837.4]
  wire  _T_749; // @[MemPrimitives.scala 82:228:@19838.4]
  wire  _T_750; // @[MemPrimitives.scala 83:102:@19839.4]
  wire [41:0] _T_752; // @[Cat.scala 30:58:@19841.4]
  wire [41:0] _T_754; // @[Cat.scala 30:58:@19843.4]
  wire [41:0] _T_755; // @[Mux.scala 31:69:@19844.4]
  wire  _T_762; // @[MemPrimitives.scala 82:210:@19852.4]
  wire  _T_763; // @[MemPrimitives.scala 82:228:@19853.4]
  wire  _T_764; // @[MemPrimitives.scala 83:102:@19854.4]
  wire  _T_768; // @[MemPrimitives.scala 82:210:@19856.4]
  wire  _T_769; // @[MemPrimitives.scala 82:228:@19857.4]
  wire  _T_770; // @[MemPrimitives.scala 83:102:@19858.4]
  wire [41:0] _T_772; // @[Cat.scala 30:58:@19860.4]
  wire [41:0] _T_774; // @[Cat.scala 30:58:@19862.4]
  wire [41:0] _T_775; // @[Mux.scala 31:69:@19863.4]
  wire  _T_782; // @[MemPrimitives.scala 82:210:@19871.4]
  wire  _T_783; // @[MemPrimitives.scala 82:228:@19872.4]
  wire  _T_784; // @[MemPrimitives.scala 83:102:@19873.4]
  wire  _T_788; // @[MemPrimitives.scala 82:210:@19875.4]
  wire  _T_789; // @[MemPrimitives.scala 82:228:@19876.4]
  wire  _T_790; // @[MemPrimitives.scala 83:102:@19877.4]
  wire [41:0] _T_792; // @[Cat.scala 30:58:@19879.4]
  wire [41:0] _T_794; // @[Cat.scala 30:58:@19881.4]
  wire [41:0] _T_795; // @[Mux.scala 31:69:@19882.4]
  wire  _T_802; // @[MemPrimitives.scala 82:210:@19890.4]
  wire  _T_803; // @[MemPrimitives.scala 82:228:@19891.4]
  wire  _T_804; // @[MemPrimitives.scala 83:102:@19892.4]
  wire  _T_808; // @[MemPrimitives.scala 82:210:@19894.4]
  wire  _T_809; // @[MemPrimitives.scala 82:228:@19895.4]
  wire  _T_810; // @[MemPrimitives.scala 83:102:@19896.4]
  wire [41:0] _T_812; // @[Cat.scala 30:58:@19898.4]
  wire [41:0] _T_814; // @[Cat.scala 30:58:@19900.4]
  wire [41:0] _T_815; // @[Mux.scala 31:69:@19901.4]
  wire  _T_820; // @[MemPrimitives.scala 82:210:@19908.4]
  wire  _T_823; // @[MemPrimitives.scala 82:228:@19910.4]
  wire  _T_824; // @[MemPrimitives.scala 83:102:@19911.4]
  wire  _T_826; // @[MemPrimitives.scala 82:210:@19912.4]
  wire  _T_829; // @[MemPrimitives.scala 82:228:@19914.4]
  wire  _T_830; // @[MemPrimitives.scala 83:102:@19915.4]
  wire [41:0] _T_832; // @[Cat.scala 30:58:@19917.4]
  wire [41:0] _T_834; // @[Cat.scala 30:58:@19919.4]
  wire [41:0] _T_835; // @[Mux.scala 31:69:@19920.4]
  wire  _T_840; // @[MemPrimitives.scala 82:210:@19927.4]
  wire  _T_843; // @[MemPrimitives.scala 82:228:@19929.4]
  wire  _T_844; // @[MemPrimitives.scala 83:102:@19930.4]
  wire  _T_846; // @[MemPrimitives.scala 82:210:@19931.4]
  wire  _T_849; // @[MemPrimitives.scala 82:228:@19933.4]
  wire  _T_850; // @[MemPrimitives.scala 83:102:@19934.4]
  wire [41:0] _T_852; // @[Cat.scala 30:58:@19936.4]
  wire [41:0] _T_854; // @[Cat.scala 30:58:@19938.4]
  wire [41:0] _T_855; // @[Mux.scala 31:69:@19939.4]
  wire  _T_863; // @[MemPrimitives.scala 82:228:@19948.4]
  wire  _T_864; // @[MemPrimitives.scala 83:102:@19949.4]
  wire  _T_869; // @[MemPrimitives.scala 82:228:@19952.4]
  wire  _T_870; // @[MemPrimitives.scala 83:102:@19953.4]
  wire [41:0] _T_872; // @[Cat.scala 30:58:@19955.4]
  wire [41:0] _T_874; // @[Cat.scala 30:58:@19957.4]
  wire [41:0] _T_875; // @[Mux.scala 31:69:@19958.4]
  wire  _T_883; // @[MemPrimitives.scala 82:228:@19967.4]
  wire  _T_884; // @[MemPrimitives.scala 83:102:@19968.4]
  wire  _T_889; // @[MemPrimitives.scala 82:228:@19971.4]
  wire  _T_890; // @[MemPrimitives.scala 83:102:@19972.4]
  wire [41:0] _T_892; // @[Cat.scala 30:58:@19974.4]
  wire [41:0] _T_894; // @[Cat.scala 30:58:@19976.4]
  wire [41:0] _T_895; // @[Mux.scala 31:69:@19977.4]
  wire  _T_903; // @[MemPrimitives.scala 82:228:@19986.4]
  wire  _T_904; // @[MemPrimitives.scala 83:102:@19987.4]
  wire  _T_909; // @[MemPrimitives.scala 82:228:@19990.4]
  wire  _T_910; // @[MemPrimitives.scala 83:102:@19991.4]
  wire [41:0] _T_912; // @[Cat.scala 30:58:@19993.4]
  wire [41:0] _T_914; // @[Cat.scala 30:58:@19995.4]
  wire [41:0] _T_915; // @[Mux.scala 31:69:@19996.4]
  wire  _T_923; // @[MemPrimitives.scala 82:228:@20005.4]
  wire  _T_924; // @[MemPrimitives.scala 83:102:@20006.4]
  wire  _T_929; // @[MemPrimitives.scala 82:228:@20009.4]
  wire  _T_930; // @[MemPrimitives.scala 83:102:@20010.4]
  wire [41:0] _T_932; // @[Cat.scala 30:58:@20012.4]
  wire [41:0] _T_934; // @[Cat.scala 30:58:@20014.4]
  wire [41:0] _T_935; // @[Mux.scala 31:69:@20015.4]
  wire  _T_940; // @[MemPrimitives.scala 82:210:@20022.4]
  wire  _T_943; // @[MemPrimitives.scala 82:228:@20024.4]
  wire  _T_944; // @[MemPrimitives.scala 83:102:@20025.4]
  wire  _T_946; // @[MemPrimitives.scala 82:210:@20026.4]
  wire  _T_949; // @[MemPrimitives.scala 82:228:@20028.4]
  wire  _T_950; // @[MemPrimitives.scala 83:102:@20029.4]
  wire [41:0] _T_952; // @[Cat.scala 30:58:@20031.4]
  wire [41:0] _T_954; // @[Cat.scala 30:58:@20033.4]
  wire [41:0] _T_955; // @[Mux.scala 31:69:@20034.4]
  wire  _T_960; // @[MemPrimitives.scala 82:210:@20041.4]
  wire  _T_963; // @[MemPrimitives.scala 82:228:@20043.4]
  wire  _T_964; // @[MemPrimitives.scala 83:102:@20044.4]
  wire  _T_966; // @[MemPrimitives.scala 82:210:@20045.4]
  wire  _T_969; // @[MemPrimitives.scala 82:228:@20047.4]
  wire  _T_970; // @[MemPrimitives.scala 83:102:@20048.4]
  wire [41:0] _T_972; // @[Cat.scala 30:58:@20050.4]
  wire [41:0] _T_974; // @[Cat.scala 30:58:@20052.4]
  wire [41:0] _T_975; // @[Mux.scala 31:69:@20053.4]
  wire  _T_983; // @[MemPrimitives.scala 82:228:@20062.4]
  wire  _T_984; // @[MemPrimitives.scala 83:102:@20063.4]
  wire  _T_989; // @[MemPrimitives.scala 82:228:@20066.4]
  wire  _T_990; // @[MemPrimitives.scala 83:102:@20067.4]
  wire [41:0] _T_992; // @[Cat.scala 30:58:@20069.4]
  wire [41:0] _T_994; // @[Cat.scala 30:58:@20071.4]
  wire [41:0] _T_995; // @[Mux.scala 31:69:@20072.4]
  wire  _T_1003; // @[MemPrimitives.scala 82:228:@20081.4]
  wire  _T_1004; // @[MemPrimitives.scala 83:102:@20082.4]
  wire  _T_1009; // @[MemPrimitives.scala 82:228:@20085.4]
  wire  _T_1010; // @[MemPrimitives.scala 83:102:@20086.4]
  wire [41:0] _T_1012; // @[Cat.scala 30:58:@20088.4]
  wire [41:0] _T_1014; // @[Cat.scala 30:58:@20090.4]
  wire [41:0] _T_1015; // @[Mux.scala 31:69:@20091.4]
  wire  _T_1023; // @[MemPrimitives.scala 82:228:@20100.4]
  wire  _T_1024; // @[MemPrimitives.scala 83:102:@20101.4]
  wire  _T_1029; // @[MemPrimitives.scala 82:228:@20104.4]
  wire  _T_1030; // @[MemPrimitives.scala 83:102:@20105.4]
  wire [41:0] _T_1032; // @[Cat.scala 30:58:@20107.4]
  wire [41:0] _T_1034; // @[Cat.scala 30:58:@20109.4]
  wire [41:0] _T_1035; // @[Mux.scala 31:69:@20110.4]
  wire  _T_1043; // @[MemPrimitives.scala 82:228:@20119.4]
  wire  _T_1044; // @[MemPrimitives.scala 83:102:@20120.4]
  wire  _T_1049; // @[MemPrimitives.scala 82:228:@20123.4]
  wire  _T_1050; // @[MemPrimitives.scala 83:102:@20124.4]
  wire [41:0] _T_1052; // @[Cat.scala 30:58:@20126.4]
  wire [41:0] _T_1054; // @[Cat.scala 30:58:@20128.4]
  wire [41:0] _T_1055; // @[Mux.scala 31:69:@20129.4]
  wire  _T_1060; // @[MemPrimitives.scala 82:210:@20136.4]
  wire  _T_1063; // @[MemPrimitives.scala 82:228:@20138.4]
  wire  _T_1064; // @[MemPrimitives.scala 83:102:@20139.4]
  wire  _T_1066; // @[MemPrimitives.scala 82:210:@20140.4]
  wire  _T_1069; // @[MemPrimitives.scala 82:228:@20142.4]
  wire  _T_1070; // @[MemPrimitives.scala 83:102:@20143.4]
  wire [41:0] _T_1072; // @[Cat.scala 30:58:@20145.4]
  wire [41:0] _T_1074; // @[Cat.scala 30:58:@20147.4]
  wire [41:0] _T_1075; // @[Mux.scala 31:69:@20148.4]
  wire  _T_1080; // @[MemPrimitives.scala 82:210:@20155.4]
  wire  _T_1083; // @[MemPrimitives.scala 82:228:@20157.4]
  wire  _T_1084; // @[MemPrimitives.scala 83:102:@20158.4]
  wire  _T_1086; // @[MemPrimitives.scala 82:210:@20159.4]
  wire  _T_1089; // @[MemPrimitives.scala 82:228:@20161.4]
  wire  _T_1090; // @[MemPrimitives.scala 83:102:@20162.4]
  wire [41:0] _T_1092; // @[Cat.scala 30:58:@20164.4]
  wire [41:0] _T_1094; // @[Cat.scala 30:58:@20166.4]
  wire [41:0] _T_1095; // @[Mux.scala 31:69:@20167.4]
  wire  _T_1103; // @[MemPrimitives.scala 82:228:@20176.4]
  wire  _T_1104; // @[MemPrimitives.scala 83:102:@20177.4]
  wire  _T_1109; // @[MemPrimitives.scala 82:228:@20180.4]
  wire  _T_1110; // @[MemPrimitives.scala 83:102:@20181.4]
  wire [41:0] _T_1112; // @[Cat.scala 30:58:@20183.4]
  wire [41:0] _T_1114; // @[Cat.scala 30:58:@20185.4]
  wire [41:0] _T_1115; // @[Mux.scala 31:69:@20186.4]
  wire  _T_1123; // @[MemPrimitives.scala 82:228:@20195.4]
  wire  _T_1124; // @[MemPrimitives.scala 83:102:@20196.4]
  wire  _T_1129; // @[MemPrimitives.scala 82:228:@20199.4]
  wire  _T_1130; // @[MemPrimitives.scala 83:102:@20200.4]
  wire [41:0] _T_1132; // @[Cat.scala 30:58:@20202.4]
  wire [41:0] _T_1134; // @[Cat.scala 30:58:@20204.4]
  wire [41:0] _T_1135; // @[Mux.scala 31:69:@20205.4]
  wire  _T_1143; // @[MemPrimitives.scala 82:228:@20214.4]
  wire  _T_1144; // @[MemPrimitives.scala 83:102:@20215.4]
  wire  _T_1149; // @[MemPrimitives.scala 82:228:@20218.4]
  wire  _T_1150; // @[MemPrimitives.scala 83:102:@20219.4]
  wire [41:0] _T_1152; // @[Cat.scala 30:58:@20221.4]
  wire [41:0] _T_1154; // @[Cat.scala 30:58:@20223.4]
  wire [41:0] _T_1155; // @[Mux.scala 31:69:@20224.4]
  wire  _T_1163; // @[MemPrimitives.scala 82:228:@20233.4]
  wire  _T_1164; // @[MemPrimitives.scala 83:102:@20234.4]
  wire  _T_1169; // @[MemPrimitives.scala 82:228:@20237.4]
  wire  _T_1170; // @[MemPrimitives.scala 83:102:@20238.4]
  wire [41:0] _T_1172; // @[Cat.scala 30:58:@20240.4]
  wire [41:0] _T_1174; // @[Cat.scala 30:58:@20242.4]
  wire [41:0] _T_1175; // @[Mux.scala 31:69:@20243.4]
  wire  _T_1180; // @[MemPrimitives.scala 110:210:@20250.4]
  wire  _T_1182; // @[MemPrimitives.scala 110:210:@20251.4]
  wire  _T_1183; // @[MemPrimitives.scala 110:228:@20252.4]
  wire  _T_1186; // @[MemPrimitives.scala 110:210:@20254.4]
  wire  _T_1188; // @[MemPrimitives.scala 110:210:@20255.4]
  wire  _T_1189; // @[MemPrimitives.scala 110:228:@20256.4]
  wire  _T_1192; // @[MemPrimitives.scala 110:210:@20258.4]
  wire  _T_1194; // @[MemPrimitives.scala 110:210:@20259.4]
  wire  _T_1195; // @[MemPrimitives.scala 110:228:@20260.4]
  wire  _T_1198; // @[MemPrimitives.scala 110:210:@20262.4]
  wire  _T_1200; // @[MemPrimitives.scala 110:210:@20263.4]
  wire  _T_1201; // @[MemPrimitives.scala 110:228:@20264.4]
  wire  _T_1204; // @[MemPrimitives.scala 110:210:@20266.4]
  wire  _T_1206; // @[MemPrimitives.scala 110:210:@20267.4]
  wire  _T_1207; // @[MemPrimitives.scala 110:228:@20268.4]
  wire  _T_1210; // @[MemPrimitives.scala 110:210:@20270.4]
  wire  _T_1212; // @[MemPrimitives.scala 110:210:@20271.4]
  wire  _T_1213; // @[MemPrimitives.scala 110:228:@20272.4]
  wire  _T_1216; // @[MemPrimitives.scala 110:210:@20274.4]
  wire  _T_1218; // @[MemPrimitives.scala 110:210:@20275.4]
  wire  _T_1219; // @[MemPrimitives.scala 110:228:@20276.4]
  wire  _T_1222; // @[MemPrimitives.scala 110:210:@20278.4]
  wire  _T_1224; // @[MemPrimitives.scala 110:210:@20279.4]
  wire  _T_1225; // @[MemPrimitives.scala 110:228:@20280.4]
  wire  _T_1228; // @[MemPrimitives.scala 110:210:@20282.4]
  wire  _T_1230; // @[MemPrimitives.scala 110:210:@20283.4]
  wire  _T_1231; // @[MemPrimitives.scala 110:228:@20284.4]
  wire  _T_1233; // @[MemPrimitives.scala 126:35:@20298.4]
  wire  _T_1234; // @[MemPrimitives.scala 126:35:@20299.4]
  wire  _T_1235; // @[MemPrimitives.scala 126:35:@20300.4]
  wire  _T_1236; // @[MemPrimitives.scala 126:35:@20301.4]
  wire  _T_1237; // @[MemPrimitives.scala 126:35:@20302.4]
  wire  _T_1238; // @[MemPrimitives.scala 126:35:@20303.4]
  wire  _T_1239; // @[MemPrimitives.scala 126:35:@20304.4]
  wire  _T_1240; // @[MemPrimitives.scala 126:35:@20305.4]
  wire  _T_1241; // @[MemPrimitives.scala 126:35:@20306.4]
  wire [10:0] _T_1243; // @[Cat.scala 30:58:@20308.4]
  wire [10:0] _T_1245; // @[Cat.scala 30:58:@20310.4]
  wire [10:0] _T_1247; // @[Cat.scala 30:58:@20312.4]
  wire [10:0] _T_1249; // @[Cat.scala 30:58:@20314.4]
  wire [10:0] _T_1251; // @[Cat.scala 30:58:@20316.4]
  wire [10:0] _T_1253; // @[Cat.scala 30:58:@20318.4]
  wire [10:0] _T_1255; // @[Cat.scala 30:58:@20320.4]
  wire [10:0] _T_1257; // @[Cat.scala 30:58:@20322.4]
  wire [10:0] _T_1259; // @[Cat.scala 30:58:@20324.4]
  wire [10:0] _T_1260; // @[Mux.scala 31:69:@20325.4]
  wire [10:0] _T_1261; // @[Mux.scala 31:69:@20326.4]
  wire [10:0] _T_1262; // @[Mux.scala 31:69:@20327.4]
  wire [10:0] _T_1263; // @[Mux.scala 31:69:@20328.4]
  wire [10:0] _T_1264; // @[Mux.scala 31:69:@20329.4]
  wire [10:0] _T_1265; // @[Mux.scala 31:69:@20330.4]
  wire [10:0] _T_1266; // @[Mux.scala 31:69:@20331.4]
  wire [10:0] _T_1267; // @[Mux.scala 31:69:@20332.4]
  wire  _T_1272; // @[MemPrimitives.scala 110:210:@20339.4]
  wire  _T_1274; // @[MemPrimitives.scala 110:210:@20340.4]
  wire  _T_1275; // @[MemPrimitives.scala 110:228:@20341.4]
  wire  _T_1278; // @[MemPrimitives.scala 110:210:@20343.4]
  wire  _T_1280; // @[MemPrimitives.scala 110:210:@20344.4]
  wire  _T_1281; // @[MemPrimitives.scala 110:228:@20345.4]
  wire  _T_1284; // @[MemPrimitives.scala 110:210:@20347.4]
  wire  _T_1286; // @[MemPrimitives.scala 110:210:@20348.4]
  wire  _T_1287; // @[MemPrimitives.scala 110:228:@20349.4]
  wire  _T_1290; // @[MemPrimitives.scala 110:210:@20351.4]
  wire  _T_1292; // @[MemPrimitives.scala 110:210:@20352.4]
  wire  _T_1293; // @[MemPrimitives.scala 110:228:@20353.4]
  wire  _T_1296; // @[MemPrimitives.scala 110:210:@20355.4]
  wire  _T_1298; // @[MemPrimitives.scala 110:210:@20356.4]
  wire  _T_1299; // @[MemPrimitives.scala 110:228:@20357.4]
  wire  _T_1302; // @[MemPrimitives.scala 110:210:@20359.4]
  wire  _T_1304; // @[MemPrimitives.scala 110:210:@20360.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@20361.4]
  wire  _T_1308; // @[MemPrimitives.scala 110:210:@20363.4]
  wire  _T_1310; // @[MemPrimitives.scala 110:210:@20364.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@20365.4]
  wire  _T_1314; // @[MemPrimitives.scala 110:210:@20367.4]
  wire  _T_1316; // @[MemPrimitives.scala 110:210:@20368.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@20369.4]
  wire  _T_1320; // @[MemPrimitives.scala 110:210:@20371.4]
  wire  _T_1322; // @[MemPrimitives.scala 110:210:@20372.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@20373.4]
  wire  _T_1325; // @[MemPrimitives.scala 126:35:@20387.4]
  wire  _T_1326; // @[MemPrimitives.scala 126:35:@20388.4]
  wire  _T_1327; // @[MemPrimitives.scala 126:35:@20389.4]
  wire  _T_1328; // @[MemPrimitives.scala 126:35:@20390.4]
  wire  _T_1329; // @[MemPrimitives.scala 126:35:@20391.4]
  wire  _T_1330; // @[MemPrimitives.scala 126:35:@20392.4]
  wire  _T_1331; // @[MemPrimitives.scala 126:35:@20393.4]
  wire  _T_1332; // @[MemPrimitives.scala 126:35:@20394.4]
  wire  _T_1333; // @[MemPrimitives.scala 126:35:@20395.4]
  wire [10:0] _T_1335; // @[Cat.scala 30:58:@20397.4]
  wire [10:0] _T_1337; // @[Cat.scala 30:58:@20399.4]
  wire [10:0] _T_1339; // @[Cat.scala 30:58:@20401.4]
  wire [10:0] _T_1341; // @[Cat.scala 30:58:@20403.4]
  wire [10:0] _T_1343; // @[Cat.scala 30:58:@20405.4]
  wire [10:0] _T_1345; // @[Cat.scala 30:58:@20407.4]
  wire [10:0] _T_1347; // @[Cat.scala 30:58:@20409.4]
  wire [10:0] _T_1349; // @[Cat.scala 30:58:@20411.4]
  wire [10:0] _T_1351; // @[Cat.scala 30:58:@20413.4]
  wire [10:0] _T_1352; // @[Mux.scala 31:69:@20414.4]
  wire [10:0] _T_1353; // @[Mux.scala 31:69:@20415.4]
  wire [10:0] _T_1354; // @[Mux.scala 31:69:@20416.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@20417.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@20418.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@20419.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@20420.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@20421.4]
  wire  _T_1366; // @[MemPrimitives.scala 110:210:@20429.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@20430.4]
  wire  _T_1372; // @[MemPrimitives.scala 110:210:@20433.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@20434.4]
  wire  _T_1378; // @[MemPrimitives.scala 110:210:@20437.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@20438.4]
  wire  _T_1384; // @[MemPrimitives.scala 110:210:@20441.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@20442.4]
  wire  _T_1390; // @[MemPrimitives.scala 110:210:@20445.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@20446.4]
  wire  _T_1396; // @[MemPrimitives.scala 110:210:@20449.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@20450.4]
  wire  _T_1402; // @[MemPrimitives.scala 110:210:@20453.4]
  wire  _T_1403; // @[MemPrimitives.scala 110:228:@20454.4]
  wire  _T_1408; // @[MemPrimitives.scala 110:210:@20457.4]
  wire  _T_1409; // @[MemPrimitives.scala 110:228:@20458.4]
  wire  _T_1414; // @[MemPrimitives.scala 110:210:@20461.4]
  wire  _T_1415; // @[MemPrimitives.scala 110:228:@20462.4]
  wire  _T_1417; // @[MemPrimitives.scala 126:35:@20476.4]
  wire  _T_1418; // @[MemPrimitives.scala 126:35:@20477.4]
  wire  _T_1419; // @[MemPrimitives.scala 126:35:@20478.4]
  wire  _T_1420; // @[MemPrimitives.scala 126:35:@20479.4]
  wire  _T_1421; // @[MemPrimitives.scala 126:35:@20480.4]
  wire  _T_1422; // @[MemPrimitives.scala 126:35:@20481.4]
  wire  _T_1423; // @[MemPrimitives.scala 126:35:@20482.4]
  wire  _T_1424; // @[MemPrimitives.scala 126:35:@20483.4]
  wire  _T_1425; // @[MemPrimitives.scala 126:35:@20484.4]
  wire [10:0] _T_1427; // @[Cat.scala 30:58:@20486.4]
  wire [10:0] _T_1429; // @[Cat.scala 30:58:@20488.4]
  wire [10:0] _T_1431; // @[Cat.scala 30:58:@20490.4]
  wire [10:0] _T_1433; // @[Cat.scala 30:58:@20492.4]
  wire [10:0] _T_1435; // @[Cat.scala 30:58:@20494.4]
  wire [10:0] _T_1437; // @[Cat.scala 30:58:@20496.4]
  wire [10:0] _T_1439; // @[Cat.scala 30:58:@20498.4]
  wire [10:0] _T_1441; // @[Cat.scala 30:58:@20500.4]
  wire [10:0] _T_1443; // @[Cat.scala 30:58:@20502.4]
  wire [10:0] _T_1444; // @[Mux.scala 31:69:@20503.4]
  wire [10:0] _T_1445; // @[Mux.scala 31:69:@20504.4]
  wire [10:0] _T_1446; // @[Mux.scala 31:69:@20505.4]
  wire [10:0] _T_1447; // @[Mux.scala 31:69:@20506.4]
  wire [10:0] _T_1448; // @[Mux.scala 31:69:@20507.4]
  wire [10:0] _T_1449; // @[Mux.scala 31:69:@20508.4]
  wire [10:0] _T_1450; // @[Mux.scala 31:69:@20509.4]
  wire [10:0] _T_1451; // @[Mux.scala 31:69:@20510.4]
  wire  _T_1458; // @[MemPrimitives.scala 110:210:@20518.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@20519.4]
  wire  _T_1464; // @[MemPrimitives.scala 110:210:@20522.4]
  wire  _T_1465; // @[MemPrimitives.scala 110:228:@20523.4]
  wire  _T_1470; // @[MemPrimitives.scala 110:210:@20526.4]
  wire  _T_1471; // @[MemPrimitives.scala 110:228:@20527.4]
  wire  _T_1476; // @[MemPrimitives.scala 110:210:@20530.4]
  wire  _T_1477; // @[MemPrimitives.scala 110:228:@20531.4]
  wire  _T_1482; // @[MemPrimitives.scala 110:210:@20534.4]
  wire  _T_1483; // @[MemPrimitives.scala 110:228:@20535.4]
  wire  _T_1488; // @[MemPrimitives.scala 110:210:@20538.4]
  wire  _T_1489; // @[MemPrimitives.scala 110:228:@20539.4]
  wire  _T_1494; // @[MemPrimitives.scala 110:210:@20542.4]
  wire  _T_1495; // @[MemPrimitives.scala 110:228:@20543.4]
  wire  _T_1500; // @[MemPrimitives.scala 110:210:@20546.4]
  wire  _T_1501; // @[MemPrimitives.scala 110:228:@20547.4]
  wire  _T_1506; // @[MemPrimitives.scala 110:210:@20550.4]
  wire  _T_1507; // @[MemPrimitives.scala 110:228:@20551.4]
  wire  _T_1509; // @[MemPrimitives.scala 126:35:@20565.4]
  wire  _T_1510; // @[MemPrimitives.scala 126:35:@20566.4]
  wire  _T_1511; // @[MemPrimitives.scala 126:35:@20567.4]
  wire  _T_1512; // @[MemPrimitives.scala 126:35:@20568.4]
  wire  _T_1513; // @[MemPrimitives.scala 126:35:@20569.4]
  wire  _T_1514; // @[MemPrimitives.scala 126:35:@20570.4]
  wire  _T_1515; // @[MemPrimitives.scala 126:35:@20571.4]
  wire  _T_1516; // @[MemPrimitives.scala 126:35:@20572.4]
  wire  _T_1517; // @[MemPrimitives.scala 126:35:@20573.4]
  wire [10:0] _T_1519; // @[Cat.scala 30:58:@20575.4]
  wire [10:0] _T_1521; // @[Cat.scala 30:58:@20577.4]
  wire [10:0] _T_1523; // @[Cat.scala 30:58:@20579.4]
  wire [10:0] _T_1525; // @[Cat.scala 30:58:@20581.4]
  wire [10:0] _T_1527; // @[Cat.scala 30:58:@20583.4]
  wire [10:0] _T_1529; // @[Cat.scala 30:58:@20585.4]
  wire [10:0] _T_1531; // @[Cat.scala 30:58:@20587.4]
  wire [10:0] _T_1533; // @[Cat.scala 30:58:@20589.4]
  wire [10:0] _T_1535; // @[Cat.scala 30:58:@20591.4]
  wire [10:0] _T_1536; // @[Mux.scala 31:69:@20592.4]
  wire [10:0] _T_1537; // @[Mux.scala 31:69:@20593.4]
  wire [10:0] _T_1538; // @[Mux.scala 31:69:@20594.4]
  wire [10:0] _T_1539; // @[Mux.scala 31:69:@20595.4]
  wire [10:0] _T_1540; // @[Mux.scala 31:69:@20596.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@20597.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@20598.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@20599.4]
  wire  _T_1550; // @[MemPrimitives.scala 110:210:@20607.4]
  wire  _T_1551; // @[MemPrimitives.scala 110:228:@20608.4]
  wire  _T_1556; // @[MemPrimitives.scala 110:210:@20611.4]
  wire  _T_1557; // @[MemPrimitives.scala 110:228:@20612.4]
  wire  _T_1562; // @[MemPrimitives.scala 110:210:@20615.4]
  wire  _T_1563; // @[MemPrimitives.scala 110:228:@20616.4]
  wire  _T_1568; // @[MemPrimitives.scala 110:210:@20619.4]
  wire  _T_1569; // @[MemPrimitives.scala 110:228:@20620.4]
  wire  _T_1574; // @[MemPrimitives.scala 110:210:@20623.4]
  wire  _T_1575; // @[MemPrimitives.scala 110:228:@20624.4]
  wire  _T_1580; // @[MemPrimitives.scala 110:210:@20627.4]
  wire  _T_1581; // @[MemPrimitives.scala 110:228:@20628.4]
  wire  _T_1586; // @[MemPrimitives.scala 110:210:@20631.4]
  wire  _T_1587; // @[MemPrimitives.scala 110:228:@20632.4]
  wire  _T_1592; // @[MemPrimitives.scala 110:210:@20635.4]
  wire  _T_1593; // @[MemPrimitives.scala 110:228:@20636.4]
  wire  _T_1598; // @[MemPrimitives.scala 110:210:@20639.4]
  wire  _T_1599; // @[MemPrimitives.scala 110:228:@20640.4]
  wire  _T_1601; // @[MemPrimitives.scala 126:35:@20654.4]
  wire  _T_1602; // @[MemPrimitives.scala 126:35:@20655.4]
  wire  _T_1603; // @[MemPrimitives.scala 126:35:@20656.4]
  wire  _T_1604; // @[MemPrimitives.scala 126:35:@20657.4]
  wire  _T_1605; // @[MemPrimitives.scala 126:35:@20658.4]
  wire  _T_1606; // @[MemPrimitives.scala 126:35:@20659.4]
  wire  _T_1607; // @[MemPrimitives.scala 126:35:@20660.4]
  wire  _T_1608; // @[MemPrimitives.scala 126:35:@20661.4]
  wire  _T_1609; // @[MemPrimitives.scala 126:35:@20662.4]
  wire [10:0] _T_1611; // @[Cat.scala 30:58:@20664.4]
  wire [10:0] _T_1613; // @[Cat.scala 30:58:@20666.4]
  wire [10:0] _T_1615; // @[Cat.scala 30:58:@20668.4]
  wire [10:0] _T_1617; // @[Cat.scala 30:58:@20670.4]
  wire [10:0] _T_1619; // @[Cat.scala 30:58:@20672.4]
  wire [10:0] _T_1621; // @[Cat.scala 30:58:@20674.4]
  wire [10:0] _T_1623; // @[Cat.scala 30:58:@20676.4]
  wire [10:0] _T_1625; // @[Cat.scala 30:58:@20678.4]
  wire [10:0] _T_1627; // @[Cat.scala 30:58:@20680.4]
  wire [10:0] _T_1628; // @[Mux.scala 31:69:@20681.4]
  wire [10:0] _T_1629; // @[Mux.scala 31:69:@20682.4]
  wire [10:0] _T_1630; // @[Mux.scala 31:69:@20683.4]
  wire [10:0] _T_1631; // @[Mux.scala 31:69:@20684.4]
  wire [10:0] _T_1632; // @[Mux.scala 31:69:@20685.4]
  wire [10:0] _T_1633; // @[Mux.scala 31:69:@20686.4]
  wire [10:0] _T_1634; // @[Mux.scala 31:69:@20687.4]
  wire [10:0] _T_1635; // @[Mux.scala 31:69:@20688.4]
  wire  _T_1642; // @[MemPrimitives.scala 110:210:@20696.4]
  wire  _T_1643; // @[MemPrimitives.scala 110:228:@20697.4]
  wire  _T_1648; // @[MemPrimitives.scala 110:210:@20700.4]
  wire  _T_1649; // @[MemPrimitives.scala 110:228:@20701.4]
  wire  _T_1654; // @[MemPrimitives.scala 110:210:@20704.4]
  wire  _T_1655; // @[MemPrimitives.scala 110:228:@20705.4]
  wire  _T_1660; // @[MemPrimitives.scala 110:210:@20708.4]
  wire  _T_1661; // @[MemPrimitives.scala 110:228:@20709.4]
  wire  _T_1666; // @[MemPrimitives.scala 110:210:@20712.4]
  wire  _T_1667; // @[MemPrimitives.scala 110:228:@20713.4]
  wire  _T_1672; // @[MemPrimitives.scala 110:210:@20716.4]
  wire  _T_1673; // @[MemPrimitives.scala 110:228:@20717.4]
  wire  _T_1678; // @[MemPrimitives.scala 110:210:@20720.4]
  wire  _T_1679; // @[MemPrimitives.scala 110:228:@20721.4]
  wire  _T_1684; // @[MemPrimitives.scala 110:210:@20724.4]
  wire  _T_1685; // @[MemPrimitives.scala 110:228:@20725.4]
  wire  _T_1690; // @[MemPrimitives.scala 110:210:@20728.4]
  wire  _T_1691; // @[MemPrimitives.scala 110:228:@20729.4]
  wire  _T_1693; // @[MemPrimitives.scala 126:35:@20743.4]
  wire  _T_1694; // @[MemPrimitives.scala 126:35:@20744.4]
  wire  _T_1695; // @[MemPrimitives.scala 126:35:@20745.4]
  wire  _T_1696; // @[MemPrimitives.scala 126:35:@20746.4]
  wire  _T_1697; // @[MemPrimitives.scala 126:35:@20747.4]
  wire  _T_1698; // @[MemPrimitives.scala 126:35:@20748.4]
  wire  _T_1699; // @[MemPrimitives.scala 126:35:@20749.4]
  wire  _T_1700; // @[MemPrimitives.scala 126:35:@20750.4]
  wire  _T_1701; // @[MemPrimitives.scala 126:35:@20751.4]
  wire [10:0] _T_1703; // @[Cat.scala 30:58:@20753.4]
  wire [10:0] _T_1705; // @[Cat.scala 30:58:@20755.4]
  wire [10:0] _T_1707; // @[Cat.scala 30:58:@20757.4]
  wire [10:0] _T_1709; // @[Cat.scala 30:58:@20759.4]
  wire [10:0] _T_1711; // @[Cat.scala 30:58:@20761.4]
  wire [10:0] _T_1713; // @[Cat.scala 30:58:@20763.4]
  wire [10:0] _T_1715; // @[Cat.scala 30:58:@20765.4]
  wire [10:0] _T_1717; // @[Cat.scala 30:58:@20767.4]
  wire [10:0] _T_1719; // @[Cat.scala 30:58:@20769.4]
  wire [10:0] _T_1720; // @[Mux.scala 31:69:@20770.4]
  wire [10:0] _T_1721; // @[Mux.scala 31:69:@20771.4]
  wire [10:0] _T_1722; // @[Mux.scala 31:69:@20772.4]
  wire [10:0] _T_1723; // @[Mux.scala 31:69:@20773.4]
  wire [10:0] _T_1724; // @[Mux.scala 31:69:@20774.4]
  wire [10:0] _T_1725; // @[Mux.scala 31:69:@20775.4]
  wire [10:0] _T_1726; // @[Mux.scala 31:69:@20776.4]
  wire [10:0] _T_1727; // @[Mux.scala 31:69:@20777.4]
  wire  _T_1732; // @[MemPrimitives.scala 110:210:@20784.4]
  wire  _T_1735; // @[MemPrimitives.scala 110:228:@20786.4]
  wire  _T_1738; // @[MemPrimitives.scala 110:210:@20788.4]
  wire  _T_1741; // @[MemPrimitives.scala 110:228:@20790.4]
  wire  _T_1744; // @[MemPrimitives.scala 110:210:@20792.4]
  wire  _T_1747; // @[MemPrimitives.scala 110:228:@20794.4]
  wire  _T_1750; // @[MemPrimitives.scala 110:210:@20796.4]
  wire  _T_1753; // @[MemPrimitives.scala 110:228:@20798.4]
  wire  _T_1756; // @[MemPrimitives.scala 110:210:@20800.4]
  wire  _T_1759; // @[MemPrimitives.scala 110:228:@20802.4]
  wire  _T_1762; // @[MemPrimitives.scala 110:210:@20804.4]
  wire  _T_1765; // @[MemPrimitives.scala 110:228:@20806.4]
  wire  _T_1768; // @[MemPrimitives.scala 110:210:@20808.4]
  wire  _T_1771; // @[MemPrimitives.scala 110:228:@20810.4]
  wire  _T_1774; // @[MemPrimitives.scala 110:210:@20812.4]
  wire  _T_1777; // @[MemPrimitives.scala 110:228:@20814.4]
  wire  _T_1780; // @[MemPrimitives.scala 110:210:@20816.4]
  wire  _T_1783; // @[MemPrimitives.scala 110:228:@20818.4]
  wire  _T_1785; // @[MemPrimitives.scala 126:35:@20832.4]
  wire  _T_1786; // @[MemPrimitives.scala 126:35:@20833.4]
  wire  _T_1787; // @[MemPrimitives.scala 126:35:@20834.4]
  wire  _T_1788; // @[MemPrimitives.scala 126:35:@20835.4]
  wire  _T_1789; // @[MemPrimitives.scala 126:35:@20836.4]
  wire  _T_1790; // @[MemPrimitives.scala 126:35:@20837.4]
  wire  _T_1791; // @[MemPrimitives.scala 126:35:@20838.4]
  wire  _T_1792; // @[MemPrimitives.scala 126:35:@20839.4]
  wire  _T_1793; // @[MemPrimitives.scala 126:35:@20840.4]
  wire [10:0] _T_1795; // @[Cat.scala 30:58:@20842.4]
  wire [10:0] _T_1797; // @[Cat.scala 30:58:@20844.4]
  wire [10:0] _T_1799; // @[Cat.scala 30:58:@20846.4]
  wire [10:0] _T_1801; // @[Cat.scala 30:58:@20848.4]
  wire [10:0] _T_1803; // @[Cat.scala 30:58:@20850.4]
  wire [10:0] _T_1805; // @[Cat.scala 30:58:@20852.4]
  wire [10:0] _T_1807; // @[Cat.scala 30:58:@20854.4]
  wire [10:0] _T_1809; // @[Cat.scala 30:58:@20856.4]
  wire [10:0] _T_1811; // @[Cat.scala 30:58:@20858.4]
  wire [10:0] _T_1812; // @[Mux.scala 31:69:@20859.4]
  wire [10:0] _T_1813; // @[Mux.scala 31:69:@20860.4]
  wire [10:0] _T_1814; // @[Mux.scala 31:69:@20861.4]
  wire [10:0] _T_1815; // @[Mux.scala 31:69:@20862.4]
  wire [10:0] _T_1816; // @[Mux.scala 31:69:@20863.4]
  wire [10:0] _T_1817; // @[Mux.scala 31:69:@20864.4]
  wire [10:0] _T_1818; // @[Mux.scala 31:69:@20865.4]
  wire [10:0] _T_1819; // @[Mux.scala 31:69:@20866.4]
  wire  _T_1824; // @[MemPrimitives.scala 110:210:@20873.4]
  wire  _T_1827; // @[MemPrimitives.scala 110:228:@20875.4]
  wire  _T_1830; // @[MemPrimitives.scala 110:210:@20877.4]
  wire  _T_1833; // @[MemPrimitives.scala 110:228:@20879.4]
  wire  _T_1836; // @[MemPrimitives.scala 110:210:@20881.4]
  wire  _T_1839; // @[MemPrimitives.scala 110:228:@20883.4]
  wire  _T_1842; // @[MemPrimitives.scala 110:210:@20885.4]
  wire  _T_1845; // @[MemPrimitives.scala 110:228:@20887.4]
  wire  _T_1848; // @[MemPrimitives.scala 110:210:@20889.4]
  wire  _T_1851; // @[MemPrimitives.scala 110:228:@20891.4]
  wire  _T_1854; // @[MemPrimitives.scala 110:210:@20893.4]
  wire  _T_1857; // @[MemPrimitives.scala 110:228:@20895.4]
  wire  _T_1860; // @[MemPrimitives.scala 110:210:@20897.4]
  wire  _T_1863; // @[MemPrimitives.scala 110:228:@20899.4]
  wire  _T_1866; // @[MemPrimitives.scala 110:210:@20901.4]
  wire  _T_1869; // @[MemPrimitives.scala 110:228:@20903.4]
  wire  _T_1872; // @[MemPrimitives.scala 110:210:@20905.4]
  wire  _T_1875; // @[MemPrimitives.scala 110:228:@20907.4]
  wire  _T_1877; // @[MemPrimitives.scala 126:35:@20921.4]
  wire  _T_1878; // @[MemPrimitives.scala 126:35:@20922.4]
  wire  _T_1879; // @[MemPrimitives.scala 126:35:@20923.4]
  wire  _T_1880; // @[MemPrimitives.scala 126:35:@20924.4]
  wire  _T_1881; // @[MemPrimitives.scala 126:35:@20925.4]
  wire  _T_1882; // @[MemPrimitives.scala 126:35:@20926.4]
  wire  _T_1883; // @[MemPrimitives.scala 126:35:@20927.4]
  wire  _T_1884; // @[MemPrimitives.scala 126:35:@20928.4]
  wire  _T_1885; // @[MemPrimitives.scala 126:35:@20929.4]
  wire [10:0] _T_1887; // @[Cat.scala 30:58:@20931.4]
  wire [10:0] _T_1889; // @[Cat.scala 30:58:@20933.4]
  wire [10:0] _T_1891; // @[Cat.scala 30:58:@20935.4]
  wire [10:0] _T_1893; // @[Cat.scala 30:58:@20937.4]
  wire [10:0] _T_1895; // @[Cat.scala 30:58:@20939.4]
  wire [10:0] _T_1897; // @[Cat.scala 30:58:@20941.4]
  wire [10:0] _T_1899; // @[Cat.scala 30:58:@20943.4]
  wire [10:0] _T_1901; // @[Cat.scala 30:58:@20945.4]
  wire [10:0] _T_1903; // @[Cat.scala 30:58:@20947.4]
  wire [10:0] _T_1904; // @[Mux.scala 31:69:@20948.4]
  wire [10:0] _T_1905; // @[Mux.scala 31:69:@20949.4]
  wire [10:0] _T_1906; // @[Mux.scala 31:69:@20950.4]
  wire [10:0] _T_1907; // @[Mux.scala 31:69:@20951.4]
  wire [10:0] _T_1908; // @[Mux.scala 31:69:@20952.4]
  wire [10:0] _T_1909; // @[Mux.scala 31:69:@20953.4]
  wire [10:0] _T_1910; // @[Mux.scala 31:69:@20954.4]
  wire [10:0] _T_1911; // @[Mux.scala 31:69:@20955.4]
  wire  _T_1919; // @[MemPrimitives.scala 110:228:@20964.4]
  wire  _T_1925; // @[MemPrimitives.scala 110:228:@20968.4]
  wire  _T_1931; // @[MemPrimitives.scala 110:228:@20972.4]
  wire  _T_1937; // @[MemPrimitives.scala 110:228:@20976.4]
  wire  _T_1943; // @[MemPrimitives.scala 110:228:@20980.4]
  wire  _T_1949; // @[MemPrimitives.scala 110:228:@20984.4]
  wire  _T_1955; // @[MemPrimitives.scala 110:228:@20988.4]
  wire  _T_1961; // @[MemPrimitives.scala 110:228:@20992.4]
  wire  _T_1967; // @[MemPrimitives.scala 110:228:@20996.4]
  wire  _T_1969; // @[MemPrimitives.scala 126:35:@21010.4]
  wire  _T_1970; // @[MemPrimitives.scala 126:35:@21011.4]
  wire  _T_1971; // @[MemPrimitives.scala 126:35:@21012.4]
  wire  _T_1972; // @[MemPrimitives.scala 126:35:@21013.4]
  wire  _T_1973; // @[MemPrimitives.scala 126:35:@21014.4]
  wire  _T_1974; // @[MemPrimitives.scala 126:35:@21015.4]
  wire  _T_1975; // @[MemPrimitives.scala 126:35:@21016.4]
  wire  _T_1976; // @[MemPrimitives.scala 126:35:@21017.4]
  wire  _T_1977; // @[MemPrimitives.scala 126:35:@21018.4]
  wire [10:0] _T_1979; // @[Cat.scala 30:58:@21020.4]
  wire [10:0] _T_1981; // @[Cat.scala 30:58:@21022.4]
  wire [10:0] _T_1983; // @[Cat.scala 30:58:@21024.4]
  wire [10:0] _T_1985; // @[Cat.scala 30:58:@21026.4]
  wire [10:0] _T_1987; // @[Cat.scala 30:58:@21028.4]
  wire [10:0] _T_1989; // @[Cat.scala 30:58:@21030.4]
  wire [10:0] _T_1991; // @[Cat.scala 30:58:@21032.4]
  wire [10:0] _T_1993; // @[Cat.scala 30:58:@21034.4]
  wire [10:0] _T_1995; // @[Cat.scala 30:58:@21036.4]
  wire [10:0] _T_1996; // @[Mux.scala 31:69:@21037.4]
  wire [10:0] _T_1997; // @[Mux.scala 31:69:@21038.4]
  wire [10:0] _T_1998; // @[Mux.scala 31:69:@21039.4]
  wire [10:0] _T_1999; // @[Mux.scala 31:69:@21040.4]
  wire [10:0] _T_2000; // @[Mux.scala 31:69:@21041.4]
  wire [10:0] _T_2001; // @[Mux.scala 31:69:@21042.4]
  wire [10:0] _T_2002; // @[Mux.scala 31:69:@21043.4]
  wire [10:0] _T_2003; // @[Mux.scala 31:69:@21044.4]
  wire  _T_2011; // @[MemPrimitives.scala 110:228:@21053.4]
  wire  _T_2017; // @[MemPrimitives.scala 110:228:@21057.4]
  wire  _T_2023; // @[MemPrimitives.scala 110:228:@21061.4]
  wire  _T_2029; // @[MemPrimitives.scala 110:228:@21065.4]
  wire  _T_2035; // @[MemPrimitives.scala 110:228:@21069.4]
  wire  _T_2041; // @[MemPrimitives.scala 110:228:@21073.4]
  wire  _T_2047; // @[MemPrimitives.scala 110:228:@21077.4]
  wire  _T_2053; // @[MemPrimitives.scala 110:228:@21081.4]
  wire  _T_2059; // @[MemPrimitives.scala 110:228:@21085.4]
  wire  _T_2061; // @[MemPrimitives.scala 126:35:@21099.4]
  wire  _T_2062; // @[MemPrimitives.scala 126:35:@21100.4]
  wire  _T_2063; // @[MemPrimitives.scala 126:35:@21101.4]
  wire  _T_2064; // @[MemPrimitives.scala 126:35:@21102.4]
  wire  _T_2065; // @[MemPrimitives.scala 126:35:@21103.4]
  wire  _T_2066; // @[MemPrimitives.scala 126:35:@21104.4]
  wire  _T_2067; // @[MemPrimitives.scala 126:35:@21105.4]
  wire  _T_2068; // @[MemPrimitives.scala 126:35:@21106.4]
  wire  _T_2069; // @[MemPrimitives.scala 126:35:@21107.4]
  wire [10:0] _T_2071; // @[Cat.scala 30:58:@21109.4]
  wire [10:0] _T_2073; // @[Cat.scala 30:58:@21111.4]
  wire [10:0] _T_2075; // @[Cat.scala 30:58:@21113.4]
  wire [10:0] _T_2077; // @[Cat.scala 30:58:@21115.4]
  wire [10:0] _T_2079; // @[Cat.scala 30:58:@21117.4]
  wire [10:0] _T_2081; // @[Cat.scala 30:58:@21119.4]
  wire [10:0] _T_2083; // @[Cat.scala 30:58:@21121.4]
  wire [10:0] _T_2085; // @[Cat.scala 30:58:@21123.4]
  wire [10:0] _T_2087; // @[Cat.scala 30:58:@21125.4]
  wire [10:0] _T_2088; // @[Mux.scala 31:69:@21126.4]
  wire [10:0] _T_2089; // @[Mux.scala 31:69:@21127.4]
  wire [10:0] _T_2090; // @[Mux.scala 31:69:@21128.4]
  wire [10:0] _T_2091; // @[Mux.scala 31:69:@21129.4]
  wire [10:0] _T_2092; // @[Mux.scala 31:69:@21130.4]
  wire [10:0] _T_2093; // @[Mux.scala 31:69:@21131.4]
  wire [10:0] _T_2094; // @[Mux.scala 31:69:@21132.4]
  wire [10:0] _T_2095; // @[Mux.scala 31:69:@21133.4]
  wire  _T_2103; // @[MemPrimitives.scala 110:228:@21142.4]
  wire  _T_2109; // @[MemPrimitives.scala 110:228:@21146.4]
  wire  _T_2115; // @[MemPrimitives.scala 110:228:@21150.4]
  wire  _T_2121; // @[MemPrimitives.scala 110:228:@21154.4]
  wire  _T_2127; // @[MemPrimitives.scala 110:228:@21158.4]
  wire  _T_2133; // @[MemPrimitives.scala 110:228:@21162.4]
  wire  _T_2139; // @[MemPrimitives.scala 110:228:@21166.4]
  wire  _T_2145; // @[MemPrimitives.scala 110:228:@21170.4]
  wire  _T_2151; // @[MemPrimitives.scala 110:228:@21174.4]
  wire  _T_2153; // @[MemPrimitives.scala 126:35:@21188.4]
  wire  _T_2154; // @[MemPrimitives.scala 126:35:@21189.4]
  wire  _T_2155; // @[MemPrimitives.scala 126:35:@21190.4]
  wire  _T_2156; // @[MemPrimitives.scala 126:35:@21191.4]
  wire  _T_2157; // @[MemPrimitives.scala 126:35:@21192.4]
  wire  _T_2158; // @[MemPrimitives.scala 126:35:@21193.4]
  wire  _T_2159; // @[MemPrimitives.scala 126:35:@21194.4]
  wire  _T_2160; // @[MemPrimitives.scala 126:35:@21195.4]
  wire  _T_2161; // @[MemPrimitives.scala 126:35:@21196.4]
  wire [10:0] _T_2163; // @[Cat.scala 30:58:@21198.4]
  wire [10:0] _T_2165; // @[Cat.scala 30:58:@21200.4]
  wire [10:0] _T_2167; // @[Cat.scala 30:58:@21202.4]
  wire [10:0] _T_2169; // @[Cat.scala 30:58:@21204.4]
  wire [10:0] _T_2171; // @[Cat.scala 30:58:@21206.4]
  wire [10:0] _T_2173; // @[Cat.scala 30:58:@21208.4]
  wire [10:0] _T_2175; // @[Cat.scala 30:58:@21210.4]
  wire [10:0] _T_2177; // @[Cat.scala 30:58:@21212.4]
  wire [10:0] _T_2179; // @[Cat.scala 30:58:@21214.4]
  wire [10:0] _T_2180; // @[Mux.scala 31:69:@21215.4]
  wire [10:0] _T_2181; // @[Mux.scala 31:69:@21216.4]
  wire [10:0] _T_2182; // @[Mux.scala 31:69:@21217.4]
  wire [10:0] _T_2183; // @[Mux.scala 31:69:@21218.4]
  wire [10:0] _T_2184; // @[Mux.scala 31:69:@21219.4]
  wire [10:0] _T_2185; // @[Mux.scala 31:69:@21220.4]
  wire [10:0] _T_2186; // @[Mux.scala 31:69:@21221.4]
  wire [10:0] _T_2187; // @[Mux.scala 31:69:@21222.4]
  wire  _T_2195; // @[MemPrimitives.scala 110:228:@21231.4]
  wire  _T_2201; // @[MemPrimitives.scala 110:228:@21235.4]
  wire  _T_2207; // @[MemPrimitives.scala 110:228:@21239.4]
  wire  _T_2213; // @[MemPrimitives.scala 110:228:@21243.4]
  wire  _T_2219; // @[MemPrimitives.scala 110:228:@21247.4]
  wire  _T_2225; // @[MemPrimitives.scala 110:228:@21251.4]
  wire  _T_2231; // @[MemPrimitives.scala 110:228:@21255.4]
  wire  _T_2237; // @[MemPrimitives.scala 110:228:@21259.4]
  wire  _T_2243; // @[MemPrimitives.scala 110:228:@21263.4]
  wire  _T_2245; // @[MemPrimitives.scala 126:35:@21277.4]
  wire  _T_2246; // @[MemPrimitives.scala 126:35:@21278.4]
  wire  _T_2247; // @[MemPrimitives.scala 126:35:@21279.4]
  wire  _T_2248; // @[MemPrimitives.scala 126:35:@21280.4]
  wire  _T_2249; // @[MemPrimitives.scala 126:35:@21281.4]
  wire  _T_2250; // @[MemPrimitives.scala 126:35:@21282.4]
  wire  _T_2251; // @[MemPrimitives.scala 126:35:@21283.4]
  wire  _T_2252; // @[MemPrimitives.scala 126:35:@21284.4]
  wire  _T_2253; // @[MemPrimitives.scala 126:35:@21285.4]
  wire [10:0] _T_2255; // @[Cat.scala 30:58:@21287.4]
  wire [10:0] _T_2257; // @[Cat.scala 30:58:@21289.4]
  wire [10:0] _T_2259; // @[Cat.scala 30:58:@21291.4]
  wire [10:0] _T_2261; // @[Cat.scala 30:58:@21293.4]
  wire [10:0] _T_2263; // @[Cat.scala 30:58:@21295.4]
  wire [10:0] _T_2265; // @[Cat.scala 30:58:@21297.4]
  wire [10:0] _T_2267; // @[Cat.scala 30:58:@21299.4]
  wire [10:0] _T_2269; // @[Cat.scala 30:58:@21301.4]
  wire [10:0] _T_2271; // @[Cat.scala 30:58:@21303.4]
  wire [10:0] _T_2272; // @[Mux.scala 31:69:@21304.4]
  wire [10:0] _T_2273; // @[Mux.scala 31:69:@21305.4]
  wire [10:0] _T_2274; // @[Mux.scala 31:69:@21306.4]
  wire [10:0] _T_2275; // @[Mux.scala 31:69:@21307.4]
  wire [10:0] _T_2276; // @[Mux.scala 31:69:@21308.4]
  wire [10:0] _T_2277; // @[Mux.scala 31:69:@21309.4]
  wire [10:0] _T_2278; // @[Mux.scala 31:69:@21310.4]
  wire [10:0] _T_2279; // @[Mux.scala 31:69:@21311.4]
  wire  _T_2284; // @[MemPrimitives.scala 110:210:@21318.4]
  wire  _T_2287; // @[MemPrimitives.scala 110:228:@21320.4]
  wire  _T_2290; // @[MemPrimitives.scala 110:210:@21322.4]
  wire  _T_2293; // @[MemPrimitives.scala 110:228:@21324.4]
  wire  _T_2296; // @[MemPrimitives.scala 110:210:@21326.4]
  wire  _T_2299; // @[MemPrimitives.scala 110:228:@21328.4]
  wire  _T_2302; // @[MemPrimitives.scala 110:210:@21330.4]
  wire  _T_2305; // @[MemPrimitives.scala 110:228:@21332.4]
  wire  _T_2308; // @[MemPrimitives.scala 110:210:@21334.4]
  wire  _T_2311; // @[MemPrimitives.scala 110:228:@21336.4]
  wire  _T_2314; // @[MemPrimitives.scala 110:210:@21338.4]
  wire  _T_2317; // @[MemPrimitives.scala 110:228:@21340.4]
  wire  _T_2320; // @[MemPrimitives.scala 110:210:@21342.4]
  wire  _T_2323; // @[MemPrimitives.scala 110:228:@21344.4]
  wire  _T_2326; // @[MemPrimitives.scala 110:210:@21346.4]
  wire  _T_2329; // @[MemPrimitives.scala 110:228:@21348.4]
  wire  _T_2332; // @[MemPrimitives.scala 110:210:@21350.4]
  wire  _T_2335; // @[MemPrimitives.scala 110:228:@21352.4]
  wire  _T_2337; // @[MemPrimitives.scala 126:35:@21366.4]
  wire  _T_2338; // @[MemPrimitives.scala 126:35:@21367.4]
  wire  _T_2339; // @[MemPrimitives.scala 126:35:@21368.4]
  wire  _T_2340; // @[MemPrimitives.scala 126:35:@21369.4]
  wire  _T_2341; // @[MemPrimitives.scala 126:35:@21370.4]
  wire  _T_2342; // @[MemPrimitives.scala 126:35:@21371.4]
  wire  _T_2343; // @[MemPrimitives.scala 126:35:@21372.4]
  wire  _T_2344; // @[MemPrimitives.scala 126:35:@21373.4]
  wire  _T_2345; // @[MemPrimitives.scala 126:35:@21374.4]
  wire [10:0] _T_2347; // @[Cat.scala 30:58:@21376.4]
  wire [10:0] _T_2349; // @[Cat.scala 30:58:@21378.4]
  wire [10:0] _T_2351; // @[Cat.scala 30:58:@21380.4]
  wire [10:0] _T_2353; // @[Cat.scala 30:58:@21382.4]
  wire [10:0] _T_2355; // @[Cat.scala 30:58:@21384.4]
  wire [10:0] _T_2357; // @[Cat.scala 30:58:@21386.4]
  wire [10:0] _T_2359; // @[Cat.scala 30:58:@21388.4]
  wire [10:0] _T_2361; // @[Cat.scala 30:58:@21390.4]
  wire [10:0] _T_2363; // @[Cat.scala 30:58:@21392.4]
  wire [10:0] _T_2364; // @[Mux.scala 31:69:@21393.4]
  wire [10:0] _T_2365; // @[Mux.scala 31:69:@21394.4]
  wire [10:0] _T_2366; // @[Mux.scala 31:69:@21395.4]
  wire [10:0] _T_2367; // @[Mux.scala 31:69:@21396.4]
  wire [10:0] _T_2368; // @[Mux.scala 31:69:@21397.4]
  wire [10:0] _T_2369; // @[Mux.scala 31:69:@21398.4]
  wire [10:0] _T_2370; // @[Mux.scala 31:69:@21399.4]
  wire [10:0] _T_2371; // @[Mux.scala 31:69:@21400.4]
  wire  _T_2376; // @[MemPrimitives.scala 110:210:@21407.4]
  wire  _T_2379; // @[MemPrimitives.scala 110:228:@21409.4]
  wire  _T_2382; // @[MemPrimitives.scala 110:210:@21411.4]
  wire  _T_2385; // @[MemPrimitives.scala 110:228:@21413.4]
  wire  _T_2388; // @[MemPrimitives.scala 110:210:@21415.4]
  wire  _T_2391; // @[MemPrimitives.scala 110:228:@21417.4]
  wire  _T_2394; // @[MemPrimitives.scala 110:210:@21419.4]
  wire  _T_2397; // @[MemPrimitives.scala 110:228:@21421.4]
  wire  _T_2400; // @[MemPrimitives.scala 110:210:@21423.4]
  wire  _T_2403; // @[MemPrimitives.scala 110:228:@21425.4]
  wire  _T_2406; // @[MemPrimitives.scala 110:210:@21427.4]
  wire  _T_2409; // @[MemPrimitives.scala 110:228:@21429.4]
  wire  _T_2412; // @[MemPrimitives.scala 110:210:@21431.4]
  wire  _T_2415; // @[MemPrimitives.scala 110:228:@21433.4]
  wire  _T_2418; // @[MemPrimitives.scala 110:210:@21435.4]
  wire  _T_2421; // @[MemPrimitives.scala 110:228:@21437.4]
  wire  _T_2424; // @[MemPrimitives.scala 110:210:@21439.4]
  wire  _T_2427; // @[MemPrimitives.scala 110:228:@21441.4]
  wire  _T_2429; // @[MemPrimitives.scala 126:35:@21455.4]
  wire  _T_2430; // @[MemPrimitives.scala 126:35:@21456.4]
  wire  _T_2431; // @[MemPrimitives.scala 126:35:@21457.4]
  wire  _T_2432; // @[MemPrimitives.scala 126:35:@21458.4]
  wire  _T_2433; // @[MemPrimitives.scala 126:35:@21459.4]
  wire  _T_2434; // @[MemPrimitives.scala 126:35:@21460.4]
  wire  _T_2435; // @[MemPrimitives.scala 126:35:@21461.4]
  wire  _T_2436; // @[MemPrimitives.scala 126:35:@21462.4]
  wire  _T_2437; // @[MemPrimitives.scala 126:35:@21463.4]
  wire [10:0] _T_2439; // @[Cat.scala 30:58:@21465.4]
  wire [10:0] _T_2441; // @[Cat.scala 30:58:@21467.4]
  wire [10:0] _T_2443; // @[Cat.scala 30:58:@21469.4]
  wire [10:0] _T_2445; // @[Cat.scala 30:58:@21471.4]
  wire [10:0] _T_2447; // @[Cat.scala 30:58:@21473.4]
  wire [10:0] _T_2449; // @[Cat.scala 30:58:@21475.4]
  wire [10:0] _T_2451; // @[Cat.scala 30:58:@21477.4]
  wire [10:0] _T_2453; // @[Cat.scala 30:58:@21479.4]
  wire [10:0] _T_2455; // @[Cat.scala 30:58:@21481.4]
  wire [10:0] _T_2456; // @[Mux.scala 31:69:@21482.4]
  wire [10:0] _T_2457; // @[Mux.scala 31:69:@21483.4]
  wire [10:0] _T_2458; // @[Mux.scala 31:69:@21484.4]
  wire [10:0] _T_2459; // @[Mux.scala 31:69:@21485.4]
  wire [10:0] _T_2460; // @[Mux.scala 31:69:@21486.4]
  wire [10:0] _T_2461; // @[Mux.scala 31:69:@21487.4]
  wire [10:0] _T_2462; // @[Mux.scala 31:69:@21488.4]
  wire [10:0] _T_2463; // @[Mux.scala 31:69:@21489.4]
  wire  _T_2471; // @[MemPrimitives.scala 110:228:@21498.4]
  wire  _T_2477; // @[MemPrimitives.scala 110:228:@21502.4]
  wire  _T_2483; // @[MemPrimitives.scala 110:228:@21506.4]
  wire  _T_2489; // @[MemPrimitives.scala 110:228:@21510.4]
  wire  _T_2495; // @[MemPrimitives.scala 110:228:@21514.4]
  wire  _T_2501; // @[MemPrimitives.scala 110:228:@21518.4]
  wire  _T_2507; // @[MemPrimitives.scala 110:228:@21522.4]
  wire  _T_2513; // @[MemPrimitives.scala 110:228:@21526.4]
  wire  _T_2519; // @[MemPrimitives.scala 110:228:@21530.4]
  wire  _T_2521; // @[MemPrimitives.scala 126:35:@21544.4]
  wire  _T_2522; // @[MemPrimitives.scala 126:35:@21545.4]
  wire  _T_2523; // @[MemPrimitives.scala 126:35:@21546.4]
  wire  _T_2524; // @[MemPrimitives.scala 126:35:@21547.4]
  wire  _T_2525; // @[MemPrimitives.scala 126:35:@21548.4]
  wire  _T_2526; // @[MemPrimitives.scala 126:35:@21549.4]
  wire  _T_2527; // @[MemPrimitives.scala 126:35:@21550.4]
  wire  _T_2528; // @[MemPrimitives.scala 126:35:@21551.4]
  wire  _T_2529; // @[MemPrimitives.scala 126:35:@21552.4]
  wire [10:0] _T_2531; // @[Cat.scala 30:58:@21554.4]
  wire [10:0] _T_2533; // @[Cat.scala 30:58:@21556.4]
  wire [10:0] _T_2535; // @[Cat.scala 30:58:@21558.4]
  wire [10:0] _T_2537; // @[Cat.scala 30:58:@21560.4]
  wire [10:0] _T_2539; // @[Cat.scala 30:58:@21562.4]
  wire [10:0] _T_2541; // @[Cat.scala 30:58:@21564.4]
  wire [10:0] _T_2543; // @[Cat.scala 30:58:@21566.4]
  wire [10:0] _T_2545; // @[Cat.scala 30:58:@21568.4]
  wire [10:0] _T_2547; // @[Cat.scala 30:58:@21570.4]
  wire [10:0] _T_2548; // @[Mux.scala 31:69:@21571.4]
  wire [10:0] _T_2549; // @[Mux.scala 31:69:@21572.4]
  wire [10:0] _T_2550; // @[Mux.scala 31:69:@21573.4]
  wire [10:0] _T_2551; // @[Mux.scala 31:69:@21574.4]
  wire [10:0] _T_2552; // @[Mux.scala 31:69:@21575.4]
  wire [10:0] _T_2553; // @[Mux.scala 31:69:@21576.4]
  wire [10:0] _T_2554; // @[Mux.scala 31:69:@21577.4]
  wire [10:0] _T_2555; // @[Mux.scala 31:69:@21578.4]
  wire  _T_2563; // @[MemPrimitives.scala 110:228:@21587.4]
  wire  _T_2569; // @[MemPrimitives.scala 110:228:@21591.4]
  wire  _T_2575; // @[MemPrimitives.scala 110:228:@21595.4]
  wire  _T_2581; // @[MemPrimitives.scala 110:228:@21599.4]
  wire  _T_2587; // @[MemPrimitives.scala 110:228:@21603.4]
  wire  _T_2593; // @[MemPrimitives.scala 110:228:@21607.4]
  wire  _T_2599; // @[MemPrimitives.scala 110:228:@21611.4]
  wire  _T_2605; // @[MemPrimitives.scala 110:228:@21615.4]
  wire  _T_2611; // @[MemPrimitives.scala 110:228:@21619.4]
  wire  _T_2613; // @[MemPrimitives.scala 126:35:@21633.4]
  wire  _T_2614; // @[MemPrimitives.scala 126:35:@21634.4]
  wire  _T_2615; // @[MemPrimitives.scala 126:35:@21635.4]
  wire  _T_2616; // @[MemPrimitives.scala 126:35:@21636.4]
  wire  _T_2617; // @[MemPrimitives.scala 126:35:@21637.4]
  wire  _T_2618; // @[MemPrimitives.scala 126:35:@21638.4]
  wire  _T_2619; // @[MemPrimitives.scala 126:35:@21639.4]
  wire  _T_2620; // @[MemPrimitives.scala 126:35:@21640.4]
  wire  _T_2621; // @[MemPrimitives.scala 126:35:@21641.4]
  wire [10:0] _T_2623; // @[Cat.scala 30:58:@21643.4]
  wire [10:0] _T_2625; // @[Cat.scala 30:58:@21645.4]
  wire [10:0] _T_2627; // @[Cat.scala 30:58:@21647.4]
  wire [10:0] _T_2629; // @[Cat.scala 30:58:@21649.4]
  wire [10:0] _T_2631; // @[Cat.scala 30:58:@21651.4]
  wire [10:0] _T_2633; // @[Cat.scala 30:58:@21653.4]
  wire [10:0] _T_2635; // @[Cat.scala 30:58:@21655.4]
  wire [10:0] _T_2637; // @[Cat.scala 30:58:@21657.4]
  wire [10:0] _T_2639; // @[Cat.scala 30:58:@21659.4]
  wire [10:0] _T_2640; // @[Mux.scala 31:69:@21660.4]
  wire [10:0] _T_2641; // @[Mux.scala 31:69:@21661.4]
  wire [10:0] _T_2642; // @[Mux.scala 31:69:@21662.4]
  wire [10:0] _T_2643; // @[Mux.scala 31:69:@21663.4]
  wire [10:0] _T_2644; // @[Mux.scala 31:69:@21664.4]
  wire [10:0] _T_2645; // @[Mux.scala 31:69:@21665.4]
  wire [10:0] _T_2646; // @[Mux.scala 31:69:@21666.4]
  wire [10:0] _T_2647; // @[Mux.scala 31:69:@21667.4]
  wire  _T_2655; // @[MemPrimitives.scala 110:228:@21676.4]
  wire  _T_2661; // @[MemPrimitives.scala 110:228:@21680.4]
  wire  _T_2667; // @[MemPrimitives.scala 110:228:@21684.4]
  wire  _T_2673; // @[MemPrimitives.scala 110:228:@21688.4]
  wire  _T_2679; // @[MemPrimitives.scala 110:228:@21692.4]
  wire  _T_2685; // @[MemPrimitives.scala 110:228:@21696.4]
  wire  _T_2691; // @[MemPrimitives.scala 110:228:@21700.4]
  wire  _T_2697; // @[MemPrimitives.scala 110:228:@21704.4]
  wire  _T_2703; // @[MemPrimitives.scala 110:228:@21708.4]
  wire  _T_2705; // @[MemPrimitives.scala 126:35:@21722.4]
  wire  _T_2706; // @[MemPrimitives.scala 126:35:@21723.4]
  wire  _T_2707; // @[MemPrimitives.scala 126:35:@21724.4]
  wire  _T_2708; // @[MemPrimitives.scala 126:35:@21725.4]
  wire  _T_2709; // @[MemPrimitives.scala 126:35:@21726.4]
  wire  _T_2710; // @[MemPrimitives.scala 126:35:@21727.4]
  wire  _T_2711; // @[MemPrimitives.scala 126:35:@21728.4]
  wire  _T_2712; // @[MemPrimitives.scala 126:35:@21729.4]
  wire  _T_2713; // @[MemPrimitives.scala 126:35:@21730.4]
  wire [10:0] _T_2715; // @[Cat.scala 30:58:@21732.4]
  wire [10:0] _T_2717; // @[Cat.scala 30:58:@21734.4]
  wire [10:0] _T_2719; // @[Cat.scala 30:58:@21736.4]
  wire [10:0] _T_2721; // @[Cat.scala 30:58:@21738.4]
  wire [10:0] _T_2723; // @[Cat.scala 30:58:@21740.4]
  wire [10:0] _T_2725; // @[Cat.scala 30:58:@21742.4]
  wire [10:0] _T_2727; // @[Cat.scala 30:58:@21744.4]
  wire [10:0] _T_2729; // @[Cat.scala 30:58:@21746.4]
  wire [10:0] _T_2731; // @[Cat.scala 30:58:@21748.4]
  wire [10:0] _T_2732; // @[Mux.scala 31:69:@21749.4]
  wire [10:0] _T_2733; // @[Mux.scala 31:69:@21750.4]
  wire [10:0] _T_2734; // @[Mux.scala 31:69:@21751.4]
  wire [10:0] _T_2735; // @[Mux.scala 31:69:@21752.4]
  wire [10:0] _T_2736; // @[Mux.scala 31:69:@21753.4]
  wire [10:0] _T_2737; // @[Mux.scala 31:69:@21754.4]
  wire [10:0] _T_2738; // @[Mux.scala 31:69:@21755.4]
  wire [10:0] _T_2739; // @[Mux.scala 31:69:@21756.4]
  wire  _T_2747; // @[MemPrimitives.scala 110:228:@21765.4]
  wire  _T_2753; // @[MemPrimitives.scala 110:228:@21769.4]
  wire  _T_2759; // @[MemPrimitives.scala 110:228:@21773.4]
  wire  _T_2765; // @[MemPrimitives.scala 110:228:@21777.4]
  wire  _T_2771; // @[MemPrimitives.scala 110:228:@21781.4]
  wire  _T_2777; // @[MemPrimitives.scala 110:228:@21785.4]
  wire  _T_2783; // @[MemPrimitives.scala 110:228:@21789.4]
  wire  _T_2789; // @[MemPrimitives.scala 110:228:@21793.4]
  wire  _T_2795; // @[MemPrimitives.scala 110:228:@21797.4]
  wire  _T_2797; // @[MemPrimitives.scala 126:35:@21811.4]
  wire  _T_2798; // @[MemPrimitives.scala 126:35:@21812.4]
  wire  _T_2799; // @[MemPrimitives.scala 126:35:@21813.4]
  wire  _T_2800; // @[MemPrimitives.scala 126:35:@21814.4]
  wire  _T_2801; // @[MemPrimitives.scala 126:35:@21815.4]
  wire  _T_2802; // @[MemPrimitives.scala 126:35:@21816.4]
  wire  _T_2803; // @[MemPrimitives.scala 126:35:@21817.4]
  wire  _T_2804; // @[MemPrimitives.scala 126:35:@21818.4]
  wire  _T_2805; // @[MemPrimitives.scala 126:35:@21819.4]
  wire [10:0] _T_2807; // @[Cat.scala 30:58:@21821.4]
  wire [10:0] _T_2809; // @[Cat.scala 30:58:@21823.4]
  wire [10:0] _T_2811; // @[Cat.scala 30:58:@21825.4]
  wire [10:0] _T_2813; // @[Cat.scala 30:58:@21827.4]
  wire [10:0] _T_2815; // @[Cat.scala 30:58:@21829.4]
  wire [10:0] _T_2817; // @[Cat.scala 30:58:@21831.4]
  wire [10:0] _T_2819; // @[Cat.scala 30:58:@21833.4]
  wire [10:0] _T_2821; // @[Cat.scala 30:58:@21835.4]
  wire [10:0] _T_2823; // @[Cat.scala 30:58:@21837.4]
  wire [10:0] _T_2824; // @[Mux.scala 31:69:@21838.4]
  wire [10:0] _T_2825; // @[Mux.scala 31:69:@21839.4]
  wire [10:0] _T_2826; // @[Mux.scala 31:69:@21840.4]
  wire [10:0] _T_2827; // @[Mux.scala 31:69:@21841.4]
  wire [10:0] _T_2828; // @[Mux.scala 31:69:@21842.4]
  wire [10:0] _T_2829; // @[Mux.scala 31:69:@21843.4]
  wire [10:0] _T_2830; // @[Mux.scala 31:69:@21844.4]
  wire [10:0] _T_2831; // @[Mux.scala 31:69:@21845.4]
  wire  _T_2836; // @[MemPrimitives.scala 110:210:@21852.4]
  wire  _T_2839; // @[MemPrimitives.scala 110:228:@21854.4]
  wire  _T_2842; // @[MemPrimitives.scala 110:210:@21856.4]
  wire  _T_2845; // @[MemPrimitives.scala 110:228:@21858.4]
  wire  _T_2848; // @[MemPrimitives.scala 110:210:@21860.4]
  wire  _T_2851; // @[MemPrimitives.scala 110:228:@21862.4]
  wire  _T_2854; // @[MemPrimitives.scala 110:210:@21864.4]
  wire  _T_2857; // @[MemPrimitives.scala 110:228:@21866.4]
  wire  _T_2860; // @[MemPrimitives.scala 110:210:@21868.4]
  wire  _T_2863; // @[MemPrimitives.scala 110:228:@21870.4]
  wire  _T_2866; // @[MemPrimitives.scala 110:210:@21872.4]
  wire  _T_2869; // @[MemPrimitives.scala 110:228:@21874.4]
  wire  _T_2872; // @[MemPrimitives.scala 110:210:@21876.4]
  wire  _T_2875; // @[MemPrimitives.scala 110:228:@21878.4]
  wire  _T_2878; // @[MemPrimitives.scala 110:210:@21880.4]
  wire  _T_2881; // @[MemPrimitives.scala 110:228:@21882.4]
  wire  _T_2884; // @[MemPrimitives.scala 110:210:@21884.4]
  wire  _T_2887; // @[MemPrimitives.scala 110:228:@21886.4]
  wire  _T_2889; // @[MemPrimitives.scala 126:35:@21900.4]
  wire  _T_2890; // @[MemPrimitives.scala 126:35:@21901.4]
  wire  _T_2891; // @[MemPrimitives.scala 126:35:@21902.4]
  wire  _T_2892; // @[MemPrimitives.scala 126:35:@21903.4]
  wire  _T_2893; // @[MemPrimitives.scala 126:35:@21904.4]
  wire  _T_2894; // @[MemPrimitives.scala 126:35:@21905.4]
  wire  _T_2895; // @[MemPrimitives.scala 126:35:@21906.4]
  wire  _T_2896; // @[MemPrimitives.scala 126:35:@21907.4]
  wire  _T_2897; // @[MemPrimitives.scala 126:35:@21908.4]
  wire [10:0] _T_2899; // @[Cat.scala 30:58:@21910.4]
  wire [10:0] _T_2901; // @[Cat.scala 30:58:@21912.4]
  wire [10:0] _T_2903; // @[Cat.scala 30:58:@21914.4]
  wire [10:0] _T_2905; // @[Cat.scala 30:58:@21916.4]
  wire [10:0] _T_2907; // @[Cat.scala 30:58:@21918.4]
  wire [10:0] _T_2909; // @[Cat.scala 30:58:@21920.4]
  wire [10:0] _T_2911; // @[Cat.scala 30:58:@21922.4]
  wire [10:0] _T_2913; // @[Cat.scala 30:58:@21924.4]
  wire [10:0] _T_2915; // @[Cat.scala 30:58:@21926.4]
  wire [10:0] _T_2916; // @[Mux.scala 31:69:@21927.4]
  wire [10:0] _T_2917; // @[Mux.scala 31:69:@21928.4]
  wire [10:0] _T_2918; // @[Mux.scala 31:69:@21929.4]
  wire [10:0] _T_2919; // @[Mux.scala 31:69:@21930.4]
  wire [10:0] _T_2920; // @[Mux.scala 31:69:@21931.4]
  wire [10:0] _T_2921; // @[Mux.scala 31:69:@21932.4]
  wire [10:0] _T_2922; // @[Mux.scala 31:69:@21933.4]
  wire [10:0] _T_2923; // @[Mux.scala 31:69:@21934.4]
  wire  _T_2928; // @[MemPrimitives.scala 110:210:@21941.4]
  wire  _T_2931; // @[MemPrimitives.scala 110:228:@21943.4]
  wire  _T_2934; // @[MemPrimitives.scala 110:210:@21945.4]
  wire  _T_2937; // @[MemPrimitives.scala 110:228:@21947.4]
  wire  _T_2940; // @[MemPrimitives.scala 110:210:@21949.4]
  wire  _T_2943; // @[MemPrimitives.scala 110:228:@21951.4]
  wire  _T_2946; // @[MemPrimitives.scala 110:210:@21953.4]
  wire  _T_2949; // @[MemPrimitives.scala 110:228:@21955.4]
  wire  _T_2952; // @[MemPrimitives.scala 110:210:@21957.4]
  wire  _T_2955; // @[MemPrimitives.scala 110:228:@21959.4]
  wire  _T_2958; // @[MemPrimitives.scala 110:210:@21961.4]
  wire  _T_2961; // @[MemPrimitives.scala 110:228:@21963.4]
  wire  _T_2964; // @[MemPrimitives.scala 110:210:@21965.4]
  wire  _T_2967; // @[MemPrimitives.scala 110:228:@21967.4]
  wire  _T_2970; // @[MemPrimitives.scala 110:210:@21969.4]
  wire  _T_2973; // @[MemPrimitives.scala 110:228:@21971.4]
  wire  _T_2976; // @[MemPrimitives.scala 110:210:@21973.4]
  wire  _T_2979; // @[MemPrimitives.scala 110:228:@21975.4]
  wire  _T_2981; // @[MemPrimitives.scala 126:35:@21989.4]
  wire  _T_2982; // @[MemPrimitives.scala 126:35:@21990.4]
  wire  _T_2983; // @[MemPrimitives.scala 126:35:@21991.4]
  wire  _T_2984; // @[MemPrimitives.scala 126:35:@21992.4]
  wire  _T_2985; // @[MemPrimitives.scala 126:35:@21993.4]
  wire  _T_2986; // @[MemPrimitives.scala 126:35:@21994.4]
  wire  _T_2987; // @[MemPrimitives.scala 126:35:@21995.4]
  wire  _T_2988; // @[MemPrimitives.scala 126:35:@21996.4]
  wire  _T_2989; // @[MemPrimitives.scala 126:35:@21997.4]
  wire [10:0] _T_2991; // @[Cat.scala 30:58:@21999.4]
  wire [10:0] _T_2993; // @[Cat.scala 30:58:@22001.4]
  wire [10:0] _T_2995; // @[Cat.scala 30:58:@22003.4]
  wire [10:0] _T_2997; // @[Cat.scala 30:58:@22005.4]
  wire [10:0] _T_2999; // @[Cat.scala 30:58:@22007.4]
  wire [10:0] _T_3001; // @[Cat.scala 30:58:@22009.4]
  wire [10:0] _T_3003; // @[Cat.scala 30:58:@22011.4]
  wire [10:0] _T_3005; // @[Cat.scala 30:58:@22013.4]
  wire [10:0] _T_3007; // @[Cat.scala 30:58:@22015.4]
  wire [10:0] _T_3008; // @[Mux.scala 31:69:@22016.4]
  wire [10:0] _T_3009; // @[Mux.scala 31:69:@22017.4]
  wire [10:0] _T_3010; // @[Mux.scala 31:69:@22018.4]
  wire [10:0] _T_3011; // @[Mux.scala 31:69:@22019.4]
  wire [10:0] _T_3012; // @[Mux.scala 31:69:@22020.4]
  wire [10:0] _T_3013; // @[Mux.scala 31:69:@22021.4]
  wire [10:0] _T_3014; // @[Mux.scala 31:69:@22022.4]
  wire [10:0] _T_3015; // @[Mux.scala 31:69:@22023.4]
  wire  _T_3023; // @[MemPrimitives.scala 110:228:@22032.4]
  wire  _T_3029; // @[MemPrimitives.scala 110:228:@22036.4]
  wire  _T_3035; // @[MemPrimitives.scala 110:228:@22040.4]
  wire  _T_3041; // @[MemPrimitives.scala 110:228:@22044.4]
  wire  _T_3047; // @[MemPrimitives.scala 110:228:@22048.4]
  wire  _T_3053; // @[MemPrimitives.scala 110:228:@22052.4]
  wire  _T_3059; // @[MemPrimitives.scala 110:228:@22056.4]
  wire  _T_3065; // @[MemPrimitives.scala 110:228:@22060.4]
  wire  _T_3071; // @[MemPrimitives.scala 110:228:@22064.4]
  wire  _T_3073; // @[MemPrimitives.scala 126:35:@22078.4]
  wire  _T_3074; // @[MemPrimitives.scala 126:35:@22079.4]
  wire  _T_3075; // @[MemPrimitives.scala 126:35:@22080.4]
  wire  _T_3076; // @[MemPrimitives.scala 126:35:@22081.4]
  wire  _T_3077; // @[MemPrimitives.scala 126:35:@22082.4]
  wire  _T_3078; // @[MemPrimitives.scala 126:35:@22083.4]
  wire  _T_3079; // @[MemPrimitives.scala 126:35:@22084.4]
  wire  _T_3080; // @[MemPrimitives.scala 126:35:@22085.4]
  wire  _T_3081; // @[MemPrimitives.scala 126:35:@22086.4]
  wire [10:0] _T_3083; // @[Cat.scala 30:58:@22088.4]
  wire [10:0] _T_3085; // @[Cat.scala 30:58:@22090.4]
  wire [10:0] _T_3087; // @[Cat.scala 30:58:@22092.4]
  wire [10:0] _T_3089; // @[Cat.scala 30:58:@22094.4]
  wire [10:0] _T_3091; // @[Cat.scala 30:58:@22096.4]
  wire [10:0] _T_3093; // @[Cat.scala 30:58:@22098.4]
  wire [10:0] _T_3095; // @[Cat.scala 30:58:@22100.4]
  wire [10:0] _T_3097; // @[Cat.scala 30:58:@22102.4]
  wire [10:0] _T_3099; // @[Cat.scala 30:58:@22104.4]
  wire [10:0] _T_3100; // @[Mux.scala 31:69:@22105.4]
  wire [10:0] _T_3101; // @[Mux.scala 31:69:@22106.4]
  wire [10:0] _T_3102; // @[Mux.scala 31:69:@22107.4]
  wire [10:0] _T_3103; // @[Mux.scala 31:69:@22108.4]
  wire [10:0] _T_3104; // @[Mux.scala 31:69:@22109.4]
  wire [10:0] _T_3105; // @[Mux.scala 31:69:@22110.4]
  wire [10:0] _T_3106; // @[Mux.scala 31:69:@22111.4]
  wire [10:0] _T_3107; // @[Mux.scala 31:69:@22112.4]
  wire  _T_3115; // @[MemPrimitives.scala 110:228:@22121.4]
  wire  _T_3121; // @[MemPrimitives.scala 110:228:@22125.4]
  wire  _T_3127; // @[MemPrimitives.scala 110:228:@22129.4]
  wire  _T_3133; // @[MemPrimitives.scala 110:228:@22133.4]
  wire  _T_3139; // @[MemPrimitives.scala 110:228:@22137.4]
  wire  _T_3145; // @[MemPrimitives.scala 110:228:@22141.4]
  wire  _T_3151; // @[MemPrimitives.scala 110:228:@22145.4]
  wire  _T_3157; // @[MemPrimitives.scala 110:228:@22149.4]
  wire  _T_3163; // @[MemPrimitives.scala 110:228:@22153.4]
  wire  _T_3165; // @[MemPrimitives.scala 126:35:@22167.4]
  wire  _T_3166; // @[MemPrimitives.scala 126:35:@22168.4]
  wire  _T_3167; // @[MemPrimitives.scala 126:35:@22169.4]
  wire  _T_3168; // @[MemPrimitives.scala 126:35:@22170.4]
  wire  _T_3169; // @[MemPrimitives.scala 126:35:@22171.4]
  wire  _T_3170; // @[MemPrimitives.scala 126:35:@22172.4]
  wire  _T_3171; // @[MemPrimitives.scala 126:35:@22173.4]
  wire  _T_3172; // @[MemPrimitives.scala 126:35:@22174.4]
  wire  _T_3173; // @[MemPrimitives.scala 126:35:@22175.4]
  wire [10:0] _T_3175; // @[Cat.scala 30:58:@22177.4]
  wire [10:0] _T_3177; // @[Cat.scala 30:58:@22179.4]
  wire [10:0] _T_3179; // @[Cat.scala 30:58:@22181.4]
  wire [10:0] _T_3181; // @[Cat.scala 30:58:@22183.4]
  wire [10:0] _T_3183; // @[Cat.scala 30:58:@22185.4]
  wire [10:0] _T_3185; // @[Cat.scala 30:58:@22187.4]
  wire [10:0] _T_3187; // @[Cat.scala 30:58:@22189.4]
  wire [10:0] _T_3189; // @[Cat.scala 30:58:@22191.4]
  wire [10:0] _T_3191; // @[Cat.scala 30:58:@22193.4]
  wire [10:0] _T_3192; // @[Mux.scala 31:69:@22194.4]
  wire [10:0] _T_3193; // @[Mux.scala 31:69:@22195.4]
  wire [10:0] _T_3194; // @[Mux.scala 31:69:@22196.4]
  wire [10:0] _T_3195; // @[Mux.scala 31:69:@22197.4]
  wire [10:0] _T_3196; // @[Mux.scala 31:69:@22198.4]
  wire [10:0] _T_3197; // @[Mux.scala 31:69:@22199.4]
  wire [10:0] _T_3198; // @[Mux.scala 31:69:@22200.4]
  wire [10:0] _T_3199; // @[Mux.scala 31:69:@22201.4]
  wire  _T_3207; // @[MemPrimitives.scala 110:228:@22210.4]
  wire  _T_3213; // @[MemPrimitives.scala 110:228:@22214.4]
  wire  _T_3219; // @[MemPrimitives.scala 110:228:@22218.4]
  wire  _T_3225; // @[MemPrimitives.scala 110:228:@22222.4]
  wire  _T_3231; // @[MemPrimitives.scala 110:228:@22226.4]
  wire  _T_3237; // @[MemPrimitives.scala 110:228:@22230.4]
  wire  _T_3243; // @[MemPrimitives.scala 110:228:@22234.4]
  wire  _T_3249; // @[MemPrimitives.scala 110:228:@22238.4]
  wire  _T_3255; // @[MemPrimitives.scala 110:228:@22242.4]
  wire  _T_3257; // @[MemPrimitives.scala 126:35:@22256.4]
  wire  _T_3258; // @[MemPrimitives.scala 126:35:@22257.4]
  wire  _T_3259; // @[MemPrimitives.scala 126:35:@22258.4]
  wire  _T_3260; // @[MemPrimitives.scala 126:35:@22259.4]
  wire  _T_3261; // @[MemPrimitives.scala 126:35:@22260.4]
  wire  _T_3262; // @[MemPrimitives.scala 126:35:@22261.4]
  wire  _T_3263; // @[MemPrimitives.scala 126:35:@22262.4]
  wire  _T_3264; // @[MemPrimitives.scala 126:35:@22263.4]
  wire  _T_3265; // @[MemPrimitives.scala 126:35:@22264.4]
  wire [10:0] _T_3267; // @[Cat.scala 30:58:@22266.4]
  wire [10:0] _T_3269; // @[Cat.scala 30:58:@22268.4]
  wire [10:0] _T_3271; // @[Cat.scala 30:58:@22270.4]
  wire [10:0] _T_3273; // @[Cat.scala 30:58:@22272.4]
  wire [10:0] _T_3275; // @[Cat.scala 30:58:@22274.4]
  wire [10:0] _T_3277; // @[Cat.scala 30:58:@22276.4]
  wire [10:0] _T_3279; // @[Cat.scala 30:58:@22278.4]
  wire [10:0] _T_3281; // @[Cat.scala 30:58:@22280.4]
  wire [10:0] _T_3283; // @[Cat.scala 30:58:@22282.4]
  wire [10:0] _T_3284; // @[Mux.scala 31:69:@22283.4]
  wire [10:0] _T_3285; // @[Mux.scala 31:69:@22284.4]
  wire [10:0] _T_3286; // @[Mux.scala 31:69:@22285.4]
  wire [10:0] _T_3287; // @[Mux.scala 31:69:@22286.4]
  wire [10:0] _T_3288; // @[Mux.scala 31:69:@22287.4]
  wire [10:0] _T_3289; // @[Mux.scala 31:69:@22288.4]
  wire [10:0] _T_3290; // @[Mux.scala 31:69:@22289.4]
  wire [10:0] _T_3291; // @[Mux.scala 31:69:@22290.4]
  wire  _T_3299; // @[MemPrimitives.scala 110:228:@22299.4]
  wire  _T_3305; // @[MemPrimitives.scala 110:228:@22303.4]
  wire  _T_3311; // @[MemPrimitives.scala 110:228:@22307.4]
  wire  _T_3317; // @[MemPrimitives.scala 110:228:@22311.4]
  wire  _T_3323; // @[MemPrimitives.scala 110:228:@22315.4]
  wire  _T_3329; // @[MemPrimitives.scala 110:228:@22319.4]
  wire  _T_3335; // @[MemPrimitives.scala 110:228:@22323.4]
  wire  _T_3341; // @[MemPrimitives.scala 110:228:@22327.4]
  wire  _T_3347; // @[MemPrimitives.scala 110:228:@22331.4]
  wire  _T_3349; // @[MemPrimitives.scala 126:35:@22345.4]
  wire  _T_3350; // @[MemPrimitives.scala 126:35:@22346.4]
  wire  _T_3351; // @[MemPrimitives.scala 126:35:@22347.4]
  wire  _T_3352; // @[MemPrimitives.scala 126:35:@22348.4]
  wire  _T_3353; // @[MemPrimitives.scala 126:35:@22349.4]
  wire  _T_3354; // @[MemPrimitives.scala 126:35:@22350.4]
  wire  _T_3355; // @[MemPrimitives.scala 126:35:@22351.4]
  wire  _T_3356; // @[MemPrimitives.scala 126:35:@22352.4]
  wire  _T_3357; // @[MemPrimitives.scala 126:35:@22353.4]
  wire [10:0] _T_3359; // @[Cat.scala 30:58:@22355.4]
  wire [10:0] _T_3361; // @[Cat.scala 30:58:@22357.4]
  wire [10:0] _T_3363; // @[Cat.scala 30:58:@22359.4]
  wire [10:0] _T_3365; // @[Cat.scala 30:58:@22361.4]
  wire [10:0] _T_3367; // @[Cat.scala 30:58:@22363.4]
  wire [10:0] _T_3369; // @[Cat.scala 30:58:@22365.4]
  wire [10:0] _T_3371; // @[Cat.scala 30:58:@22367.4]
  wire [10:0] _T_3373; // @[Cat.scala 30:58:@22369.4]
  wire [10:0] _T_3375; // @[Cat.scala 30:58:@22371.4]
  wire [10:0] _T_3376; // @[Mux.scala 31:69:@22372.4]
  wire [10:0] _T_3377; // @[Mux.scala 31:69:@22373.4]
  wire [10:0] _T_3378; // @[Mux.scala 31:69:@22374.4]
  wire [10:0] _T_3379; // @[Mux.scala 31:69:@22375.4]
  wire [10:0] _T_3380; // @[Mux.scala 31:69:@22376.4]
  wire [10:0] _T_3381; // @[Mux.scala 31:69:@22377.4]
  wire [10:0] _T_3382; // @[Mux.scala 31:69:@22378.4]
  wire [10:0] _T_3383; // @[Mux.scala 31:69:@22379.4]
  wire  _T_3479; // @[package.scala 96:25:@22508.4 package.scala 96:25:@22509.4]
  wire [31:0] _T_3483; // @[Mux.scala 31:69:@22518.4]
  wire  _T_3476; // @[package.scala 96:25:@22500.4 package.scala 96:25:@22501.4]
  wire [31:0] _T_3484; // @[Mux.scala 31:69:@22519.4]
  wire  _T_3473; // @[package.scala 96:25:@22492.4 package.scala 96:25:@22493.4]
  wire [31:0] _T_3485; // @[Mux.scala 31:69:@22520.4]
  wire  _T_3470; // @[package.scala 96:25:@22484.4 package.scala 96:25:@22485.4]
  wire [31:0] _T_3486; // @[Mux.scala 31:69:@22521.4]
  wire  _T_3467; // @[package.scala 96:25:@22476.4 package.scala 96:25:@22477.4]
  wire [31:0] _T_3487; // @[Mux.scala 31:69:@22522.4]
  wire  _T_3464; // @[package.scala 96:25:@22468.4 package.scala 96:25:@22469.4]
  wire [31:0] _T_3488; // @[Mux.scala 31:69:@22523.4]
  wire  _T_3461; // @[package.scala 96:25:@22460.4 package.scala 96:25:@22461.4]
  wire [31:0] _T_3489; // @[Mux.scala 31:69:@22524.4]
  wire  _T_3458; // @[package.scala 96:25:@22452.4 package.scala 96:25:@22453.4]
  wire [31:0] _T_3490; // @[Mux.scala 31:69:@22525.4]
  wire  _T_3455; // @[package.scala 96:25:@22444.4 package.scala 96:25:@22445.4]
  wire [31:0] _T_3491; // @[Mux.scala 31:69:@22526.4]
  wire  _T_3452; // @[package.scala 96:25:@22436.4 package.scala 96:25:@22437.4]
  wire [31:0] _T_3492; // @[Mux.scala 31:69:@22527.4]
  wire  _T_3449; // @[package.scala 96:25:@22428.4 package.scala 96:25:@22429.4]
  wire  _T_3586; // @[package.scala 96:25:@22652.4 package.scala 96:25:@22653.4]
  wire [31:0] _T_3590; // @[Mux.scala 31:69:@22662.4]
  wire  _T_3583; // @[package.scala 96:25:@22644.4 package.scala 96:25:@22645.4]
  wire [31:0] _T_3591; // @[Mux.scala 31:69:@22663.4]
  wire  _T_3580; // @[package.scala 96:25:@22636.4 package.scala 96:25:@22637.4]
  wire [31:0] _T_3592; // @[Mux.scala 31:69:@22664.4]
  wire  _T_3577; // @[package.scala 96:25:@22628.4 package.scala 96:25:@22629.4]
  wire [31:0] _T_3593; // @[Mux.scala 31:69:@22665.4]
  wire  _T_3574; // @[package.scala 96:25:@22620.4 package.scala 96:25:@22621.4]
  wire [31:0] _T_3594; // @[Mux.scala 31:69:@22666.4]
  wire  _T_3571; // @[package.scala 96:25:@22612.4 package.scala 96:25:@22613.4]
  wire [31:0] _T_3595; // @[Mux.scala 31:69:@22667.4]
  wire  _T_3568; // @[package.scala 96:25:@22604.4 package.scala 96:25:@22605.4]
  wire [31:0] _T_3596; // @[Mux.scala 31:69:@22668.4]
  wire  _T_3565; // @[package.scala 96:25:@22596.4 package.scala 96:25:@22597.4]
  wire [31:0] _T_3597; // @[Mux.scala 31:69:@22669.4]
  wire  _T_3562; // @[package.scala 96:25:@22588.4 package.scala 96:25:@22589.4]
  wire [31:0] _T_3598; // @[Mux.scala 31:69:@22670.4]
  wire  _T_3559; // @[package.scala 96:25:@22580.4 package.scala 96:25:@22581.4]
  wire [31:0] _T_3599; // @[Mux.scala 31:69:@22671.4]
  wire  _T_3556; // @[package.scala 96:25:@22572.4 package.scala 96:25:@22573.4]
  wire  _T_3693; // @[package.scala 96:25:@22796.4 package.scala 96:25:@22797.4]
  wire [31:0] _T_3697; // @[Mux.scala 31:69:@22806.4]
  wire  _T_3690; // @[package.scala 96:25:@22788.4 package.scala 96:25:@22789.4]
  wire [31:0] _T_3698; // @[Mux.scala 31:69:@22807.4]
  wire  _T_3687; // @[package.scala 96:25:@22780.4 package.scala 96:25:@22781.4]
  wire [31:0] _T_3699; // @[Mux.scala 31:69:@22808.4]
  wire  _T_3684; // @[package.scala 96:25:@22772.4 package.scala 96:25:@22773.4]
  wire [31:0] _T_3700; // @[Mux.scala 31:69:@22809.4]
  wire  _T_3681; // @[package.scala 96:25:@22764.4 package.scala 96:25:@22765.4]
  wire [31:0] _T_3701; // @[Mux.scala 31:69:@22810.4]
  wire  _T_3678; // @[package.scala 96:25:@22756.4 package.scala 96:25:@22757.4]
  wire [31:0] _T_3702; // @[Mux.scala 31:69:@22811.4]
  wire  _T_3675; // @[package.scala 96:25:@22748.4 package.scala 96:25:@22749.4]
  wire [31:0] _T_3703; // @[Mux.scala 31:69:@22812.4]
  wire  _T_3672; // @[package.scala 96:25:@22740.4 package.scala 96:25:@22741.4]
  wire [31:0] _T_3704; // @[Mux.scala 31:69:@22813.4]
  wire  _T_3669; // @[package.scala 96:25:@22732.4 package.scala 96:25:@22733.4]
  wire [31:0] _T_3705; // @[Mux.scala 31:69:@22814.4]
  wire  _T_3666; // @[package.scala 96:25:@22724.4 package.scala 96:25:@22725.4]
  wire [31:0] _T_3706; // @[Mux.scala 31:69:@22815.4]
  wire  _T_3663; // @[package.scala 96:25:@22716.4 package.scala 96:25:@22717.4]
  wire  _T_3800; // @[package.scala 96:25:@22940.4 package.scala 96:25:@22941.4]
  wire [31:0] _T_3804; // @[Mux.scala 31:69:@22950.4]
  wire  _T_3797; // @[package.scala 96:25:@22932.4 package.scala 96:25:@22933.4]
  wire [31:0] _T_3805; // @[Mux.scala 31:69:@22951.4]
  wire  _T_3794; // @[package.scala 96:25:@22924.4 package.scala 96:25:@22925.4]
  wire [31:0] _T_3806; // @[Mux.scala 31:69:@22952.4]
  wire  _T_3791; // @[package.scala 96:25:@22916.4 package.scala 96:25:@22917.4]
  wire [31:0] _T_3807; // @[Mux.scala 31:69:@22953.4]
  wire  _T_3788; // @[package.scala 96:25:@22908.4 package.scala 96:25:@22909.4]
  wire [31:0] _T_3808; // @[Mux.scala 31:69:@22954.4]
  wire  _T_3785; // @[package.scala 96:25:@22900.4 package.scala 96:25:@22901.4]
  wire [31:0] _T_3809; // @[Mux.scala 31:69:@22955.4]
  wire  _T_3782; // @[package.scala 96:25:@22892.4 package.scala 96:25:@22893.4]
  wire [31:0] _T_3810; // @[Mux.scala 31:69:@22956.4]
  wire  _T_3779; // @[package.scala 96:25:@22884.4 package.scala 96:25:@22885.4]
  wire [31:0] _T_3811; // @[Mux.scala 31:69:@22957.4]
  wire  _T_3776; // @[package.scala 96:25:@22876.4 package.scala 96:25:@22877.4]
  wire [31:0] _T_3812; // @[Mux.scala 31:69:@22958.4]
  wire  _T_3773; // @[package.scala 96:25:@22868.4 package.scala 96:25:@22869.4]
  wire [31:0] _T_3813; // @[Mux.scala 31:69:@22959.4]
  wire  _T_3770; // @[package.scala 96:25:@22860.4 package.scala 96:25:@22861.4]
  wire  _T_3907; // @[package.scala 96:25:@23084.4 package.scala 96:25:@23085.4]
  wire [31:0] _T_3911; // @[Mux.scala 31:69:@23094.4]
  wire  _T_3904; // @[package.scala 96:25:@23076.4 package.scala 96:25:@23077.4]
  wire [31:0] _T_3912; // @[Mux.scala 31:69:@23095.4]
  wire  _T_3901; // @[package.scala 96:25:@23068.4 package.scala 96:25:@23069.4]
  wire [31:0] _T_3913; // @[Mux.scala 31:69:@23096.4]
  wire  _T_3898; // @[package.scala 96:25:@23060.4 package.scala 96:25:@23061.4]
  wire [31:0] _T_3914; // @[Mux.scala 31:69:@23097.4]
  wire  _T_3895; // @[package.scala 96:25:@23052.4 package.scala 96:25:@23053.4]
  wire [31:0] _T_3915; // @[Mux.scala 31:69:@23098.4]
  wire  _T_3892; // @[package.scala 96:25:@23044.4 package.scala 96:25:@23045.4]
  wire [31:0] _T_3916; // @[Mux.scala 31:69:@23099.4]
  wire  _T_3889; // @[package.scala 96:25:@23036.4 package.scala 96:25:@23037.4]
  wire [31:0] _T_3917; // @[Mux.scala 31:69:@23100.4]
  wire  _T_3886; // @[package.scala 96:25:@23028.4 package.scala 96:25:@23029.4]
  wire [31:0] _T_3918; // @[Mux.scala 31:69:@23101.4]
  wire  _T_3883; // @[package.scala 96:25:@23020.4 package.scala 96:25:@23021.4]
  wire [31:0] _T_3919; // @[Mux.scala 31:69:@23102.4]
  wire  _T_3880; // @[package.scala 96:25:@23012.4 package.scala 96:25:@23013.4]
  wire [31:0] _T_3920; // @[Mux.scala 31:69:@23103.4]
  wire  _T_3877; // @[package.scala 96:25:@23004.4 package.scala 96:25:@23005.4]
  wire  _T_4014; // @[package.scala 96:25:@23228.4 package.scala 96:25:@23229.4]
  wire [31:0] _T_4018; // @[Mux.scala 31:69:@23238.4]
  wire  _T_4011; // @[package.scala 96:25:@23220.4 package.scala 96:25:@23221.4]
  wire [31:0] _T_4019; // @[Mux.scala 31:69:@23239.4]
  wire  _T_4008; // @[package.scala 96:25:@23212.4 package.scala 96:25:@23213.4]
  wire [31:0] _T_4020; // @[Mux.scala 31:69:@23240.4]
  wire  _T_4005; // @[package.scala 96:25:@23204.4 package.scala 96:25:@23205.4]
  wire [31:0] _T_4021; // @[Mux.scala 31:69:@23241.4]
  wire  _T_4002; // @[package.scala 96:25:@23196.4 package.scala 96:25:@23197.4]
  wire [31:0] _T_4022; // @[Mux.scala 31:69:@23242.4]
  wire  _T_3999; // @[package.scala 96:25:@23188.4 package.scala 96:25:@23189.4]
  wire [31:0] _T_4023; // @[Mux.scala 31:69:@23243.4]
  wire  _T_3996; // @[package.scala 96:25:@23180.4 package.scala 96:25:@23181.4]
  wire [31:0] _T_4024; // @[Mux.scala 31:69:@23244.4]
  wire  _T_3993; // @[package.scala 96:25:@23172.4 package.scala 96:25:@23173.4]
  wire [31:0] _T_4025; // @[Mux.scala 31:69:@23245.4]
  wire  _T_3990; // @[package.scala 96:25:@23164.4 package.scala 96:25:@23165.4]
  wire [31:0] _T_4026; // @[Mux.scala 31:69:@23246.4]
  wire  _T_3987; // @[package.scala 96:25:@23156.4 package.scala 96:25:@23157.4]
  wire [31:0] _T_4027; // @[Mux.scala 31:69:@23247.4]
  wire  _T_3984; // @[package.scala 96:25:@23148.4 package.scala 96:25:@23149.4]
  wire  _T_4121; // @[package.scala 96:25:@23372.4 package.scala 96:25:@23373.4]
  wire [31:0] _T_4125; // @[Mux.scala 31:69:@23382.4]
  wire  _T_4118; // @[package.scala 96:25:@23364.4 package.scala 96:25:@23365.4]
  wire [31:0] _T_4126; // @[Mux.scala 31:69:@23383.4]
  wire  _T_4115; // @[package.scala 96:25:@23356.4 package.scala 96:25:@23357.4]
  wire [31:0] _T_4127; // @[Mux.scala 31:69:@23384.4]
  wire  _T_4112; // @[package.scala 96:25:@23348.4 package.scala 96:25:@23349.4]
  wire [31:0] _T_4128; // @[Mux.scala 31:69:@23385.4]
  wire  _T_4109; // @[package.scala 96:25:@23340.4 package.scala 96:25:@23341.4]
  wire [31:0] _T_4129; // @[Mux.scala 31:69:@23386.4]
  wire  _T_4106; // @[package.scala 96:25:@23332.4 package.scala 96:25:@23333.4]
  wire [31:0] _T_4130; // @[Mux.scala 31:69:@23387.4]
  wire  _T_4103; // @[package.scala 96:25:@23324.4 package.scala 96:25:@23325.4]
  wire [31:0] _T_4131; // @[Mux.scala 31:69:@23388.4]
  wire  _T_4100; // @[package.scala 96:25:@23316.4 package.scala 96:25:@23317.4]
  wire [31:0] _T_4132; // @[Mux.scala 31:69:@23389.4]
  wire  _T_4097; // @[package.scala 96:25:@23308.4 package.scala 96:25:@23309.4]
  wire [31:0] _T_4133; // @[Mux.scala 31:69:@23390.4]
  wire  _T_4094; // @[package.scala 96:25:@23300.4 package.scala 96:25:@23301.4]
  wire [31:0] _T_4134; // @[Mux.scala 31:69:@23391.4]
  wire  _T_4091; // @[package.scala 96:25:@23292.4 package.scala 96:25:@23293.4]
  wire  _T_4228; // @[package.scala 96:25:@23516.4 package.scala 96:25:@23517.4]
  wire [31:0] _T_4232; // @[Mux.scala 31:69:@23526.4]
  wire  _T_4225; // @[package.scala 96:25:@23508.4 package.scala 96:25:@23509.4]
  wire [31:0] _T_4233; // @[Mux.scala 31:69:@23527.4]
  wire  _T_4222; // @[package.scala 96:25:@23500.4 package.scala 96:25:@23501.4]
  wire [31:0] _T_4234; // @[Mux.scala 31:69:@23528.4]
  wire  _T_4219; // @[package.scala 96:25:@23492.4 package.scala 96:25:@23493.4]
  wire [31:0] _T_4235; // @[Mux.scala 31:69:@23529.4]
  wire  _T_4216; // @[package.scala 96:25:@23484.4 package.scala 96:25:@23485.4]
  wire [31:0] _T_4236; // @[Mux.scala 31:69:@23530.4]
  wire  _T_4213; // @[package.scala 96:25:@23476.4 package.scala 96:25:@23477.4]
  wire [31:0] _T_4237; // @[Mux.scala 31:69:@23531.4]
  wire  _T_4210; // @[package.scala 96:25:@23468.4 package.scala 96:25:@23469.4]
  wire [31:0] _T_4238; // @[Mux.scala 31:69:@23532.4]
  wire  _T_4207; // @[package.scala 96:25:@23460.4 package.scala 96:25:@23461.4]
  wire [31:0] _T_4239; // @[Mux.scala 31:69:@23533.4]
  wire  _T_4204; // @[package.scala 96:25:@23452.4 package.scala 96:25:@23453.4]
  wire [31:0] _T_4240; // @[Mux.scala 31:69:@23534.4]
  wire  _T_4201; // @[package.scala 96:25:@23444.4 package.scala 96:25:@23445.4]
  wire [31:0] _T_4241; // @[Mux.scala 31:69:@23535.4]
  wire  _T_4198; // @[package.scala 96:25:@23436.4 package.scala 96:25:@23437.4]
  wire  _T_4335; // @[package.scala 96:25:@23660.4 package.scala 96:25:@23661.4]
  wire [31:0] _T_4339; // @[Mux.scala 31:69:@23670.4]
  wire  _T_4332; // @[package.scala 96:25:@23652.4 package.scala 96:25:@23653.4]
  wire [31:0] _T_4340; // @[Mux.scala 31:69:@23671.4]
  wire  _T_4329; // @[package.scala 96:25:@23644.4 package.scala 96:25:@23645.4]
  wire [31:0] _T_4341; // @[Mux.scala 31:69:@23672.4]
  wire  _T_4326; // @[package.scala 96:25:@23636.4 package.scala 96:25:@23637.4]
  wire [31:0] _T_4342; // @[Mux.scala 31:69:@23673.4]
  wire  _T_4323; // @[package.scala 96:25:@23628.4 package.scala 96:25:@23629.4]
  wire [31:0] _T_4343; // @[Mux.scala 31:69:@23674.4]
  wire  _T_4320; // @[package.scala 96:25:@23620.4 package.scala 96:25:@23621.4]
  wire [31:0] _T_4344; // @[Mux.scala 31:69:@23675.4]
  wire  _T_4317; // @[package.scala 96:25:@23612.4 package.scala 96:25:@23613.4]
  wire [31:0] _T_4345; // @[Mux.scala 31:69:@23676.4]
  wire  _T_4314; // @[package.scala 96:25:@23604.4 package.scala 96:25:@23605.4]
  wire [31:0] _T_4346; // @[Mux.scala 31:69:@23677.4]
  wire  _T_4311; // @[package.scala 96:25:@23596.4 package.scala 96:25:@23597.4]
  wire [31:0] _T_4347; // @[Mux.scala 31:69:@23678.4]
  wire  _T_4308; // @[package.scala 96:25:@23588.4 package.scala 96:25:@23589.4]
  wire [31:0] _T_4348; // @[Mux.scala 31:69:@23679.4]
  wire  _T_4305; // @[package.scala 96:25:@23580.4 package.scala 96:25:@23581.4]
  wire  _T_4442; // @[package.scala 96:25:@23804.4 package.scala 96:25:@23805.4]
  wire [31:0] _T_4446; // @[Mux.scala 31:69:@23814.4]
  wire  _T_4439; // @[package.scala 96:25:@23796.4 package.scala 96:25:@23797.4]
  wire [31:0] _T_4447; // @[Mux.scala 31:69:@23815.4]
  wire  _T_4436; // @[package.scala 96:25:@23788.4 package.scala 96:25:@23789.4]
  wire [31:0] _T_4448; // @[Mux.scala 31:69:@23816.4]
  wire  _T_4433; // @[package.scala 96:25:@23780.4 package.scala 96:25:@23781.4]
  wire [31:0] _T_4449; // @[Mux.scala 31:69:@23817.4]
  wire  _T_4430; // @[package.scala 96:25:@23772.4 package.scala 96:25:@23773.4]
  wire [31:0] _T_4450; // @[Mux.scala 31:69:@23818.4]
  wire  _T_4427; // @[package.scala 96:25:@23764.4 package.scala 96:25:@23765.4]
  wire [31:0] _T_4451; // @[Mux.scala 31:69:@23819.4]
  wire  _T_4424; // @[package.scala 96:25:@23756.4 package.scala 96:25:@23757.4]
  wire [31:0] _T_4452; // @[Mux.scala 31:69:@23820.4]
  wire  _T_4421; // @[package.scala 96:25:@23748.4 package.scala 96:25:@23749.4]
  wire [31:0] _T_4453; // @[Mux.scala 31:69:@23821.4]
  wire  _T_4418; // @[package.scala 96:25:@23740.4 package.scala 96:25:@23741.4]
  wire [31:0] _T_4454; // @[Mux.scala 31:69:@23822.4]
  wire  _T_4415; // @[package.scala 96:25:@23732.4 package.scala 96:25:@23733.4]
  wire [31:0] _T_4455; // @[Mux.scala 31:69:@23823.4]
  wire  _T_4412; // @[package.scala 96:25:@23724.4 package.scala 96:25:@23725.4]
  wire  _T_4549; // @[package.scala 96:25:@23948.4 package.scala 96:25:@23949.4]
  wire [31:0] _T_4553; // @[Mux.scala 31:69:@23958.4]
  wire  _T_4546; // @[package.scala 96:25:@23940.4 package.scala 96:25:@23941.4]
  wire [31:0] _T_4554; // @[Mux.scala 31:69:@23959.4]
  wire  _T_4543; // @[package.scala 96:25:@23932.4 package.scala 96:25:@23933.4]
  wire [31:0] _T_4555; // @[Mux.scala 31:69:@23960.4]
  wire  _T_4540; // @[package.scala 96:25:@23924.4 package.scala 96:25:@23925.4]
  wire [31:0] _T_4556; // @[Mux.scala 31:69:@23961.4]
  wire  _T_4537; // @[package.scala 96:25:@23916.4 package.scala 96:25:@23917.4]
  wire [31:0] _T_4557; // @[Mux.scala 31:69:@23962.4]
  wire  _T_4534; // @[package.scala 96:25:@23908.4 package.scala 96:25:@23909.4]
  wire [31:0] _T_4558; // @[Mux.scala 31:69:@23963.4]
  wire  _T_4531; // @[package.scala 96:25:@23900.4 package.scala 96:25:@23901.4]
  wire [31:0] _T_4559; // @[Mux.scala 31:69:@23964.4]
  wire  _T_4528; // @[package.scala 96:25:@23892.4 package.scala 96:25:@23893.4]
  wire [31:0] _T_4560; // @[Mux.scala 31:69:@23965.4]
  wire  _T_4525; // @[package.scala 96:25:@23884.4 package.scala 96:25:@23885.4]
  wire [31:0] _T_4561; // @[Mux.scala 31:69:@23966.4]
  wire  _T_4522; // @[package.scala 96:25:@23876.4 package.scala 96:25:@23877.4]
  wire [31:0] _T_4562; // @[Mux.scala 31:69:@23967.4]
  wire  _T_4519; // @[package.scala 96:25:@23868.4 package.scala 96:25:@23869.4]
  wire  _T_4656; // @[package.scala 96:25:@24092.4 package.scala 96:25:@24093.4]
  wire [31:0] _T_4660; // @[Mux.scala 31:69:@24102.4]
  wire  _T_4653; // @[package.scala 96:25:@24084.4 package.scala 96:25:@24085.4]
  wire [31:0] _T_4661; // @[Mux.scala 31:69:@24103.4]
  wire  _T_4650; // @[package.scala 96:25:@24076.4 package.scala 96:25:@24077.4]
  wire [31:0] _T_4662; // @[Mux.scala 31:69:@24104.4]
  wire  _T_4647; // @[package.scala 96:25:@24068.4 package.scala 96:25:@24069.4]
  wire [31:0] _T_4663; // @[Mux.scala 31:69:@24105.4]
  wire  _T_4644; // @[package.scala 96:25:@24060.4 package.scala 96:25:@24061.4]
  wire [31:0] _T_4664; // @[Mux.scala 31:69:@24106.4]
  wire  _T_4641; // @[package.scala 96:25:@24052.4 package.scala 96:25:@24053.4]
  wire [31:0] _T_4665; // @[Mux.scala 31:69:@24107.4]
  wire  _T_4638; // @[package.scala 96:25:@24044.4 package.scala 96:25:@24045.4]
  wire [31:0] _T_4666; // @[Mux.scala 31:69:@24108.4]
  wire  _T_4635; // @[package.scala 96:25:@24036.4 package.scala 96:25:@24037.4]
  wire [31:0] _T_4667; // @[Mux.scala 31:69:@24109.4]
  wire  _T_4632; // @[package.scala 96:25:@24028.4 package.scala 96:25:@24029.4]
  wire [31:0] _T_4668; // @[Mux.scala 31:69:@24110.4]
  wire  _T_4629; // @[package.scala 96:25:@24020.4 package.scala 96:25:@24021.4]
  wire [31:0] _T_4669; // @[Mux.scala 31:69:@24111.4]
  wire  _T_4626; // @[package.scala 96:25:@24012.4 package.scala 96:25:@24013.4]
  wire  _T_4763; // @[package.scala 96:25:@24236.4 package.scala 96:25:@24237.4]
  wire [31:0] _T_4767; // @[Mux.scala 31:69:@24246.4]
  wire  _T_4760; // @[package.scala 96:25:@24228.4 package.scala 96:25:@24229.4]
  wire [31:0] _T_4768; // @[Mux.scala 31:69:@24247.4]
  wire  _T_4757; // @[package.scala 96:25:@24220.4 package.scala 96:25:@24221.4]
  wire [31:0] _T_4769; // @[Mux.scala 31:69:@24248.4]
  wire  _T_4754; // @[package.scala 96:25:@24212.4 package.scala 96:25:@24213.4]
  wire [31:0] _T_4770; // @[Mux.scala 31:69:@24249.4]
  wire  _T_4751; // @[package.scala 96:25:@24204.4 package.scala 96:25:@24205.4]
  wire [31:0] _T_4771; // @[Mux.scala 31:69:@24250.4]
  wire  _T_4748; // @[package.scala 96:25:@24196.4 package.scala 96:25:@24197.4]
  wire [31:0] _T_4772; // @[Mux.scala 31:69:@24251.4]
  wire  _T_4745; // @[package.scala 96:25:@24188.4 package.scala 96:25:@24189.4]
  wire [31:0] _T_4773; // @[Mux.scala 31:69:@24252.4]
  wire  _T_4742; // @[package.scala 96:25:@24180.4 package.scala 96:25:@24181.4]
  wire [31:0] _T_4774; // @[Mux.scala 31:69:@24253.4]
  wire  _T_4739; // @[package.scala 96:25:@24172.4 package.scala 96:25:@24173.4]
  wire [31:0] _T_4775; // @[Mux.scala 31:69:@24254.4]
  wire  _T_4736; // @[package.scala 96:25:@24164.4 package.scala 96:25:@24165.4]
  wire [31:0] _T_4776; // @[Mux.scala 31:69:@24255.4]
  wire  _T_4733; // @[package.scala 96:25:@24156.4 package.scala 96:25:@24157.4]
  wire  _T_4870; // @[package.scala 96:25:@24380.4 package.scala 96:25:@24381.4]
  wire [31:0] _T_4874; // @[Mux.scala 31:69:@24390.4]
  wire  _T_4867; // @[package.scala 96:25:@24372.4 package.scala 96:25:@24373.4]
  wire [31:0] _T_4875; // @[Mux.scala 31:69:@24391.4]
  wire  _T_4864; // @[package.scala 96:25:@24364.4 package.scala 96:25:@24365.4]
  wire [31:0] _T_4876; // @[Mux.scala 31:69:@24392.4]
  wire  _T_4861; // @[package.scala 96:25:@24356.4 package.scala 96:25:@24357.4]
  wire [31:0] _T_4877; // @[Mux.scala 31:69:@24393.4]
  wire  _T_4858; // @[package.scala 96:25:@24348.4 package.scala 96:25:@24349.4]
  wire [31:0] _T_4878; // @[Mux.scala 31:69:@24394.4]
  wire  _T_4855; // @[package.scala 96:25:@24340.4 package.scala 96:25:@24341.4]
  wire [31:0] _T_4879; // @[Mux.scala 31:69:@24395.4]
  wire  _T_4852; // @[package.scala 96:25:@24332.4 package.scala 96:25:@24333.4]
  wire [31:0] _T_4880; // @[Mux.scala 31:69:@24396.4]
  wire  _T_4849; // @[package.scala 96:25:@24324.4 package.scala 96:25:@24325.4]
  wire [31:0] _T_4881; // @[Mux.scala 31:69:@24397.4]
  wire  _T_4846; // @[package.scala 96:25:@24316.4 package.scala 96:25:@24317.4]
  wire [31:0] _T_4882; // @[Mux.scala 31:69:@24398.4]
  wire  _T_4843; // @[package.scala 96:25:@24308.4 package.scala 96:25:@24309.4]
  wire [31:0] _T_4883; // @[Mux.scala 31:69:@24399.4]
  wire  _T_4840; // @[package.scala 96:25:@24300.4 package.scala 96:25:@24301.4]
  wire  _T_4977; // @[package.scala 96:25:@24524.4 package.scala 96:25:@24525.4]
  wire [31:0] _T_4981; // @[Mux.scala 31:69:@24534.4]
  wire  _T_4974; // @[package.scala 96:25:@24516.4 package.scala 96:25:@24517.4]
  wire [31:0] _T_4982; // @[Mux.scala 31:69:@24535.4]
  wire  _T_4971; // @[package.scala 96:25:@24508.4 package.scala 96:25:@24509.4]
  wire [31:0] _T_4983; // @[Mux.scala 31:69:@24536.4]
  wire  _T_4968; // @[package.scala 96:25:@24500.4 package.scala 96:25:@24501.4]
  wire [31:0] _T_4984; // @[Mux.scala 31:69:@24537.4]
  wire  _T_4965; // @[package.scala 96:25:@24492.4 package.scala 96:25:@24493.4]
  wire [31:0] _T_4985; // @[Mux.scala 31:69:@24538.4]
  wire  _T_4962; // @[package.scala 96:25:@24484.4 package.scala 96:25:@24485.4]
  wire [31:0] _T_4986; // @[Mux.scala 31:69:@24539.4]
  wire  _T_4959; // @[package.scala 96:25:@24476.4 package.scala 96:25:@24477.4]
  wire [31:0] _T_4987; // @[Mux.scala 31:69:@24540.4]
  wire  _T_4956; // @[package.scala 96:25:@24468.4 package.scala 96:25:@24469.4]
  wire [31:0] _T_4988; // @[Mux.scala 31:69:@24541.4]
  wire  _T_4953; // @[package.scala 96:25:@24460.4 package.scala 96:25:@24461.4]
  wire [31:0] _T_4989; // @[Mux.scala 31:69:@24542.4]
  wire  _T_4950; // @[package.scala 96:25:@24452.4 package.scala 96:25:@24453.4]
  wire [31:0] _T_4990; // @[Mux.scala 31:69:@24543.4]
  wire  _T_4947; // @[package.scala 96:25:@24444.4 package.scala 96:25:@24445.4]
  wire  _T_5084; // @[package.scala 96:25:@24668.4 package.scala 96:25:@24669.4]
  wire [31:0] _T_5088; // @[Mux.scala 31:69:@24678.4]
  wire  _T_5081; // @[package.scala 96:25:@24660.4 package.scala 96:25:@24661.4]
  wire [31:0] _T_5089; // @[Mux.scala 31:69:@24679.4]
  wire  _T_5078; // @[package.scala 96:25:@24652.4 package.scala 96:25:@24653.4]
  wire [31:0] _T_5090; // @[Mux.scala 31:69:@24680.4]
  wire  _T_5075; // @[package.scala 96:25:@24644.4 package.scala 96:25:@24645.4]
  wire [31:0] _T_5091; // @[Mux.scala 31:69:@24681.4]
  wire  _T_5072; // @[package.scala 96:25:@24636.4 package.scala 96:25:@24637.4]
  wire [31:0] _T_5092; // @[Mux.scala 31:69:@24682.4]
  wire  _T_5069; // @[package.scala 96:25:@24628.4 package.scala 96:25:@24629.4]
  wire [31:0] _T_5093; // @[Mux.scala 31:69:@24683.4]
  wire  _T_5066; // @[package.scala 96:25:@24620.4 package.scala 96:25:@24621.4]
  wire [31:0] _T_5094; // @[Mux.scala 31:69:@24684.4]
  wire  _T_5063; // @[package.scala 96:25:@24612.4 package.scala 96:25:@24613.4]
  wire [31:0] _T_5095; // @[Mux.scala 31:69:@24685.4]
  wire  _T_5060; // @[package.scala 96:25:@24604.4 package.scala 96:25:@24605.4]
  wire [31:0] _T_5096; // @[Mux.scala 31:69:@24686.4]
  wire  _T_5057; // @[package.scala 96:25:@24596.4 package.scala 96:25:@24597.4]
  wire [31:0] _T_5097; // @[Mux.scala 31:69:@24687.4]
  wire  _T_5054; // @[package.scala 96:25:@24588.4 package.scala 96:25:@24589.4]
  wire  _T_5191; // @[package.scala 96:25:@24812.4 package.scala 96:25:@24813.4]
  wire [31:0] _T_5195; // @[Mux.scala 31:69:@24822.4]
  wire  _T_5188; // @[package.scala 96:25:@24804.4 package.scala 96:25:@24805.4]
  wire [31:0] _T_5196; // @[Mux.scala 31:69:@24823.4]
  wire  _T_5185; // @[package.scala 96:25:@24796.4 package.scala 96:25:@24797.4]
  wire [31:0] _T_5197; // @[Mux.scala 31:69:@24824.4]
  wire  _T_5182; // @[package.scala 96:25:@24788.4 package.scala 96:25:@24789.4]
  wire [31:0] _T_5198; // @[Mux.scala 31:69:@24825.4]
  wire  _T_5179; // @[package.scala 96:25:@24780.4 package.scala 96:25:@24781.4]
  wire [31:0] _T_5199; // @[Mux.scala 31:69:@24826.4]
  wire  _T_5176; // @[package.scala 96:25:@24772.4 package.scala 96:25:@24773.4]
  wire [31:0] _T_5200; // @[Mux.scala 31:69:@24827.4]
  wire  _T_5173; // @[package.scala 96:25:@24764.4 package.scala 96:25:@24765.4]
  wire [31:0] _T_5201; // @[Mux.scala 31:69:@24828.4]
  wire  _T_5170; // @[package.scala 96:25:@24756.4 package.scala 96:25:@24757.4]
  wire [31:0] _T_5202; // @[Mux.scala 31:69:@24829.4]
  wire  _T_5167; // @[package.scala 96:25:@24748.4 package.scala 96:25:@24749.4]
  wire [31:0] _T_5203; // @[Mux.scala 31:69:@24830.4]
  wire  _T_5164; // @[package.scala 96:25:@24740.4 package.scala 96:25:@24741.4]
  wire [31:0] _T_5204; // @[Mux.scala 31:69:@24831.4]
  wire  _T_5161; // @[package.scala 96:25:@24732.4 package.scala 96:25:@24733.4]
  wire  _T_5298; // @[package.scala 96:25:@24956.4 package.scala 96:25:@24957.4]
  wire [31:0] _T_5302; // @[Mux.scala 31:69:@24966.4]
  wire  _T_5295; // @[package.scala 96:25:@24948.4 package.scala 96:25:@24949.4]
  wire [31:0] _T_5303; // @[Mux.scala 31:69:@24967.4]
  wire  _T_5292; // @[package.scala 96:25:@24940.4 package.scala 96:25:@24941.4]
  wire [31:0] _T_5304; // @[Mux.scala 31:69:@24968.4]
  wire  _T_5289; // @[package.scala 96:25:@24932.4 package.scala 96:25:@24933.4]
  wire [31:0] _T_5305; // @[Mux.scala 31:69:@24969.4]
  wire  _T_5286; // @[package.scala 96:25:@24924.4 package.scala 96:25:@24925.4]
  wire [31:0] _T_5306; // @[Mux.scala 31:69:@24970.4]
  wire  _T_5283; // @[package.scala 96:25:@24916.4 package.scala 96:25:@24917.4]
  wire [31:0] _T_5307; // @[Mux.scala 31:69:@24971.4]
  wire  _T_5280; // @[package.scala 96:25:@24908.4 package.scala 96:25:@24909.4]
  wire [31:0] _T_5308; // @[Mux.scala 31:69:@24972.4]
  wire  _T_5277; // @[package.scala 96:25:@24900.4 package.scala 96:25:@24901.4]
  wire [31:0] _T_5309; // @[Mux.scala 31:69:@24973.4]
  wire  _T_5274; // @[package.scala 96:25:@24892.4 package.scala 96:25:@24893.4]
  wire [31:0] _T_5310; // @[Mux.scala 31:69:@24974.4]
  wire  _T_5271; // @[package.scala 96:25:@24884.4 package.scala 96:25:@24885.4]
  wire [31:0] _T_5311; // @[Mux.scala 31:69:@24975.4]
  wire  _T_5268; // @[package.scala 96:25:@24876.4 package.scala 96:25:@24877.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@19410.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@19426.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@19442.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@19458.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@19474.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@19490.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@19506.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@19522.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@19538.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@19554.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@19570.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@19586.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@19602.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@19618.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@19634.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@19650.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  Mem1D_5 Mem1D_16 ( // @[MemPrimitives.scala 64:21:@19666.4]
    .clock(Mem1D_16_clock),
    .reset(Mem1D_16_reset),
    .io_r_ofs_0(Mem1D_16_io_r_ofs_0),
    .io_r_backpressure(Mem1D_16_io_r_backpressure),
    .io_w_ofs_0(Mem1D_16_io_w_ofs_0),
    .io_w_data_0(Mem1D_16_io_w_data_0),
    .io_w_en_0(Mem1D_16_io_w_en_0),
    .io_output(Mem1D_16_io_output)
  );
  Mem1D_5 Mem1D_17 ( // @[MemPrimitives.scala 64:21:@19682.4]
    .clock(Mem1D_17_clock),
    .reset(Mem1D_17_reset),
    .io_r_ofs_0(Mem1D_17_io_r_ofs_0),
    .io_r_backpressure(Mem1D_17_io_r_backpressure),
    .io_w_ofs_0(Mem1D_17_io_w_ofs_0),
    .io_w_data_0(Mem1D_17_io_w_data_0),
    .io_w_en_0(Mem1D_17_io_w_en_0),
    .io_output(Mem1D_17_io_output)
  );
  Mem1D_5 Mem1D_18 ( // @[MemPrimitives.scala 64:21:@19698.4]
    .clock(Mem1D_18_clock),
    .reset(Mem1D_18_reset),
    .io_r_ofs_0(Mem1D_18_io_r_ofs_0),
    .io_r_backpressure(Mem1D_18_io_r_backpressure),
    .io_w_ofs_0(Mem1D_18_io_w_ofs_0),
    .io_w_data_0(Mem1D_18_io_w_data_0),
    .io_w_en_0(Mem1D_18_io_w_en_0),
    .io_output(Mem1D_18_io_output)
  );
  Mem1D_5 Mem1D_19 ( // @[MemPrimitives.scala 64:21:@19714.4]
    .clock(Mem1D_19_clock),
    .reset(Mem1D_19_reset),
    .io_r_ofs_0(Mem1D_19_io_r_ofs_0),
    .io_r_backpressure(Mem1D_19_io_r_backpressure),
    .io_w_ofs_0(Mem1D_19_io_w_ofs_0),
    .io_w_data_0(Mem1D_19_io_w_data_0),
    .io_w_en_0(Mem1D_19_io_w_en_0),
    .io_output(Mem1D_19_io_output)
  );
  Mem1D_5 Mem1D_20 ( // @[MemPrimitives.scala 64:21:@19730.4]
    .clock(Mem1D_20_clock),
    .reset(Mem1D_20_reset),
    .io_r_ofs_0(Mem1D_20_io_r_ofs_0),
    .io_r_backpressure(Mem1D_20_io_r_backpressure),
    .io_w_ofs_0(Mem1D_20_io_w_ofs_0),
    .io_w_data_0(Mem1D_20_io_w_data_0),
    .io_w_en_0(Mem1D_20_io_w_en_0),
    .io_output(Mem1D_20_io_output)
  );
  Mem1D_5 Mem1D_21 ( // @[MemPrimitives.scala 64:21:@19746.4]
    .clock(Mem1D_21_clock),
    .reset(Mem1D_21_reset),
    .io_r_ofs_0(Mem1D_21_io_r_ofs_0),
    .io_r_backpressure(Mem1D_21_io_r_backpressure),
    .io_w_ofs_0(Mem1D_21_io_w_ofs_0),
    .io_w_data_0(Mem1D_21_io_w_data_0),
    .io_w_en_0(Mem1D_21_io_w_en_0),
    .io_output(Mem1D_21_io_output)
  );
  Mem1D_5 Mem1D_22 ( // @[MemPrimitives.scala 64:21:@19762.4]
    .clock(Mem1D_22_clock),
    .reset(Mem1D_22_reset),
    .io_r_ofs_0(Mem1D_22_io_r_ofs_0),
    .io_r_backpressure(Mem1D_22_io_r_backpressure),
    .io_w_ofs_0(Mem1D_22_io_w_ofs_0),
    .io_w_data_0(Mem1D_22_io_w_data_0),
    .io_w_en_0(Mem1D_22_io_w_en_0),
    .io_output(Mem1D_22_io_output)
  );
  Mem1D_5 Mem1D_23 ( // @[MemPrimitives.scala 64:21:@19778.4]
    .clock(Mem1D_23_clock),
    .reset(Mem1D_23_reset),
    .io_r_ofs_0(Mem1D_23_io_r_ofs_0),
    .io_r_backpressure(Mem1D_23_io_r_backpressure),
    .io_w_ofs_0(Mem1D_23_io_w_ofs_0),
    .io_w_data_0(Mem1D_23_io_w_data_0),
    .io_w_en_0(Mem1D_23_io_w_en_0),
    .io_output(Mem1D_23_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@20286.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_ins_6(StickySelects_io_ins_6),
    .io_ins_7(StickySelects_io_ins_7),
    .io_ins_8(StickySelects_io_ins_8),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5),
    .io_outs_6(StickySelects_io_outs_6),
    .io_outs_7(StickySelects_io_outs_7),
    .io_outs_8(StickySelects_io_outs_8)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@20375.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_ins_6(StickySelects_1_io_ins_6),
    .io_ins_7(StickySelects_1_io_ins_7),
    .io_ins_8(StickySelects_1_io_ins_8),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5),
    .io_outs_6(StickySelects_1_io_outs_6),
    .io_outs_7(StickySelects_1_io_outs_7),
    .io_outs_8(StickySelects_1_io_outs_8)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@20464.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_ins_6(StickySelects_2_io_ins_6),
    .io_ins_7(StickySelects_2_io_ins_7),
    .io_ins_8(StickySelects_2_io_ins_8),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5),
    .io_outs_6(StickySelects_2_io_outs_6),
    .io_outs_7(StickySelects_2_io_outs_7),
    .io_outs_8(StickySelects_2_io_outs_8)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@20553.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_ins_6(StickySelects_3_io_ins_6),
    .io_ins_7(StickySelects_3_io_ins_7),
    .io_ins_8(StickySelects_3_io_ins_8),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5),
    .io_outs_6(StickySelects_3_io_outs_6),
    .io_outs_7(StickySelects_3_io_outs_7),
    .io_outs_8(StickySelects_3_io_outs_8)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@20642.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_ins_6(StickySelects_4_io_ins_6),
    .io_ins_7(StickySelects_4_io_ins_7),
    .io_ins_8(StickySelects_4_io_ins_8),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5),
    .io_outs_6(StickySelects_4_io_outs_6),
    .io_outs_7(StickySelects_4_io_outs_7),
    .io_outs_8(StickySelects_4_io_outs_8)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@20731.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_ins_6(StickySelects_5_io_ins_6),
    .io_ins_7(StickySelects_5_io_ins_7),
    .io_ins_8(StickySelects_5_io_ins_8),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5),
    .io_outs_6(StickySelects_5_io_outs_6),
    .io_outs_7(StickySelects_5_io_outs_7),
    .io_outs_8(StickySelects_5_io_outs_8)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@20820.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_ins_6(StickySelects_6_io_ins_6),
    .io_ins_7(StickySelects_6_io_ins_7),
    .io_ins_8(StickySelects_6_io_ins_8),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5),
    .io_outs_6(StickySelects_6_io_outs_6),
    .io_outs_7(StickySelects_6_io_outs_7),
    .io_outs_8(StickySelects_6_io_outs_8)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@20909.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_ins_6(StickySelects_7_io_ins_6),
    .io_ins_7(StickySelects_7_io_ins_7),
    .io_ins_8(StickySelects_7_io_ins_8),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5),
    .io_outs_6(StickySelects_7_io_outs_6),
    .io_outs_7(StickySelects_7_io_outs_7),
    .io_outs_8(StickySelects_7_io_outs_8)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@20998.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_ins_6(StickySelects_8_io_ins_6),
    .io_ins_7(StickySelects_8_io_ins_7),
    .io_ins_8(StickySelects_8_io_ins_8),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5),
    .io_outs_6(StickySelects_8_io_outs_6),
    .io_outs_7(StickySelects_8_io_outs_7),
    .io_outs_8(StickySelects_8_io_outs_8)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@21087.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_ins_6(StickySelects_9_io_ins_6),
    .io_ins_7(StickySelects_9_io_ins_7),
    .io_ins_8(StickySelects_9_io_ins_8),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5),
    .io_outs_6(StickySelects_9_io_outs_6),
    .io_outs_7(StickySelects_9_io_outs_7),
    .io_outs_8(StickySelects_9_io_outs_8)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@21176.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_ins_6(StickySelects_10_io_ins_6),
    .io_ins_7(StickySelects_10_io_ins_7),
    .io_ins_8(StickySelects_10_io_ins_8),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5),
    .io_outs_6(StickySelects_10_io_outs_6),
    .io_outs_7(StickySelects_10_io_outs_7),
    .io_outs_8(StickySelects_10_io_outs_8)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@21265.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_ins_6(StickySelects_11_io_ins_6),
    .io_ins_7(StickySelects_11_io_ins_7),
    .io_ins_8(StickySelects_11_io_ins_8),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5),
    .io_outs_6(StickySelects_11_io_outs_6),
    .io_outs_7(StickySelects_11_io_outs_7),
    .io_outs_8(StickySelects_11_io_outs_8)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@21354.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_ins_6(StickySelects_12_io_ins_6),
    .io_ins_7(StickySelects_12_io_ins_7),
    .io_ins_8(StickySelects_12_io_ins_8),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5),
    .io_outs_6(StickySelects_12_io_outs_6),
    .io_outs_7(StickySelects_12_io_outs_7),
    .io_outs_8(StickySelects_12_io_outs_8)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@21443.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_ins_6(StickySelects_13_io_ins_6),
    .io_ins_7(StickySelects_13_io_ins_7),
    .io_ins_8(StickySelects_13_io_ins_8),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5),
    .io_outs_6(StickySelects_13_io_outs_6),
    .io_outs_7(StickySelects_13_io_outs_7),
    .io_outs_8(StickySelects_13_io_outs_8)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@21532.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_ins_6(StickySelects_14_io_ins_6),
    .io_ins_7(StickySelects_14_io_ins_7),
    .io_ins_8(StickySelects_14_io_ins_8),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5),
    .io_outs_6(StickySelects_14_io_outs_6),
    .io_outs_7(StickySelects_14_io_outs_7),
    .io_outs_8(StickySelects_14_io_outs_8)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@21621.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_ins_6(StickySelects_15_io_ins_6),
    .io_ins_7(StickySelects_15_io_ins_7),
    .io_ins_8(StickySelects_15_io_ins_8),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5),
    .io_outs_6(StickySelects_15_io_outs_6),
    .io_outs_7(StickySelects_15_io_outs_7),
    .io_outs_8(StickySelects_15_io_outs_8)
  );
  StickySelects_1 StickySelects_16 ( // @[MemPrimitives.scala 124:33:@21710.4]
    .clock(StickySelects_16_clock),
    .reset(StickySelects_16_reset),
    .io_ins_0(StickySelects_16_io_ins_0),
    .io_ins_1(StickySelects_16_io_ins_1),
    .io_ins_2(StickySelects_16_io_ins_2),
    .io_ins_3(StickySelects_16_io_ins_3),
    .io_ins_4(StickySelects_16_io_ins_4),
    .io_ins_5(StickySelects_16_io_ins_5),
    .io_ins_6(StickySelects_16_io_ins_6),
    .io_ins_7(StickySelects_16_io_ins_7),
    .io_ins_8(StickySelects_16_io_ins_8),
    .io_outs_0(StickySelects_16_io_outs_0),
    .io_outs_1(StickySelects_16_io_outs_1),
    .io_outs_2(StickySelects_16_io_outs_2),
    .io_outs_3(StickySelects_16_io_outs_3),
    .io_outs_4(StickySelects_16_io_outs_4),
    .io_outs_5(StickySelects_16_io_outs_5),
    .io_outs_6(StickySelects_16_io_outs_6),
    .io_outs_7(StickySelects_16_io_outs_7),
    .io_outs_8(StickySelects_16_io_outs_8)
  );
  StickySelects_1 StickySelects_17 ( // @[MemPrimitives.scala 124:33:@21799.4]
    .clock(StickySelects_17_clock),
    .reset(StickySelects_17_reset),
    .io_ins_0(StickySelects_17_io_ins_0),
    .io_ins_1(StickySelects_17_io_ins_1),
    .io_ins_2(StickySelects_17_io_ins_2),
    .io_ins_3(StickySelects_17_io_ins_3),
    .io_ins_4(StickySelects_17_io_ins_4),
    .io_ins_5(StickySelects_17_io_ins_5),
    .io_ins_6(StickySelects_17_io_ins_6),
    .io_ins_7(StickySelects_17_io_ins_7),
    .io_ins_8(StickySelects_17_io_ins_8),
    .io_outs_0(StickySelects_17_io_outs_0),
    .io_outs_1(StickySelects_17_io_outs_1),
    .io_outs_2(StickySelects_17_io_outs_2),
    .io_outs_3(StickySelects_17_io_outs_3),
    .io_outs_4(StickySelects_17_io_outs_4),
    .io_outs_5(StickySelects_17_io_outs_5),
    .io_outs_6(StickySelects_17_io_outs_6),
    .io_outs_7(StickySelects_17_io_outs_7),
    .io_outs_8(StickySelects_17_io_outs_8)
  );
  StickySelects_1 StickySelects_18 ( // @[MemPrimitives.scala 124:33:@21888.4]
    .clock(StickySelects_18_clock),
    .reset(StickySelects_18_reset),
    .io_ins_0(StickySelects_18_io_ins_0),
    .io_ins_1(StickySelects_18_io_ins_1),
    .io_ins_2(StickySelects_18_io_ins_2),
    .io_ins_3(StickySelects_18_io_ins_3),
    .io_ins_4(StickySelects_18_io_ins_4),
    .io_ins_5(StickySelects_18_io_ins_5),
    .io_ins_6(StickySelects_18_io_ins_6),
    .io_ins_7(StickySelects_18_io_ins_7),
    .io_ins_8(StickySelects_18_io_ins_8),
    .io_outs_0(StickySelects_18_io_outs_0),
    .io_outs_1(StickySelects_18_io_outs_1),
    .io_outs_2(StickySelects_18_io_outs_2),
    .io_outs_3(StickySelects_18_io_outs_3),
    .io_outs_4(StickySelects_18_io_outs_4),
    .io_outs_5(StickySelects_18_io_outs_5),
    .io_outs_6(StickySelects_18_io_outs_6),
    .io_outs_7(StickySelects_18_io_outs_7),
    .io_outs_8(StickySelects_18_io_outs_8)
  );
  StickySelects_1 StickySelects_19 ( // @[MemPrimitives.scala 124:33:@21977.4]
    .clock(StickySelects_19_clock),
    .reset(StickySelects_19_reset),
    .io_ins_0(StickySelects_19_io_ins_0),
    .io_ins_1(StickySelects_19_io_ins_1),
    .io_ins_2(StickySelects_19_io_ins_2),
    .io_ins_3(StickySelects_19_io_ins_3),
    .io_ins_4(StickySelects_19_io_ins_4),
    .io_ins_5(StickySelects_19_io_ins_5),
    .io_ins_6(StickySelects_19_io_ins_6),
    .io_ins_7(StickySelects_19_io_ins_7),
    .io_ins_8(StickySelects_19_io_ins_8),
    .io_outs_0(StickySelects_19_io_outs_0),
    .io_outs_1(StickySelects_19_io_outs_1),
    .io_outs_2(StickySelects_19_io_outs_2),
    .io_outs_3(StickySelects_19_io_outs_3),
    .io_outs_4(StickySelects_19_io_outs_4),
    .io_outs_5(StickySelects_19_io_outs_5),
    .io_outs_6(StickySelects_19_io_outs_6),
    .io_outs_7(StickySelects_19_io_outs_7),
    .io_outs_8(StickySelects_19_io_outs_8)
  );
  StickySelects_1 StickySelects_20 ( // @[MemPrimitives.scala 124:33:@22066.4]
    .clock(StickySelects_20_clock),
    .reset(StickySelects_20_reset),
    .io_ins_0(StickySelects_20_io_ins_0),
    .io_ins_1(StickySelects_20_io_ins_1),
    .io_ins_2(StickySelects_20_io_ins_2),
    .io_ins_3(StickySelects_20_io_ins_3),
    .io_ins_4(StickySelects_20_io_ins_4),
    .io_ins_5(StickySelects_20_io_ins_5),
    .io_ins_6(StickySelects_20_io_ins_6),
    .io_ins_7(StickySelects_20_io_ins_7),
    .io_ins_8(StickySelects_20_io_ins_8),
    .io_outs_0(StickySelects_20_io_outs_0),
    .io_outs_1(StickySelects_20_io_outs_1),
    .io_outs_2(StickySelects_20_io_outs_2),
    .io_outs_3(StickySelects_20_io_outs_3),
    .io_outs_4(StickySelects_20_io_outs_4),
    .io_outs_5(StickySelects_20_io_outs_5),
    .io_outs_6(StickySelects_20_io_outs_6),
    .io_outs_7(StickySelects_20_io_outs_7),
    .io_outs_8(StickySelects_20_io_outs_8)
  );
  StickySelects_1 StickySelects_21 ( // @[MemPrimitives.scala 124:33:@22155.4]
    .clock(StickySelects_21_clock),
    .reset(StickySelects_21_reset),
    .io_ins_0(StickySelects_21_io_ins_0),
    .io_ins_1(StickySelects_21_io_ins_1),
    .io_ins_2(StickySelects_21_io_ins_2),
    .io_ins_3(StickySelects_21_io_ins_3),
    .io_ins_4(StickySelects_21_io_ins_4),
    .io_ins_5(StickySelects_21_io_ins_5),
    .io_ins_6(StickySelects_21_io_ins_6),
    .io_ins_7(StickySelects_21_io_ins_7),
    .io_ins_8(StickySelects_21_io_ins_8),
    .io_outs_0(StickySelects_21_io_outs_0),
    .io_outs_1(StickySelects_21_io_outs_1),
    .io_outs_2(StickySelects_21_io_outs_2),
    .io_outs_3(StickySelects_21_io_outs_3),
    .io_outs_4(StickySelects_21_io_outs_4),
    .io_outs_5(StickySelects_21_io_outs_5),
    .io_outs_6(StickySelects_21_io_outs_6),
    .io_outs_7(StickySelects_21_io_outs_7),
    .io_outs_8(StickySelects_21_io_outs_8)
  );
  StickySelects_1 StickySelects_22 ( // @[MemPrimitives.scala 124:33:@22244.4]
    .clock(StickySelects_22_clock),
    .reset(StickySelects_22_reset),
    .io_ins_0(StickySelects_22_io_ins_0),
    .io_ins_1(StickySelects_22_io_ins_1),
    .io_ins_2(StickySelects_22_io_ins_2),
    .io_ins_3(StickySelects_22_io_ins_3),
    .io_ins_4(StickySelects_22_io_ins_4),
    .io_ins_5(StickySelects_22_io_ins_5),
    .io_ins_6(StickySelects_22_io_ins_6),
    .io_ins_7(StickySelects_22_io_ins_7),
    .io_ins_8(StickySelects_22_io_ins_8),
    .io_outs_0(StickySelects_22_io_outs_0),
    .io_outs_1(StickySelects_22_io_outs_1),
    .io_outs_2(StickySelects_22_io_outs_2),
    .io_outs_3(StickySelects_22_io_outs_3),
    .io_outs_4(StickySelects_22_io_outs_4),
    .io_outs_5(StickySelects_22_io_outs_5),
    .io_outs_6(StickySelects_22_io_outs_6),
    .io_outs_7(StickySelects_22_io_outs_7),
    .io_outs_8(StickySelects_22_io_outs_8)
  );
  StickySelects_1 StickySelects_23 ( // @[MemPrimitives.scala 124:33:@22333.4]
    .clock(StickySelects_23_clock),
    .reset(StickySelects_23_reset),
    .io_ins_0(StickySelects_23_io_ins_0),
    .io_ins_1(StickySelects_23_io_ins_1),
    .io_ins_2(StickySelects_23_io_ins_2),
    .io_ins_3(StickySelects_23_io_ins_3),
    .io_ins_4(StickySelects_23_io_ins_4),
    .io_ins_5(StickySelects_23_io_ins_5),
    .io_ins_6(StickySelects_23_io_ins_6),
    .io_ins_7(StickySelects_23_io_ins_7),
    .io_ins_8(StickySelects_23_io_ins_8),
    .io_outs_0(StickySelects_23_io_outs_0),
    .io_outs_1(StickySelects_23_io_outs_1),
    .io_outs_2(StickySelects_23_io_outs_2),
    .io_outs_3(StickySelects_23_io_outs_3),
    .io_outs_4(StickySelects_23_io_outs_4),
    .io_outs_5(StickySelects_23_io_outs_5),
    .io_outs_6(StickySelects_23_io_outs_6),
    .io_outs_7(StickySelects_23_io_outs_7),
    .io_outs_8(StickySelects_23_io_outs_8)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@22423.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@22431.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@22439.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@22447.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@22455.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@22463.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@22471.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@22479.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@22487.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@22495.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@22503.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@22511.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@22567.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@22575.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@22583.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@22591.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@22599.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@22607.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@22615.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@22623.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@22631.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@22639.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@22647.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@22655.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@22711.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@22719.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@22727.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@22735.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@22743.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@22751.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@22759.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@22767.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@22775.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@22783.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@22791.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@22799.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@22855.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@22863.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@22871.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@22879.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@22887.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@22895.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@22903.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@22911.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@22919.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@22927.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@22935.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@22943.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@22999.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@23007.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@23015.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@23023.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@23031.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@23039.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@23047.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@23055.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@23063.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@23071.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@23079.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@23087.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@23143.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@23151.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@23159.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@23167.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@23175.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@23183.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@23191.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@23199.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@23207.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@23215.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@23223.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@23231.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@23287.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@23295.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@23303.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@23311.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@23319.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@23327.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@23335.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@23343.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@23351.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@23359.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@23367.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@23375.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@23431.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@23439.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@23447.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@23455.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@23463.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@23471.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@23479.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@23487.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@23495.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@23503.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@23511.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@23519.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@23575.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@23583.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@23591.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@23599.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@23607.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@23615.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@23623.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@23631.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@23639.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@23647.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@23655.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@23663.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_108 ( // @[package.scala 93:22:@23719.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_109 ( // @[package.scala 93:22:@23727.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_110 ( // @[package.scala 93:22:@23735.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_111 ( // @[package.scala 93:22:@23743.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_112 ( // @[package.scala 93:22:@23751.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_113 ( // @[package.scala 93:22:@23759.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_114 ( // @[package.scala 93:22:@23767.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_115 ( // @[package.scala 93:22:@23775.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_116 ( // @[package.scala 93:22:@23783.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_117 ( // @[package.scala 93:22:@23791.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_118 ( // @[package.scala 93:22:@23799.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_119 ( // @[package.scala 93:22:@23807.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_120 ( // @[package.scala 93:22:@23863.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_121 ( // @[package.scala 93:22:@23871.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_122 ( // @[package.scala 93:22:@23879.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_123 ( // @[package.scala 93:22:@23887.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_124 ( // @[package.scala 93:22:@23895.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_125 ( // @[package.scala 93:22:@23903.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_126 ( // @[package.scala 93:22:@23911.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_127 ( // @[package.scala 93:22:@23919.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_128 ( // @[package.scala 93:22:@23927.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_129 ( // @[package.scala 93:22:@23935.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_130 ( // @[package.scala 93:22:@23943.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_131 ( // @[package.scala 93:22:@23951.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_132 ( // @[package.scala 93:22:@24007.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_133 ( // @[package.scala 93:22:@24015.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_134 ( // @[package.scala 93:22:@24023.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_135 ( // @[package.scala 93:22:@24031.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_136 ( // @[package.scala 93:22:@24039.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_137 ( // @[package.scala 93:22:@24047.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_138 ( // @[package.scala 93:22:@24055.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_139 ( // @[package.scala 93:22:@24063.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_140 ( // @[package.scala 93:22:@24071.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_141 ( // @[package.scala 93:22:@24079.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_142 ( // @[package.scala 93:22:@24087.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_143 ( // @[package.scala 93:22:@24095.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_144 ( // @[package.scala 93:22:@24151.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_145 ( // @[package.scala 93:22:@24159.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_146 ( // @[package.scala 93:22:@24167.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_147 ( // @[package.scala 93:22:@24175.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_148 ( // @[package.scala 93:22:@24183.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_149 ( // @[package.scala 93:22:@24191.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_150 ( // @[package.scala 93:22:@24199.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_151 ( // @[package.scala 93:22:@24207.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_152 ( // @[package.scala 93:22:@24215.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_153 ( // @[package.scala 93:22:@24223.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_154 ( // @[package.scala 93:22:@24231.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_155 ( // @[package.scala 93:22:@24239.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_156 ( // @[package.scala 93:22:@24295.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_157 ( // @[package.scala 93:22:@24303.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_158 ( // @[package.scala 93:22:@24311.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_159 ( // @[package.scala 93:22:@24319.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_160 ( // @[package.scala 93:22:@24327.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_161 ( // @[package.scala 93:22:@24335.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_162 ( // @[package.scala 93:22:@24343.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_163 ( // @[package.scala 93:22:@24351.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_164 ( // @[package.scala 93:22:@24359.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_165 ( // @[package.scala 93:22:@24367.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_166 ( // @[package.scala 93:22:@24375.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_167 ( // @[package.scala 93:22:@24383.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_168 ( // @[package.scala 93:22:@24439.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_169 ( // @[package.scala 93:22:@24447.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_170 ( // @[package.scala 93:22:@24455.4]
    .clock(RetimeWrapper_170_clock),
    .reset(RetimeWrapper_170_reset),
    .io_flow(RetimeWrapper_170_io_flow),
    .io_in(RetimeWrapper_170_io_in),
    .io_out(RetimeWrapper_170_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_171 ( // @[package.scala 93:22:@24463.4]
    .clock(RetimeWrapper_171_clock),
    .reset(RetimeWrapper_171_reset),
    .io_flow(RetimeWrapper_171_io_flow),
    .io_in(RetimeWrapper_171_io_in),
    .io_out(RetimeWrapper_171_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_172 ( // @[package.scala 93:22:@24471.4]
    .clock(RetimeWrapper_172_clock),
    .reset(RetimeWrapper_172_reset),
    .io_flow(RetimeWrapper_172_io_flow),
    .io_in(RetimeWrapper_172_io_in),
    .io_out(RetimeWrapper_172_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_173 ( // @[package.scala 93:22:@24479.4]
    .clock(RetimeWrapper_173_clock),
    .reset(RetimeWrapper_173_reset),
    .io_flow(RetimeWrapper_173_io_flow),
    .io_in(RetimeWrapper_173_io_in),
    .io_out(RetimeWrapper_173_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_174 ( // @[package.scala 93:22:@24487.4]
    .clock(RetimeWrapper_174_clock),
    .reset(RetimeWrapper_174_reset),
    .io_flow(RetimeWrapper_174_io_flow),
    .io_in(RetimeWrapper_174_io_in),
    .io_out(RetimeWrapper_174_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_175 ( // @[package.scala 93:22:@24495.4]
    .clock(RetimeWrapper_175_clock),
    .reset(RetimeWrapper_175_reset),
    .io_flow(RetimeWrapper_175_io_flow),
    .io_in(RetimeWrapper_175_io_in),
    .io_out(RetimeWrapper_175_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_176 ( // @[package.scala 93:22:@24503.4]
    .clock(RetimeWrapper_176_clock),
    .reset(RetimeWrapper_176_reset),
    .io_flow(RetimeWrapper_176_io_flow),
    .io_in(RetimeWrapper_176_io_in),
    .io_out(RetimeWrapper_176_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_177 ( // @[package.scala 93:22:@24511.4]
    .clock(RetimeWrapper_177_clock),
    .reset(RetimeWrapper_177_reset),
    .io_flow(RetimeWrapper_177_io_flow),
    .io_in(RetimeWrapper_177_io_in),
    .io_out(RetimeWrapper_177_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_178 ( // @[package.scala 93:22:@24519.4]
    .clock(RetimeWrapper_178_clock),
    .reset(RetimeWrapper_178_reset),
    .io_flow(RetimeWrapper_178_io_flow),
    .io_in(RetimeWrapper_178_io_in),
    .io_out(RetimeWrapper_178_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_179 ( // @[package.scala 93:22:@24527.4]
    .clock(RetimeWrapper_179_clock),
    .reset(RetimeWrapper_179_reset),
    .io_flow(RetimeWrapper_179_io_flow),
    .io_in(RetimeWrapper_179_io_in),
    .io_out(RetimeWrapper_179_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_180 ( // @[package.scala 93:22:@24583.4]
    .clock(RetimeWrapper_180_clock),
    .reset(RetimeWrapper_180_reset),
    .io_flow(RetimeWrapper_180_io_flow),
    .io_in(RetimeWrapper_180_io_in),
    .io_out(RetimeWrapper_180_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_181 ( // @[package.scala 93:22:@24591.4]
    .clock(RetimeWrapper_181_clock),
    .reset(RetimeWrapper_181_reset),
    .io_flow(RetimeWrapper_181_io_flow),
    .io_in(RetimeWrapper_181_io_in),
    .io_out(RetimeWrapper_181_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_182 ( // @[package.scala 93:22:@24599.4]
    .clock(RetimeWrapper_182_clock),
    .reset(RetimeWrapper_182_reset),
    .io_flow(RetimeWrapper_182_io_flow),
    .io_in(RetimeWrapper_182_io_in),
    .io_out(RetimeWrapper_182_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_183 ( // @[package.scala 93:22:@24607.4]
    .clock(RetimeWrapper_183_clock),
    .reset(RetimeWrapper_183_reset),
    .io_flow(RetimeWrapper_183_io_flow),
    .io_in(RetimeWrapper_183_io_in),
    .io_out(RetimeWrapper_183_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_184 ( // @[package.scala 93:22:@24615.4]
    .clock(RetimeWrapper_184_clock),
    .reset(RetimeWrapper_184_reset),
    .io_flow(RetimeWrapper_184_io_flow),
    .io_in(RetimeWrapper_184_io_in),
    .io_out(RetimeWrapper_184_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_185 ( // @[package.scala 93:22:@24623.4]
    .clock(RetimeWrapper_185_clock),
    .reset(RetimeWrapper_185_reset),
    .io_flow(RetimeWrapper_185_io_flow),
    .io_in(RetimeWrapper_185_io_in),
    .io_out(RetimeWrapper_185_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_186 ( // @[package.scala 93:22:@24631.4]
    .clock(RetimeWrapper_186_clock),
    .reset(RetimeWrapper_186_reset),
    .io_flow(RetimeWrapper_186_io_flow),
    .io_in(RetimeWrapper_186_io_in),
    .io_out(RetimeWrapper_186_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_187 ( // @[package.scala 93:22:@24639.4]
    .clock(RetimeWrapper_187_clock),
    .reset(RetimeWrapper_187_reset),
    .io_flow(RetimeWrapper_187_io_flow),
    .io_in(RetimeWrapper_187_io_in),
    .io_out(RetimeWrapper_187_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_188 ( // @[package.scala 93:22:@24647.4]
    .clock(RetimeWrapper_188_clock),
    .reset(RetimeWrapper_188_reset),
    .io_flow(RetimeWrapper_188_io_flow),
    .io_in(RetimeWrapper_188_io_in),
    .io_out(RetimeWrapper_188_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_189 ( // @[package.scala 93:22:@24655.4]
    .clock(RetimeWrapper_189_clock),
    .reset(RetimeWrapper_189_reset),
    .io_flow(RetimeWrapper_189_io_flow),
    .io_in(RetimeWrapper_189_io_in),
    .io_out(RetimeWrapper_189_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_190 ( // @[package.scala 93:22:@24663.4]
    .clock(RetimeWrapper_190_clock),
    .reset(RetimeWrapper_190_reset),
    .io_flow(RetimeWrapper_190_io_flow),
    .io_in(RetimeWrapper_190_io_in),
    .io_out(RetimeWrapper_190_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_191 ( // @[package.scala 93:22:@24671.4]
    .clock(RetimeWrapper_191_clock),
    .reset(RetimeWrapper_191_reset),
    .io_flow(RetimeWrapper_191_io_flow),
    .io_in(RetimeWrapper_191_io_in),
    .io_out(RetimeWrapper_191_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_192 ( // @[package.scala 93:22:@24727.4]
    .clock(RetimeWrapper_192_clock),
    .reset(RetimeWrapper_192_reset),
    .io_flow(RetimeWrapper_192_io_flow),
    .io_in(RetimeWrapper_192_io_in),
    .io_out(RetimeWrapper_192_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_193 ( // @[package.scala 93:22:@24735.4]
    .clock(RetimeWrapper_193_clock),
    .reset(RetimeWrapper_193_reset),
    .io_flow(RetimeWrapper_193_io_flow),
    .io_in(RetimeWrapper_193_io_in),
    .io_out(RetimeWrapper_193_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_194 ( // @[package.scala 93:22:@24743.4]
    .clock(RetimeWrapper_194_clock),
    .reset(RetimeWrapper_194_reset),
    .io_flow(RetimeWrapper_194_io_flow),
    .io_in(RetimeWrapper_194_io_in),
    .io_out(RetimeWrapper_194_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_195 ( // @[package.scala 93:22:@24751.4]
    .clock(RetimeWrapper_195_clock),
    .reset(RetimeWrapper_195_reset),
    .io_flow(RetimeWrapper_195_io_flow),
    .io_in(RetimeWrapper_195_io_in),
    .io_out(RetimeWrapper_195_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_196 ( // @[package.scala 93:22:@24759.4]
    .clock(RetimeWrapper_196_clock),
    .reset(RetimeWrapper_196_reset),
    .io_flow(RetimeWrapper_196_io_flow),
    .io_in(RetimeWrapper_196_io_in),
    .io_out(RetimeWrapper_196_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_197 ( // @[package.scala 93:22:@24767.4]
    .clock(RetimeWrapper_197_clock),
    .reset(RetimeWrapper_197_reset),
    .io_flow(RetimeWrapper_197_io_flow),
    .io_in(RetimeWrapper_197_io_in),
    .io_out(RetimeWrapper_197_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_198 ( // @[package.scala 93:22:@24775.4]
    .clock(RetimeWrapper_198_clock),
    .reset(RetimeWrapper_198_reset),
    .io_flow(RetimeWrapper_198_io_flow),
    .io_in(RetimeWrapper_198_io_in),
    .io_out(RetimeWrapper_198_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_199 ( // @[package.scala 93:22:@24783.4]
    .clock(RetimeWrapper_199_clock),
    .reset(RetimeWrapper_199_reset),
    .io_flow(RetimeWrapper_199_io_flow),
    .io_in(RetimeWrapper_199_io_in),
    .io_out(RetimeWrapper_199_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_200 ( // @[package.scala 93:22:@24791.4]
    .clock(RetimeWrapper_200_clock),
    .reset(RetimeWrapper_200_reset),
    .io_flow(RetimeWrapper_200_io_flow),
    .io_in(RetimeWrapper_200_io_in),
    .io_out(RetimeWrapper_200_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_201 ( // @[package.scala 93:22:@24799.4]
    .clock(RetimeWrapper_201_clock),
    .reset(RetimeWrapper_201_reset),
    .io_flow(RetimeWrapper_201_io_flow),
    .io_in(RetimeWrapper_201_io_in),
    .io_out(RetimeWrapper_201_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_202 ( // @[package.scala 93:22:@24807.4]
    .clock(RetimeWrapper_202_clock),
    .reset(RetimeWrapper_202_reset),
    .io_flow(RetimeWrapper_202_io_flow),
    .io_in(RetimeWrapper_202_io_in),
    .io_out(RetimeWrapper_202_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_203 ( // @[package.scala 93:22:@24815.4]
    .clock(RetimeWrapper_203_clock),
    .reset(RetimeWrapper_203_reset),
    .io_flow(RetimeWrapper_203_io_flow),
    .io_in(RetimeWrapper_203_io_in),
    .io_out(RetimeWrapper_203_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_204 ( // @[package.scala 93:22:@24871.4]
    .clock(RetimeWrapper_204_clock),
    .reset(RetimeWrapper_204_reset),
    .io_flow(RetimeWrapper_204_io_flow),
    .io_in(RetimeWrapper_204_io_in),
    .io_out(RetimeWrapper_204_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_205 ( // @[package.scala 93:22:@24879.4]
    .clock(RetimeWrapper_205_clock),
    .reset(RetimeWrapper_205_reset),
    .io_flow(RetimeWrapper_205_io_flow),
    .io_in(RetimeWrapper_205_io_in),
    .io_out(RetimeWrapper_205_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_206 ( // @[package.scala 93:22:@24887.4]
    .clock(RetimeWrapper_206_clock),
    .reset(RetimeWrapper_206_reset),
    .io_flow(RetimeWrapper_206_io_flow),
    .io_in(RetimeWrapper_206_io_in),
    .io_out(RetimeWrapper_206_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_207 ( // @[package.scala 93:22:@24895.4]
    .clock(RetimeWrapper_207_clock),
    .reset(RetimeWrapper_207_reset),
    .io_flow(RetimeWrapper_207_io_flow),
    .io_in(RetimeWrapper_207_io_in),
    .io_out(RetimeWrapper_207_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_208 ( // @[package.scala 93:22:@24903.4]
    .clock(RetimeWrapper_208_clock),
    .reset(RetimeWrapper_208_reset),
    .io_flow(RetimeWrapper_208_io_flow),
    .io_in(RetimeWrapper_208_io_in),
    .io_out(RetimeWrapper_208_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_209 ( // @[package.scala 93:22:@24911.4]
    .clock(RetimeWrapper_209_clock),
    .reset(RetimeWrapper_209_reset),
    .io_flow(RetimeWrapper_209_io_flow),
    .io_in(RetimeWrapper_209_io_in),
    .io_out(RetimeWrapper_209_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_210 ( // @[package.scala 93:22:@24919.4]
    .clock(RetimeWrapper_210_clock),
    .reset(RetimeWrapper_210_reset),
    .io_flow(RetimeWrapper_210_io_flow),
    .io_in(RetimeWrapper_210_io_in),
    .io_out(RetimeWrapper_210_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_211 ( // @[package.scala 93:22:@24927.4]
    .clock(RetimeWrapper_211_clock),
    .reset(RetimeWrapper_211_reset),
    .io_flow(RetimeWrapper_211_io_flow),
    .io_in(RetimeWrapper_211_io_in),
    .io_out(RetimeWrapper_211_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_212 ( // @[package.scala 93:22:@24935.4]
    .clock(RetimeWrapper_212_clock),
    .reset(RetimeWrapper_212_reset),
    .io_flow(RetimeWrapper_212_io_flow),
    .io_in(RetimeWrapper_212_io_in),
    .io_out(RetimeWrapper_212_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_213 ( // @[package.scala 93:22:@24943.4]
    .clock(RetimeWrapper_213_clock),
    .reset(RetimeWrapper_213_reset),
    .io_flow(RetimeWrapper_213_io_flow),
    .io_in(RetimeWrapper_213_io_in),
    .io_out(RetimeWrapper_213_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_214 ( // @[package.scala 93:22:@24951.4]
    .clock(RetimeWrapper_214_clock),
    .reset(RetimeWrapper_214_reset),
    .io_flow(RetimeWrapper_214_io_flow),
    .io_in(RetimeWrapper_214_io_in),
    .io_out(RetimeWrapper_214_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_215 ( // @[package.scala 93:22:@24959.4]
    .clock(RetimeWrapper_215_clock),
    .reset(RetimeWrapper_215_reset),
    .io_flow(RetimeWrapper_215_io_flow),
    .io_in(RetimeWrapper_215_io_in),
    .io_out(RetimeWrapper_215_io_out)
  );
  assign _T_700 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@19794.4]
  assign _T_702 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@19795.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 82:228:@19796.4]
  assign _T_704 = io_wPort_0_en_0 & _T_703; // @[MemPrimitives.scala 83:102:@19797.4]
  assign _T_706 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@19798.4]
  assign _T_708 = io_wPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@19799.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 82:228:@19800.4]
  assign _T_710 = io_wPort_2_en_0 & _T_709; // @[MemPrimitives.scala 83:102:@19801.4]
  assign _T_712 = {_T_704,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19803.4]
  assign _T_714 = {_T_710,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@19805.4]
  assign _T_715 = _T_704 ? _T_712 : _T_714; // @[Mux.scala 31:69:@19806.4]
  assign _T_720 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@19813.4]
  assign _T_722 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@19814.4]
  assign _T_723 = _T_720 & _T_722; // @[MemPrimitives.scala 82:228:@19815.4]
  assign _T_724 = io_wPort_1_en_0 & _T_723; // @[MemPrimitives.scala 83:102:@19816.4]
  assign _T_726 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@19817.4]
  assign _T_728 = io_wPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@19818.4]
  assign _T_729 = _T_726 & _T_728; // @[MemPrimitives.scala 82:228:@19819.4]
  assign _T_730 = io_wPort_3_en_0 & _T_729; // @[MemPrimitives.scala 83:102:@19820.4]
  assign _T_732 = {_T_724,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19822.4]
  assign _T_734 = {_T_730,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@19824.4]
  assign _T_735 = _T_724 ? _T_732 : _T_734; // @[Mux.scala 31:69:@19825.4]
  assign _T_742 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@19833.4]
  assign _T_743 = _T_700 & _T_742; // @[MemPrimitives.scala 82:228:@19834.4]
  assign _T_744 = io_wPort_0_en_0 & _T_743; // @[MemPrimitives.scala 83:102:@19835.4]
  assign _T_748 = io_wPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@19837.4]
  assign _T_749 = _T_706 & _T_748; // @[MemPrimitives.scala 82:228:@19838.4]
  assign _T_750 = io_wPort_2_en_0 & _T_749; // @[MemPrimitives.scala 83:102:@19839.4]
  assign _T_752 = {_T_744,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19841.4]
  assign _T_754 = {_T_750,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@19843.4]
  assign _T_755 = _T_744 ? _T_752 : _T_754; // @[Mux.scala 31:69:@19844.4]
  assign _T_762 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@19852.4]
  assign _T_763 = _T_720 & _T_762; // @[MemPrimitives.scala 82:228:@19853.4]
  assign _T_764 = io_wPort_1_en_0 & _T_763; // @[MemPrimitives.scala 83:102:@19854.4]
  assign _T_768 = io_wPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@19856.4]
  assign _T_769 = _T_726 & _T_768; // @[MemPrimitives.scala 82:228:@19857.4]
  assign _T_770 = io_wPort_3_en_0 & _T_769; // @[MemPrimitives.scala 83:102:@19858.4]
  assign _T_772 = {_T_764,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19860.4]
  assign _T_774 = {_T_770,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@19862.4]
  assign _T_775 = _T_764 ? _T_772 : _T_774; // @[Mux.scala 31:69:@19863.4]
  assign _T_782 = io_wPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@19871.4]
  assign _T_783 = _T_700 & _T_782; // @[MemPrimitives.scala 82:228:@19872.4]
  assign _T_784 = io_wPort_0_en_0 & _T_783; // @[MemPrimitives.scala 83:102:@19873.4]
  assign _T_788 = io_wPort_2_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@19875.4]
  assign _T_789 = _T_706 & _T_788; // @[MemPrimitives.scala 82:228:@19876.4]
  assign _T_790 = io_wPort_2_en_0 & _T_789; // @[MemPrimitives.scala 83:102:@19877.4]
  assign _T_792 = {_T_784,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19879.4]
  assign _T_794 = {_T_790,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@19881.4]
  assign _T_795 = _T_784 ? _T_792 : _T_794; // @[Mux.scala 31:69:@19882.4]
  assign _T_802 = io_wPort_1_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@19890.4]
  assign _T_803 = _T_720 & _T_802; // @[MemPrimitives.scala 82:228:@19891.4]
  assign _T_804 = io_wPort_1_en_0 & _T_803; // @[MemPrimitives.scala 83:102:@19892.4]
  assign _T_808 = io_wPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@19894.4]
  assign _T_809 = _T_726 & _T_808; // @[MemPrimitives.scala 82:228:@19895.4]
  assign _T_810 = io_wPort_3_en_0 & _T_809; // @[MemPrimitives.scala 83:102:@19896.4]
  assign _T_812 = {_T_804,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19898.4]
  assign _T_814 = {_T_810,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@19900.4]
  assign _T_815 = _T_804 ? _T_812 : _T_814; // @[Mux.scala 31:69:@19901.4]
  assign _T_820 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@19908.4]
  assign _T_823 = _T_820 & _T_702; // @[MemPrimitives.scala 82:228:@19910.4]
  assign _T_824 = io_wPort_0_en_0 & _T_823; // @[MemPrimitives.scala 83:102:@19911.4]
  assign _T_826 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@19912.4]
  assign _T_829 = _T_826 & _T_708; // @[MemPrimitives.scala 82:228:@19914.4]
  assign _T_830 = io_wPort_2_en_0 & _T_829; // @[MemPrimitives.scala 83:102:@19915.4]
  assign _T_832 = {_T_824,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19917.4]
  assign _T_834 = {_T_830,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@19919.4]
  assign _T_835 = _T_824 ? _T_832 : _T_834; // @[Mux.scala 31:69:@19920.4]
  assign _T_840 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@19927.4]
  assign _T_843 = _T_840 & _T_722; // @[MemPrimitives.scala 82:228:@19929.4]
  assign _T_844 = io_wPort_1_en_0 & _T_843; // @[MemPrimitives.scala 83:102:@19930.4]
  assign _T_846 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@19931.4]
  assign _T_849 = _T_846 & _T_728; // @[MemPrimitives.scala 82:228:@19933.4]
  assign _T_850 = io_wPort_3_en_0 & _T_849; // @[MemPrimitives.scala 83:102:@19934.4]
  assign _T_852 = {_T_844,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19936.4]
  assign _T_854 = {_T_850,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@19938.4]
  assign _T_855 = _T_844 ? _T_852 : _T_854; // @[Mux.scala 31:69:@19939.4]
  assign _T_863 = _T_820 & _T_742; // @[MemPrimitives.scala 82:228:@19948.4]
  assign _T_864 = io_wPort_0_en_0 & _T_863; // @[MemPrimitives.scala 83:102:@19949.4]
  assign _T_869 = _T_826 & _T_748; // @[MemPrimitives.scala 82:228:@19952.4]
  assign _T_870 = io_wPort_2_en_0 & _T_869; // @[MemPrimitives.scala 83:102:@19953.4]
  assign _T_872 = {_T_864,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19955.4]
  assign _T_874 = {_T_870,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@19957.4]
  assign _T_875 = _T_864 ? _T_872 : _T_874; // @[Mux.scala 31:69:@19958.4]
  assign _T_883 = _T_840 & _T_762; // @[MemPrimitives.scala 82:228:@19967.4]
  assign _T_884 = io_wPort_1_en_0 & _T_883; // @[MemPrimitives.scala 83:102:@19968.4]
  assign _T_889 = _T_846 & _T_768; // @[MemPrimitives.scala 82:228:@19971.4]
  assign _T_890 = io_wPort_3_en_0 & _T_889; // @[MemPrimitives.scala 83:102:@19972.4]
  assign _T_892 = {_T_884,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@19974.4]
  assign _T_894 = {_T_890,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@19976.4]
  assign _T_895 = _T_884 ? _T_892 : _T_894; // @[Mux.scala 31:69:@19977.4]
  assign _T_903 = _T_820 & _T_782; // @[MemPrimitives.scala 82:228:@19986.4]
  assign _T_904 = io_wPort_0_en_0 & _T_903; // @[MemPrimitives.scala 83:102:@19987.4]
  assign _T_909 = _T_826 & _T_788; // @[MemPrimitives.scala 82:228:@19990.4]
  assign _T_910 = io_wPort_2_en_0 & _T_909; // @[MemPrimitives.scala 83:102:@19991.4]
  assign _T_912 = {_T_904,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@19993.4]
  assign _T_914 = {_T_910,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@19995.4]
  assign _T_915 = _T_904 ? _T_912 : _T_914; // @[Mux.scala 31:69:@19996.4]
  assign _T_923 = _T_840 & _T_802; // @[MemPrimitives.scala 82:228:@20005.4]
  assign _T_924 = io_wPort_1_en_0 & _T_923; // @[MemPrimitives.scala 83:102:@20006.4]
  assign _T_929 = _T_846 & _T_808; // @[MemPrimitives.scala 82:228:@20009.4]
  assign _T_930 = io_wPort_3_en_0 & _T_929; // @[MemPrimitives.scala 83:102:@20010.4]
  assign _T_932 = {_T_924,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20012.4]
  assign _T_934 = {_T_930,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20014.4]
  assign _T_935 = _T_924 ? _T_932 : _T_934; // @[Mux.scala 31:69:@20015.4]
  assign _T_940 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20022.4]
  assign _T_943 = _T_940 & _T_702; // @[MemPrimitives.scala 82:228:@20024.4]
  assign _T_944 = io_wPort_0_en_0 & _T_943; // @[MemPrimitives.scala 83:102:@20025.4]
  assign _T_946 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20026.4]
  assign _T_949 = _T_946 & _T_708; // @[MemPrimitives.scala 82:228:@20028.4]
  assign _T_950 = io_wPort_2_en_0 & _T_949; // @[MemPrimitives.scala 83:102:@20029.4]
  assign _T_952 = {_T_944,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20031.4]
  assign _T_954 = {_T_950,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20033.4]
  assign _T_955 = _T_944 ? _T_952 : _T_954; // @[Mux.scala 31:69:@20034.4]
  assign _T_960 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20041.4]
  assign _T_963 = _T_960 & _T_722; // @[MemPrimitives.scala 82:228:@20043.4]
  assign _T_964 = io_wPort_1_en_0 & _T_963; // @[MemPrimitives.scala 83:102:@20044.4]
  assign _T_966 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@20045.4]
  assign _T_969 = _T_966 & _T_728; // @[MemPrimitives.scala 82:228:@20047.4]
  assign _T_970 = io_wPort_3_en_0 & _T_969; // @[MemPrimitives.scala 83:102:@20048.4]
  assign _T_972 = {_T_964,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20050.4]
  assign _T_974 = {_T_970,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20052.4]
  assign _T_975 = _T_964 ? _T_972 : _T_974; // @[Mux.scala 31:69:@20053.4]
  assign _T_983 = _T_940 & _T_742; // @[MemPrimitives.scala 82:228:@20062.4]
  assign _T_984 = io_wPort_0_en_0 & _T_983; // @[MemPrimitives.scala 83:102:@20063.4]
  assign _T_989 = _T_946 & _T_748; // @[MemPrimitives.scala 82:228:@20066.4]
  assign _T_990 = io_wPort_2_en_0 & _T_989; // @[MemPrimitives.scala 83:102:@20067.4]
  assign _T_992 = {_T_984,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20069.4]
  assign _T_994 = {_T_990,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20071.4]
  assign _T_995 = _T_984 ? _T_992 : _T_994; // @[Mux.scala 31:69:@20072.4]
  assign _T_1003 = _T_960 & _T_762; // @[MemPrimitives.scala 82:228:@20081.4]
  assign _T_1004 = io_wPort_1_en_0 & _T_1003; // @[MemPrimitives.scala 83:102:@20082.4]
  assign _T_1009 = _T_966 & _T_768; // @[MemPrimitives.scala 82:228:@20085.4]
  assign _T_1010 = io_wPort_3_en_0 & _T_1009; // @[MemPrimitives.scala 83:102:@20086.4]
  assign _T_1012 = {_T_1004,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20088.4]
  assign _T_1014 = {_T_1010,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20090.4]
  assign _T_1015 = _T_1004 ? _T_1012 : _T_1014; // @[Mux.scala 31:69:@20091.4]
  assign _T_1023 = _T_940 & _T_782; // @[MemPrimitives.scala 82:228:@20100.4]
  assign _T_1024 = io_wPort_0_en_0 & _T_1023; // @[MemPrimitives.scala 83:102:@20101.4]
  assign _T_1029 = _T_946 & _T_788; // @[MemPrimitives.scala 82:228:@20104.4]
  assign _T_1030 = io_wPort_2_en_0 & _T_1029; // @[MemPrimitives.scala 83:102:@20105.4]
  assign _T_1032 = {_T_1024,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20107.4]
  assign _T_1034 = {_T_1030,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20109.4]
  assign _T_1035 = _T_1024 ? _T_1032 : _T_1034; // @[Mux.scala 31:69:@20110.4]
  assign _T_1043 = _T_960 & _T_802; // @[MemPrimitives.scala 82:228:@20119.4]
  assign _T_1044 = io_wPort_1_en_0 & _T_1043; // @[MemPrimitives.scala 83:102:@20120.4]
  assign _T_1049 = _T_966 & _T_808; // @[MemPrimitives.scala 82:228:@20123.4]
  assign _T_1050 = io_wPort_3_en_0 & _T_1049; // @[MemPrimitives.scala 83:102:@20124.4]
  assign _T_1052 = {_T_1044,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20126.4]
  assign _T_1054 = {_T_1050,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20128.4]
  assign _T_1055 = _T_1044 ? _T_1052 : _T_1054; // @[Mux.scala 31:69:@20129.4]
  assign _T_1060 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20136.4]
  assign _T_1063 = _T_1060 & _T_702; // @[MemPrimitives.scala 82:228:@20138.4]
  assign _T_1064 = io_wPort_0_en_0 & _T_1063; // @[MemPrimitives.scala 83:102:@20139.4]
  assign _T_1066 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20140.4]
  assign _T_1069 = _T_1066 & _T_708; // @[MemPrimitives.scala 82:228:@20142.4]
  assign _T_1070 = io_wPort_2_en_0 & _T_1069; // @[MemPrimitives.scala 83:102:@20143.4]
  assign _T_1072 = {_T_1064,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20145.4]
  assign _T_1074 = {_T_1070,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20147.4]
  assign _T_1075 = _T_1064 ? _T_1072 : _T_1074; // @[Mux.scala 31:69:@20148.4]
  assign _T_1080 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20155.4]
  assign _T_1083 = _T_1080 & _T_722; // @[MemPrimitives.scala 82:228:@20157.4]
  assign _T_1084 = io_wPort_1_en_0 & _T_1083; // @[MemPrimitives.scala 83:102:@20158.4]
  assign _T_1086 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@20159.4]
  assign _T_1089 = _T_1086 & _T_728; // @[MemPrimitives.scala 82:228:@20161.4]
  assign _T_1090 = io_wPort_3_en_0 & _T_1089; // @[MemPrimitives.scala 83:102:@20162.4]
  assign _T_1092 = {_T_1084,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20164.4]
  assign _T_1094 = {_T_1090,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20166.4]
  assign _T_1095 = _T_1084 ? _T_1092 : _T_1094; // @[Mux.scala 31:69:@20167.4]
  assign _T_1103 = _T_1060 & _T_742; // @[MemPrimitives.scala 82:228:@20176.4]
  assign _T_1104 = io_wPort_0_en_0 & _T_1103; // @[MemPrimitives.scala 83:102:@20177.4]
  assign _T_1109 = _T_1066 & _T_748; // @[MemPrimitives.scala 82:228:@20180.4]
  assign _T_1110 = io_wPort_2_en_0 & _T_1109; // @[MemPrimitives.scala 83:102:@20181.4]
  assign _T_1112 = {_T_1104,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20183.4]
  assign _T_1114 = {_T_1110,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20185.4]
  assign _T_1115 = _T_1104 ? _T_1112 : _T_1114; // @[Mux.scala 31:69:@20186.4]
  assign _T_1123 = _T_1080 & _T_762; // @[MemPrimitives.scala 82:228:@20195.4]
  assign _T_1124 = io_wPort_1_en_0 & _T_1123; // @[MemPrimitives.scala 83:102:@20196.4]
  assign _T_1129 = _T_1086 & _T_768; // @[MemPrimitives.scala 82:228:@20199.4]
  assign _T_1130 = io_wPort_3_en_0 & _T_1129; // @[MemPrimitives.scala 83:102:@20200.4]
  assign _T_1132 = {_T_1124,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20202.4]
  assign _T_1134 = {_T_1130,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20204.4]
  assign _T_1135 = _T_1124 ? _T_1132 : _T_1134; // @[Mux.scala 31:69:@20205.4]
  assign _T_1143 = _T_1060 & _T_782; // @[MemPrimitives.scala 82:228:@20214.4]
  assign _T_1144 = io_wPort_0_en_0 & _T_1143; // @[MemPrimitives.scala 83:102:@20215.4]
  assign _T_1149 = _T_1066 & _T_788; // @[MemPrimitives.scala 82:228:@20218.4]
  assign _T_1150 = io_wPort_2_en_0 & _T_1149; // @[MemPrimitives.scala 83:102:@20219.4]
  assign _T_1152 = {_T_1144,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@20221.4]
  assign _T_1154 = {_T_1150,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@20223.4]
  assign _T_1155 = _T_1144 ? _T_1152 : _T_1154; // @[Mux.scala 31:69:@20224.4]
  assign _T_1163 = _T_1080 & _T_802; // @[MemPrimitives.scala 82:228:@20233.4]
  assign _T_1164 = io_wPort_1_en_0 & _T_1163; // @[MemPrimitives.scala 83:102:@20234.4]
  assign _T_1169 = _T_1086 & _T_808; // @[MemPrimitives.scala 82:228:@20237.4]
  assign _T_1170 = io_wPort_3_en_0 & _T_1169; // @[MemPrimitives.scala 83:102:@20238.4]
  assign _T_1172 = {_T_1164,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@20240.4]
  assign _T_1174 = {_T_1170,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@20242.4]
  assign _T_1175 = _T_1164 ? _T_1172 : _T_1174; // @[Mux.scala 31:69:@20243.4]
  assign _T_1180 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20250.4]
  assign _T_1182 = io_rPort_1_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20251.4]
  assign _T_1183 = _T_1180 & _T_1182; // @[MemPrimitives.scala 110:228:@20252.4]
  assign _T_1186 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20254.4]
  assign _T_1188 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20255.4]
  assign _T_1189 = _T_1186 & _T_1188; // @[MemPrimitives.scala 110:228:@20256.4]
  assign _T_1192 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20258.4]
  assign _T_1194 = io_rPort_5_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20259.4]
  assign _T_1195 = _T_1192 & _T_1194; // @[MemPrimitives.scala 110:228:@20260.4]
  assign _T_1198 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20262.4]
  assign _T_1200 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20263.4]
  assign _T_1201 = _T_1198 & _T_1200; // @[MemPrimitives.scala 110:228:@20264.4]
  assign _T_1204 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20266.4]
  assign _T_1206 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20267.4]
  assign _T_1207 = _T_1204 & _T_1206; // @[MemPrimitives.scala 110:228:@20268.4]
  assign _T_1210 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20270.4]
  assign _T_1212 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20271.4]
  assign _T_1213 = _T_1210 & _T_1212; // @[MemPrimitives.scala 110:228:@20272.4]
  assign _T_1216 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20274.4]
  assign _T_1218 = io_rPort_11_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20275.4]
  assign _T_1219 = _T_1216 & _T_1218; // @[MemPrimitives.scala 110:228:@20276.4]
  assign _T_1222 = io_rPort_13_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20278.4]
  assign _T_1224 = io_rPort_13_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20279.4]
  assign _T_1225 = _T_1222 & _T_1224; // @[MemPrimitives.scala 110:228:@20280.4]
  assign _T_1228 = io_rPort_16_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20282.4]
  assign _T_1230 = io_rPort_16_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@20283.4]
  assign _T_1231 = _T_1228 & _T_1230; // @[MemPrimitives.scala 110:228:@20284.4]
  assign _T_1233 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@20298.4]
  assign _T_1234 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@20299.4]
  assign _T_1235 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@20300.4]
  assign _T_1236 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@20301.4]
  assign _T_1237 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@20302.4]
  assign _T_1238 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@20303.4]
  assign _T_1239 = StickySelects_io_outs_6; // @[MemPrimitives.scala 126:35:@20304.4]
  assign _T_1240 = StickySelects_io_outs_7; // @[MemPrimitives.scala 126:35:@20305.4]
  assign _T_1241 = StickySelects_io_outs_8; // @[MemPrimitives.scala 126:35:@20306.4]
  assign _T_1243 = {_T_1233,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@20308.4]
  assign _T_1245 = {_T_1234,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@20310.4]
  assign _T_1247 = {_T_1235,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@20312.4]
  assign _T_1249 = {_T_1236,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@20314.4]
  assign _T_1251 = {_T_1237,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@20316.4]
  assign _T_1253 = {_T_1238,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@20318.4]
  assign _T_1255 = {_T_1239,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@20320.4]
  assign _T_1257 = {_T_1240,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@20322.4]
  assign _T_1259 = {_T_1241,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@20324.4]
  assign _T_1260 = _T_1240 ? _T_1257 : _T_1259; // @[Mux.scala 31:69:@20325.4]
  assign _T_1261 = _T_1239 ? _T_1255 : _T_1260; // @[Mux.scala 31:69:@20326.4]
  assign _T_1262 = _T_1238 ? _T_1253 : _T_1261; // @[Mux.scala 31:69:@20327.4]
  assign _T_1263 = _T_1237 ? _T_1251 : _T_1262; // @[Mux.scala 31:69:@20328.4]
  assign _T_1264 = _T_1236 ? _T_1249 : _T_1263; // @[Mux.scala 31:69:@20329.4]
  assign _T_1265 = _T_1235 ? _T_1247 : _T_1264; // @[Mux.scala 31:69:@20330.4]
  assign _T_1266 = _T_1234 ? _T_1245 : _T_1265; // @[Mux.scala 31:69:@20331.4]
  assign _T_1267 = _T_1233 ? _T_1243 : _T_1266; // @[Mux.scala 31:69:@20332.4]
  assign _T_1272 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20339.4]
  assign _T_1274 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20340.4]
  assign _T_1275 = _T_1272 & _T_1274; // @[MemPrimitives.scala 110:228:@20341.4]
  assign _T_1278 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20343.4]
  assign _T_1280 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20344.4]
  assign _T_1281 = _T_1278 & _T_1280; // @[MemPrimitives.scala 110:228:@20345.4]
  assign _T_1284 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20347.4]
  assign _T_1286 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20348.4]
  assign _T_1287 = _T_1284 & _T_1286; // @[MemPrimitives.scala 110:228:@20349.4]
  assign _T_1290 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20351.4]
  assign _T_1292 = io_rPort_6_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20352.4]
  assign _T_1293 = _T_1290 & _T_1292; // @[MemPrimitives.scala 110:228:@20353.4]
  assign _T_1296 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20355.4]
  assign _T_1298 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20356.4]
  assign _T_1299 = _T_1296 & _T_1298; // @[MemPrimitives.scala 110:228:@20357.4]
  assign _T_1302 = io_rPort_12_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20359.4]
  assign _T_1304 = io_rPort_12_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20360.4]
  assign _T_1305 = _T_1302 & _T_1304; // @[MemPrimitives.scala 110:228:@20361.4]
  assign _T_1308 = io_rPort_14_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20363.4]
  assign _T_1310 = io_rPort_14_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20364.4]
  assign _T_1311 = _T_1308 & _T_1310; // @[MemPrimitives.scala 110:228:@20365.4]
  assign _T_1314 = io_rPort_15_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20367.4]
  assign _T_1316 = io_rPort_15_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20368.4]
  assign _T_1317 = _T_1314 & _T_1316; // @[MemPrimitives.scala 110:228:@20369.4]
  assign _T_1320 = io_rPort_17_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@20371.4]
  assign _T_1322 = io_rPort_17_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@20372.4]
  assign _T_1323 = _T_1320 & _T_1322; // @[MemPrimitives.scala 110:228:@20373.4]
  assign _T_1325 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@20387.4]
  assign _T_1326 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@20388.4]
  assign _T_1327 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@20389.4]
  assign _T_1328 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@20390.4]
  assign _T_1329 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@20391.4]
  assign _T_1330 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@20392.4]
  assign _T_1331 = StickySelects_1_io_outs_6; // @[MemPrimitives.scala 126:35:@20393.4]
  assign _T_1332 = StickySelects_1_io_outs_7; // @[MemPrimitives.scala 126:35:@20394.4]
  assign _T_1333 = StickySelects_1_io_outs_8; // @[MemPrimitives.scala 126:35:@20395.4]
  assign _T_1335 = {_T_1325,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@20397.4]
  assign _T_1337 = {_T_1326,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@20399.4]
  assign _T_1339 = {_T_1327,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@20401.4]
  assign _T_1341 = {_T_1328,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@20403.4]
  assign _T_1343 = {_T_1329,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@20405.4]
  assign _T_1345 = {_T_1330,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@20407.4]
  assign _T_1347 = {_T_1331,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@20409.4]
  assign _T_1349 = {_T_1332,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@20411.4]
  assign _T_1351 = {_T_1333,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@20413.4]
  assign _T_1352 = _T_1332 ? _T_1349 : _T_1351; // @[Mux.scala 31:69:@20414.4]
  assign _T_1353 = _T_1331 ? _T_1347 : _T_1352; // @[Mux.scala 31:69:@20415.4]
  assign _T_1354 = _T_1330 ? _T_1345 : _T_1353; // @[Mux.scala 31:69:@20416.4]
  assign _T_1355 = _T_1329 ? _T_1343 : _T_1354; // @[Mux.scala 31:69:@20417.4]
  assign _T_1356 = _T_1328 ? _T_1341 : _T_1355; // @[Mux.scala 31:69:@20418.4]
  assign _T_1357 = _T_1327 ? _T_1339 : _T_1356; // @[Mux.scala 31:69:@20419.4]
  assign _T_1358 = _T_1326 ? _T_1337 : _T_1357; // @[Mux.scala 31:69:@20420.4]
  assign _T_1359 = _T_1325 ? _T_1335 : _T_1358; // @[Mux.scala 31:69:@20421.4]
  assign _T_1366 = io_rPort_1_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20429.4]
  assign _T_1367 = _T_1180 & _T_1366; // @[MemPrimitives.scala 110:228:@20430.4]
  assign _T_1372 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20433.4]
  assign _T_1373 = _T_1186 & _T_1372; // @[MemPrimitives.scala 110:228:@20434.4]
  assign _T_1378 = io_rPort_5_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20437.4]
  assign _T_1379 = _T_1192 & _T_1378; // @[MemPrimitives.scala 110:228:@20438.4]
  assign _T_1384 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20441.4]
  assign _T_1385 = _T_1198 & _T_1384; // @[MemPrimitives.scala 110:228:@20442.4]
  assign _T_1390 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20445.4]
  assign _T_1391 = _T_1204 & _T_1390; // @[MemPrimitives.scala 110:228:@20446.4]
  assign _T_1396 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20449.4]
  assign _T_1397 = _T_1210 & _T_1396; // @[MemPrimitives.scala 110:228:@20450.4]
  assign _T_1402 = io_rPort_11_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20453.4]
  assign _T_1403 = _T_1216 & _T_1402; // @[MemPrimitives.scala 110:228:@20454.4]
  assign _T_1408 = io_rPort_13_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20457.4]
  assign _T_1409 = _T_1222 & _T_1408; // @[MemPrimitives.scala 110:228:@20458.4]
  assign _T_1414 = io_rPort_16_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@20461.4]
  assign _T_1415 = _T_1228 & _T_1414; // @[MemPrimitives.scala 110:228:@20462.4]
  assign _T_1417 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@20476.4]
  assign _T_1418 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@20477.4]
  assign _T_1419 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@20478.4]
  assign _T_1420 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@20479.4]
  assign _T_1421 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@20480.4]
  assign _T_1422 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@20481.4]
  assign _T_1423 = StickySelects_2_io_outs_6; // @[MemPrimitives.scala 126:35:@20482.4]
  assign _T_1424 = StickySelects_2_io_outs_7; // @[MemPrimitives.scala 126:35:@20483.4]
  assign _T_1425 = StickySelects_2_io_outs_8; // @[MemPrimitives.scala 126:35:@20484.4]
  assign _T_1427 = {_T_1417,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@20486.4]
  assign _T_1429 = {_T_1418,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@20488.4]
  assign _T_1431 = {_T_1419,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@20490.4]
  assign _T_1433 = {_T_1420,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@20492.4]
  assign _T_1435 = {_T_1421,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@20494.4]
  assign _T_1437 = {_T_1422,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@20496.4]
  assign _T_1439 = {_T_1423,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@20498.4]
  assign _T_1441 = {_T_1424,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@20500.4]
  assign _T_1443 = {_T_1425,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@20502.4]
  assign _T_1444 = _T_1424 ? _T_1441 : _T_1443; // @[Mux.scala 31:69:@20503.4]
  assign _T_1445 = _T_1423 ? _T_1439 : _T_1444; // @[Mux.scala 31:69:@20504.4]
  assign _T_1446 = _T_1422 ? _T_1437 : _T_1445; // @[Mux.scala 31:69:@20505.4]
  assign _T_1447 = _T_1421 ? _T_1435 : _T_1446; // @[Mux.scala 31:69:@20506.4]
  assign _T_1448 = _T_1420 ? _T_1433 : _T_1447; // @[Mux.scala 31:69:@20507.4]
  assign _T_1449 = _T_1419 ? _T_1431 : _T_1448; // @[Mux.scala 31:69:@20508.4]
  assign _T_1450 = _T_1418 ? _T_1429 : _T_1449; // @[Mux.scala 31:69:@20509.4]
  assign _T_1451 = _T_1417 ? _T_1427 : _T_1450; // @[Mux.scala 31:69:@20510.4]
  assign _T_1458 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20518.4]
  assign _T_1459 = _T_1272 & _T_1458; // @[MemPrimitives.scala 110:228:@20519.4]
  assign _T_1464 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20522.4]
  assign _T_1465 = _T_1278 & _T_1464; // @[MemPrimitives.scala 110:228:@20523.4]
  assign _T_1470 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20526.4]
  assign _T_1471 = _T_1284 & _T_1470; // @[MemPrimitives.scala 110:228:@20527.4]
  assign _T_1476 = io_rPort_6_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20530.4]
  assign _T_1477 = _T_1290 & _T_1476; // @[MemPrimitives.scala 110:228:@20531.4]
  assign _T_1482 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20534.4]
  assign _T_1483 = _T_1296 & _T_1482; // @[MemPrimitives.scala 110:228:@20535.4]
  assign _T_1488 = io_rPort_12_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20538.4]
  assign _T_1489 = _T_1302 & _T_1488; // @[MemPrimitives.scala 110:228:@20539.4]
  assign _T_1494 = io_rPort_14_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20542.4]
  assign _T_1495 = _T_1308 & _T_1494; // @[MemPrimitives.scala 110:228:@20543.4]
  assign _T_1500 = io_rPort_15_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20546.4]
  assign _T_1501 = _T_1314 & _T_1500; // @[MemPrimitives.scala 110:228:@20547.4]
  assign _T_1506 = io_rPort_17_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@20550.4]
  assign _T_1507 = _T_1320 & _T_1506; // @[MemPrimitives.scala 110:228:@20551.4]
  assign _T_1509 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@20565.4]
  assign _T_1510 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@20566.4]
  assign _T_1511 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@20567.4]
  assign _T_1512 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@20568.4]
  assign _T_1513 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@20569.4]
  assign _T_1514 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@20570.4]
  assign _T_1515 = StickySelects_3_io_outs_6; // @[MemPrimitives.scala 126:35:@20571.4]
  assign _T_1516 = StickySelects_3_io_outs_7; // @[MemPrimitives.scala 126:35:@20572.4]
  assign _T_1517 = StickySelects_3_io_outs_8; // @[MemPrimitives.scala 126:35:@20573.4]
  assign _T_1519 = {_T_1509,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@20575.4]
  assign _T_1521 = {_T_1510,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@20577.4]
  assign _T_1523 = {_T_1511,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@20579.4]
  assign _T_1525 = {_T_1512,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@20581.4]
  assign _T_1527 = {_T_1513,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@20583.4]
  assign _T_1529 = {_T_1514,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@20585.4]
  assign _T_1531 = {_T_1515,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@20587.4]
  assign _T_1533 = {_T_1516,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@20589.4]
  assign _T_1535 = {_T_1517,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@20591.4]
  assign _T_1536 = _T_1516 ? _T_1533 : _T_1535; // @[Mux.scala 31:69:@20592.4]
  assign _T_1537 = _T_1515 ? _T_1531 : _T_1536; // @[Mux.scala 31:69:@20593.4]
  assign _T_1538 = _T_1514 ? _T_1529 : _T_1537; // @[Mux.scala 31:69:@20594.4]
  assign _T_1539 = _T_1513 ? _T_1527 : _T_1538; // @[Mux.scala 31:69:@20595.4]
  assign _T_1540 = _T_1512 ? _T_1525 : _T_1539; // @[Mux.scala 31:69:@20596.4]
  assign _T_1541 = _T_1511 ? _T_1523 : _T_1540; // @[Mux.scala 31:69:@20597.4]
  assign _T_1542 = _T_1510 ? _T_1521 : _T_1541; // @[Mux.scala 31:69:@20598.4]
  assign _T_1543 = _T_1509 ? _T_1519 : _T_1542; // @[Mux.scala 31:69:@20599.4]
  assign _T_1550 = io_rPort_1_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20607.4]
  assign _T_1551 = _T_1180 & _T_1550; // @[MemPrimitives.scala 110:228:@20608.4]
  assign _T_1556 = io_rPort_4_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20611.4]
  assign _T_1557 = _T_1186 & _T_1556; // @[MemPrimitives.scala 110:228:@20612.4]
  assign _T_1562 = io_rPort_5_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20615.4]
  assign _T_1563 = _T_1192 & _T_1562; // @[MemPrimitives.scala 110:228:@20616.4]
  assign _T_1568 = io_rPort_7_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20619.4]
  assign _T_1569 = _T_1198 & _T_1568; // @[MemPrimitives.scala 110:228:@20620.4]
  assign _T_1574 = io_rPort_8_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20623.4]
  assign _T_1575 = _T_1204 & _T_1574; // @[MemPrimitives.scala 110:228:@20624.4]
  assign _T_1580 = io_rPort_10_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20627.4]
  assign _T_1581 = _T_1210 & _T_1580; // @[MemPrimitives.scala 110:228:@20628.4]
  assign _T_1586 = io_rPort_11_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20631.4]
  assign _T_1587 = _T_1216 & _T_1586; // @[MemPrimitives.scala 110:228:@20632.4]
  assign _T_1592 = io_rPort_13_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20635.4]
  assign _T_1593 = _T_1222 & _T_1592; // @[MemPrimitives.scala 110:228:@20636.4]
  assign _T_1598 = io_rPort_16_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@20639.4]
  assign _T_1599 = _T_1228 & _T_1598; // @[MemPrimitives.scala 110:228:@20640.4]
  assign _T_1601 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@20654.4]
  assign _T_1602 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@20655.4]
  assign _T_1603 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@20656.4]
  assign _T_1604 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@20657.4]
  assign _T_1605 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@20658.4]
  assign _T_1606 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@20659.4]
  assign _T_1607 = StickySelects_4_io_outs_6; // @[MemPrimitives.scala 126:35:@20660.4]
  assign _T_1608 = StickySelects_4_io_outs_7; // @[MemPrimitives.scala 126:35:@20661.4]
  assign _T_1609 = StickySelects_4_io_outs_8; // @[MemPrimitives.scala 126:35:@20662.4]
  assign _T_1611 = {_T_1601,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@20664.4]
  assign _T_1613 = {_T_1602,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@20666.4]
  assign _T_1615 = {_T_1603,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@20668.4]
  assign _T_1617 = {_T_1604,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@20670.4]
  assign _T_1619 = {_T_1605,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@20672.4]
  assign _T_1621 = {_T_1606,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@20674.4]
  assign _T_1623 = {_T_1607,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@20676.4]
  assign _T_1625 = {_T_1608,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@20678.4]
  assign _T_1627 = {_T_1609,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@20680.4]
  assign _T_1628 = _T_1608 ? _T_1625 : _T_1627; // @[Mux.scala 31:69:@20681.4]
  assign _T_1629 = _T_1607 ? _T_1623 : _T_1628; // @[Mux.scala 31:69:@20682.4]
  assign _T_1630 = _T_1606 ? _T_1621 : _T_1629; // @[Mux.scala 31:69:@20683.4]
  assign _T_1631 = _T_1605 ? _T_1619 : _T_1630; // @[Mux.scala 31:69:@20684.4]
  assign _T_1632 = _T_1604 ? _T_1617 : _T_1631; // @[Mux.scala 31:69:@20685.4]
  assign _T_1633 = _T_1603 ? _T_1615 : _T_1632; // @[Mux.scala 31:69:@20686.4]
  assign _T_1634 = _T_1602 ? _T_1613 : _T_1633; // @[Mux.scala 31:69:@20687.4]
  assign _T_1635 = _T_1601 ? _T_1611 : _T_1634; // @[Mux.scala 31:69:@20688.4]
  assign _T_1642 = io_rPort_0_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20696.4]
  assign _T_1643 = _T_1272 & _T_1642; // @[MemPrimitives.scala 110:228:@20697.4]
  assign _T_1648 = io_rPort_2_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20700.4]
  assign _T_1649 = _T_1278 & _T_1648; // @[MemPrimitives.scala 110:228:@20701.4]
  assign _T_1654 = io_rPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20704.4]
  assign _T_1655 = _T_1284 & _T_1654; // @[MemPrimitives.scala 110:228:@20705.4]
  assign _T_1660 = io_rPort_6_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20708.4]
  assign _T_1661 = _T_1290 & _T_1660; // @[MemPrimitives.scala 110:228:@20709.4]
  assign _T_1666 = io_rPort_9_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20712.4]
  assign _T_1667 = _T_1296 & _T_1666; // @[MemPrimitives.scala 110:228:@20713.4]
  assign _T_1672 = io_rPort_12_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20716.4]
  assign _T_1673 = _T_1302 & _T_1672; // @[MemPrimitives.scala 110:228:@20717.4]
  assign _T_1678 = io_rPort_14_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20720.4]
  assign _T_1679 = _T_1308 & _T_1678; // @[MemPrimitives.scala 110:228:@20721.4]
  assign _T_1684 = io_rPort_15_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20724.4]
  assign _T_1685 = _T_1314 & _T_1684; // @[MemPrimitives.scala 110:228:@20725.4]
  assign _T_1690 = io_rPort_17_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@20728.4]
  assign _T_1691 = _T_1320 & _T_1690; // @[MemPrimitives.scala 110:228:@20729.4]
  assign _T_1693 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@20743.4]
  assign _T_1694 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@20744.4]
  assign _T_1695 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@20745.4]
  assign _T_1696 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@20746.4]
  assign _T_1697 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@20747.4]
  assign _T_1698 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@20748.4]
  assign _T_1699 = StickySelects_5_io_outs_6; // @[MemPrimitives.scala 126:35:@20749.4]
  assign _T_1700 = StickySelects_5_io_outs_7; // @[MemPrimitives.scala 126:35:@20750.4]
  assign _T_1701 = StickySelects_5_io_outs_8; // @[MemPrimitives.scala 126:35:@20751.4]
  assign _T_1703 = {_T_1693,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@20753.4]
  assign _T_1705 = {_T_1694,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@20755.4]
  assign _T_1707 = {_T_1695,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@20757.4]
  assign _T_1709 = {_T_1696,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@20759.4]
  assign _T_1711 = {_T_1697,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@20761.4]
  assign _T_1713 = {_T_1698,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@20763.4]
  assign _T_1715 = {_T_1699,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@20765.4]
  assign _T_1717 = {_T_1700,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@20767.4]
  assign _T_1719 = {_T_1701,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@20769.4]
  assign _T_1720 = _T_1700 ? _T_1717 : _T_1719; // @[Mux.scala 31:69:@20770.4]
  assign _T_1721 = _T_1699 ? _T_1715 : _T_1720; // @[Mux.scala 31:69:@20771.4]
  assign _T_1722 = _T_1698 ? _T_1713 : _T_1721; // @[Mux.scala 31:69:@20772.4]
  assign _T_1723 = _T_1697 ? _T_1711 : _T_1722; // @[Mux.scala 31:69:@20773.4]
  assign _T_1724 = _T_1696 ? _T_1709 : _T_1723; // @[Mux.scala 31:69:@20774.4]
  assign _T_1725 = _T_1695 ? _T_1707 : _T_1724; // @[Mux.scala 31:69:@20775.4]
  assign _T_1726 = _T_1694 ? _T_1705 : _T_1725; // @[Mux.scala 31:69:@20776.4]
  assign _T_1727 = _T_1693 ? _T_1703 : _T_1726; // @[Mux.scala 31:69:@20777.4]
  assign _T_1732 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20784.4]
  assign _T_1735 = _T_1732 & _T_1182; // @[MemPrimitives.scala 110:228:@20786.4]
  assign _T_1738 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20788.4]
  assign _T_1741 = _T_1738 & _T_1188; // @[MemPrimitives.scala 110:228:@20790.4]
  assign _T_1744 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20792.4]
  assign _T_1747 = _T_1744 & _T_1194; // @[MemPrimitives.scala 110:228:@20794.4]
  assign _T_1750 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20796.4]
  assign _T_1753 = _T_1750 & _T_1200; // @[MemPrimitives.scala 110:228:@20798.4]
  assign _T_1756 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20800.4]
  assign _T_1759 = _T_1756 & _T_1206; // @[MemPrimitives.scala 110:228:@20802.4]
  assign _T_1762 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20804.4]
  assign _T_1765 = _T_1762 & _T_1212; // @[MemPrimitives.scala 110:228:@20806.4]
  assign _T_1768 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20808.4]
  assign _T_1771 = _T_1768 & _T_1218; // @[MemPrimitives.scala 110:228:@20810.4]
  assign _T_1774 = io_rPort_13_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20812.4]
  assign _T_1777 = _T_1774 & _T_1224; // @[MemPrimitives.scala 110:228:@20814.4]
  assign _T_1780 = io_rPort_16_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20816.4]
  assign _T_1783 = _T_1780 & _T_1230; // @[MemPrimitives.scala 110:228:@20818.4]
  assign _T_1785 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@20832.4]
  assign _T_1786 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@20833.4]
  assign _T_1787 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@20834.4]
  assign _T_1788 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@20835.4]
  assign _T_1789 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@20836.4]
  assign _T_1790 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@20837.4]
  assign _T_1791 = StickySelects_6_io_outs_6; // @[MemPrimitives.scala 126:35:@20838.4]
  assign _T_1792 = StickySelects_6_io_outs_7; // @[MemPrimitives.scala 126:35:@20839.4]
  assign _T_1793 = StickySelects_6_io_outs_8; // @[MemPrimitives.scala 126:35:@20840.4]
  assign _T_1795 = {_T_1785,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@20842.4]
  assign _T_1797 = {_T_1786,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@20844.4]
  assign _T_1799 = {_T_1787,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@20846.4]
  assign _T_1801 = {_T_1788,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@20848.4]
  assign _T_1803 = {_T_1789,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@20850.4]
  assign _T_1805 = {_T_1790,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@20852.4]
  assign _T_1807 = {_T_1791,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@20854.4]
  assign _T_1809 = {_T_1792,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@20856.4]
  assign _T_1811 = {_T_1793,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@20858.4]
  assign _T_1812 = _T_1792 ? _T_1809 : _T_1811; // @[Mux.scala 31:69:@20859.4]
  assign _T_1813 = _T_1791 ? _T_1807 : _T_1812; // @[Mux.scala 31:69:@20860.4]
  assign _T_1814 = _T_1790 ? _T_1805 : _T_1813; // @[Mux.scala 31:69:@20861.4]
  assign _T_1815 = _T_1789 ? _T_1803 : _T_1814; // @[Mux.scala 31:69:@20862.4]
  assign _T_1816 = _T_1788 ? _T_1801 : _T_1815; // @[Mux.scala 31:69:@20863.4]
  assign _T_1817 = _T_1787 ? _T_1799 : _T_1816; // @[Mux.scala 31:69:@20864.4]
  assign _T_1818 = _T_1786 ? _T_1797 : _T_1817; // @[Mux.scala 31:69:@20865.4]
  assign _T_1819 = _T_1785 ? _T_1795 : _T_1818; // @[Mux.scala 31:69:@20866.4]
  assign _T_1824 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20873.4]
  assign _T_1827 = _T_1824 & _T_1274; // @[MemPrimitives.scala 110:228:@20875.4]
  assign _T_1830 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20877.4]
  assign _T_1833 = _T_1830 & _T_1280; // @[MemPrimitives.scala 110:228:@20879.4]
  assign _T_1836 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20881.4]
  assign _T_1839 = _T_1836 & _T_1286; // @[MemPrimitives.scala 110:228:@20883.4]
  assign _T_1842 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20885.4]
  assign _T_1845 = _T_1842 & _T_1292; // @[MemPrimitives.scala 110:228:@20887.4]
  assign _T_1848 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20889.4]
  assign _T_1851 = _T_1848 & _T_1298; // @[MemPrimitives.scala 110:228:@20891.4]
  assign _T_1854 = io_rPort_12_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20893.4]
  assign _T_1857 = _T_1854 & _T_1304; // @[MemPrimitives.scala 110:228:@20895.4]
  assign _T_1860 = io_rPort_14_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20897.4]
  assign _T_1863 = _T_1860 & _T_1310; // @[MemPrimitives.scala 110:228:@20899.4]
  assign _T_1866 = io_rPort_15_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20901.4]
  assign _T_1869 = _T_1866 & _T_1316; // @[MemPrimitives.scala 110:228:@20903.4]
  assign _T_1872 = io_rPort_17_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@20905.4]
  assign _T_1875 = _T_1872 & _T_1322; // @[MemPrimitives.scala 110:228:@20907.4]
  assign _T_1877 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@20921.4]
  assign _T_1878 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@20922.4]
  assign _T_1879 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@20923.4]
  assign _T_1880 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@20924.4]
  assign _T_1881 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@20925.4]
  assign _T_1882 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@20926.4]
  assign _T_1883 = StickySelects_7_io_outs_6; // @[MemPrimitives.scala 126:35:@20927.4]
  assign _T_1884 = StickySelects_7_io_outs_7; // @[MemPrimitives.scala 126:35:@20928.4]
  assign _T_1885 = StickySelects_7_io_outs_8; // @[MemPrimitives.scala 126:35:@20929.4]
  assign _T_1887 = {_T_1877,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@20931.4]
  assign _T_1889 = {_T_1878,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@20933.4]
  assign _T_1891 = {_T_1879,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@20935.4]
  assign _T_1893 = {_T_1880,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@20937.4]
  assign _T_1895 = {_T_1881,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@20939.4]
  assign _T_1897 = {_T_1882,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@20941.4]
  assign _T_1899 = {_T_1883,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@20943.4]
  assign _T_1901 = {_T_1884,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@20945.4]
  assign _T_1903 = {_T_1885,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@20947.4]
  assign _T_1904 = _T_1884 ? _T_1901 : _T_1903; // @[Mux.scala 31:69:@20948.4]
  assign _T_1905 = _T_1883 ? _T_1899 : _T_1904; // @[Mux.scala 31:69:@20949.4]
  assign _T_1906 = _T_1882 ? _T_1897 : _T_1905; // @[Mux.scala 31:69:@20950.4]
  assign _T_1907 = _T_1881 ? _T_1895 : _T_1906; // @[Mux.scala 31:69:@20951.4]
  assign _T_1908 = _T_1880 ? _T_1893 : _T_1907; // @[Mux.scala 31:69:@20952.4]
  assign _T_1909 = _T_1879 ? _T_1891 : _T_1908; // @[Mux.scala 31:69:@20953.4]
  assign _T_1910 = _T_1878 ? _T_1889 : _T_1909; // @[Mux.scala 31:69:@20954.4]
  assign _T_1911 = _T_1877 ? _T_1887 : _T_1910; // @[Mux.scala 31:69:@20955.4]
  assign _T_1919 = _T_1732 & _T_1366; // @[MemPrimitives.scala 110:228:@20964.4]
  assign _T_1925 = _T_1738 & _T_1372; // @[MemPrimitives.scala 110:228:@20968.4]
  assign _T_1931 = _T_1744 & _T_1378; // @[MemPrimitives.scala 110:228:@20972.4]
  assign _T_1937 = _T_1750 & _T_1384; // @[MemPrimitives.scala 110:228:@20976.4]
  assign _T_1943 = _T_1756 & _T_1390; // @[MemPrimitives.scala 110:228:@20980.4]
  assign _T_1949 = _T_1762 & _T_1396; // @[MemPrimitives.scala 110:228:@20984.4]
  assign _T_1955 = _T_1768 & _T_1402; // @[MemPrimitives.scala 110:228:@20988.4]
  assign _T_1961 = _T_1774 & _T_1408; // @[MemPrimitives.scala 110:228:@20992.4]
  assign _T_1967 = _T_1780 & _T_1414; // @[MemPrimitives.scala 110:228:@20996.4]
  assign _T_1969 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@21010.4]
  assign _T_1970 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@21011.4]
  assign _T_1971 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@21012.4]
  assign _T_1972 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@21013.4]
  assign _T_1973 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@21014.4]
  assign _T_1974 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@21015.4]
  assign _T_1975 = StickySelects_8_io_outs_6; // @[MemPrimitives.scala 126:35:@21016.4]
  assign _T_1976 = StickySelects_8_io_outs_7; // @[MemPrimitives.scala 126:35:@21017.4]
  assign _T_1977 = StickySelects_8_io_outs_8; // @[MemPrimitives.scala 126:35:@21018.4]
  assign _T_1979 = {_T_1969,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21020.4]
  assign _T_1981 = {_T_1970,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21022.4]
  assign _T_1983 = {_T_1971,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21024.4]
  assign _T_1985 = {_T_1972,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21026.4]
  assign _T_1987 = {_T_1973,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21028.4]
  assign _T_1989 = {_T_1974,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21030.4]
  assign _T_1991 = {_T_1975,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21032.4]
  assign _T_1993 = {_T_1976,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21034.4]
  assign _T_1995 = {_T_1977,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21036.4]
  assign _T_1996 = _T_1976 ? _T_1993 : _T_1995; // @[Mux.scala 31:69:@21037.4]
  assign _T_1997 = _T_1975 ? _T_1991 : _T_1996; // @[Mux.scala 31:69:@21038.4]
  assign _T_1998 = _T_1974 ? _T_1989 : _T_1997; // @[Mux.scala 31:69:@21039.4]
  assign _T_1999 = _T_1973 ? _T_1987 : _T_1998; // @[Mux.scala 31:69:@21040.4]
  assign _T_2000 = _T_1972 ? _T_1985 : _T_1999; // @[Mux.scala 31:69:@21041.4]
  assign _T_2001 = _T_1971 ? _T_1983 : _T_2000; // @[Mux.scala 31:69:@21042.4]
  assign _T_2002 = _T_1970 ? _T_1981 : _T_2001; // @[Mux.scala 31:69:@21043.4]
  assign _T_2003 = _T_1969 ? _T_1979 : _T_2002; // @[Mux.scala 31:69:@21044.4]
  assign _T_2011 = _T_1824 & _T_1458; // @[MemPrimitives.scala 110:228:@21053.4]
  assign _T_2017 = _T_1830 & _T_1464; // @[MemPrimitives.scala 110:228:@21057.4]
  assign _T_2023 = _T_1836 & _T_1470; // @[MemPrimitives.scala 110:228:@21061.4]
  assign _T_2029 = _T_1842 & _T_1476; // @[MemPrimitives.scala 110:228:@21065.4]
  assign _T_2035 = _T_1848 & _T_1482; // @[MemPrimitives.scala 110:228:@21069.4]
  assign _T_2041 = _T_1854 & _T_1488; // @[MemPrimitives.scala 110:228:@21073.4]
  assign _T_2047 = _T_1860 & _T_1494; // @[MemPrimitives.scala 110:228:@21077.4]
  assign _T_2053 = _T_1866 & _T_1500; // @[MemPrimitives.scala 110:228:@21081.4]
  assign _T_2059 = _T_1872 & _T_1506; // @[MemPrimitives.scala 110:228:@21085.4]
  assign _T_2061 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@21099.4]
  assign _T_2062 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@21100.4]
  assign _T_2063 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@21101.4]
  assign _T_2064 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@21102.4]
  assign _T_2065 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@21103.4]
  assign _T_2066 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@21104.4]
  assign _T_2067 = StickySelects_9_io_outs_6; // @[MemPrimitives.scala 126:35:@21105.4]
  assign _T_2068 = StickySelects_9_io_outs_7; // @[MemPrimitives.scala 126:35:@21106.4]
  assign _T_2069 = StickySelects_9_io_outs_8; // @[MemPrimitives.scala 126:35:@21107.4]
  assign _T_2071 = {_T_2061,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21109.4]
  assign _T_2073 = {_T_2062,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21111.4]
  assign _T_2075 = {_T_2063,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21113.4]
  assign _T_2077 = {_T_2064,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21115.4]
  assign _T_2079 = {_T_2065,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21117.4]
  assign _T_2081 = {_T_2066,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21119.4]
  assign _T_2083 = {_T_2067,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21121.4]
  assign _T_2085 = {_T_2068,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21123.4]
  assign _T_2087 = {_T_2069,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21125.4]
  assign _T_2088 = _T_2068 ? _T_2085 : _T_2087; // @[Mux.scala 31:69:@21126.4]
  assign _T_2089 = _T_2067 ? _T_2083 : _T_2088; // @[Mux.scala 31:69:@21127.4]
  assign _T_2090 = _T_2066 ? _T_2081 : _T_2089; // @[Mux.scala 31:69:@21128.4]
  assign _T_2091 = _T_2065 ? _T_2079 : _T_2090; // @[Mux.scala 31:69:@21129.4]
  assign _T_2092 = _T_2064 ? _T_2077 : _T_2091; // @[Mux.scala 31:69:@21130.4]
  assign _T_2093 = _T_2063 ? _T_2075 : _T_2092; // @[Mux.scala 31:69:@21131.4]
  assign _T_2094 = _T_2062 ? _T_2073 : _T_2093; // @[Mux.scala 31:69:@21132.4]
  assign _T_2095 = _T_2061 ? _T_2071 : _T_2094; // @[Mux.scala 31:69:@21133.4]
  assign _T_2103 = _T_1732 & _T_1550; // @[MemPrimitives.scala 110:228:@21142.4]
  assign _T_2109 = _T_1738 & _T_1556; // @[MemPrimitives.scala 110:228:@21146.4]
  assign _T_2115 = _T_1744 & _T_1562; // @[MemPrimitives.scala 110:228:@21150.4]
  assign _T_2121 = _T_1750 & _T_1568; // @[MemPrimitives.scala 110:228:@21154.4]
  assign _T_2127 = _T_1756 & _T_1574; // @[MemPrimitives.scala 110:228:@21158.4]
  assign _T_2133 = _T_1762 & _T_1580; // @[MemPrimitives.scala 110:228:@21162.4]
  assign _T_2139 = _T_1768 & _T_1586; // @[MemPrimitives.scala 110:228:@21166.4]
  assign _T_2145 = _T_1774 & _T_1592; // @[MemPrimitives.scala 110:228:@21170.4]
  assign _T_2151 = _T_1780 & _T_1598; // @[MemPrimitives.scala 110:228:@21174.4]
  assign _T_2153 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@21188.4]
  assign _T_2154 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@21189.4]
  assign _T_2155 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@21190.4]
  assign _T_2156 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@21191.4]
  assign _T_2157 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@21192.4]
  assign _T_2158 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@21193.4]
  assign _T_2159 = StickySelects_10_io_outs_6; // @[MemPrimitives.scala 126:35:@21194.4]
  assign _T_2160 = StickySelects_10_io_outs_7; // @[MemPrimitives.scala 126:35:@21195.4]
  assign _T_2161 = StickySelects_10_io_outs_8; // @[MemPrimitives.scala 126:35:@21196.4]
  assign _T_2163 = {_T_2153,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21198.4]
  assign _T_2165 = {_T_2154,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21200.4]
  assign _T_2167 = {_T_2155,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21202.4]
  assign _T_2169 = {_T_2156,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21204.4]
  assign _T_2171 = {_T_2157,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21206.4]
  assign _T_2173 = {_T_2158,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21208.4]
  assign _T_2175 = {_T_2159,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21210.4]
  assign _T_2177 = {_T_2160,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21212.4]
  assign _T_2179 = {_T_2161,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21214.4]
  assign _T_2180 = _T_2160 ? _T_2177 : _T_2179; // @[Mux.scala 31:69:@21215.4]
  assign _T_2181 = _T_2159 ? _T_2175 : _T_2180; // @[Mux.scala 31:69:@21216.4]
  assign _T_2182 = _T_2158 ? _T_2173 : _T_2181; // @[Mux.scala 31:69:@21217.4]
  assign _T_2183 = _T_2157 ? _T_2171 : _T_2182; // @[Mux.scala 31:69:@21218.4]
  assign _T_2184 = _T_2156 ? _T_2169 : _T_2183; // @[Mux.scala 31:69:@21219.4]
  assign _T_2185 = _T_2155 ? _T_2167 : _T_2184; // @[Mux.scala 31:69:@21220.4]
  assign _T_2186 = _T_2154 ? _T_2165 : _T_2185; // @[Mux.scala 31:69:@21221.4]
  assign _T_2187 = _T_2153 ? _T_2163 : _T_2186; // @[Mux.scala 31:69:@21222.4]
  assign _T_2195 = _T_1824 & _T_1642; // @[MemPrimitives.scala 110:228:@21231.4]
  assign _T_2201 = _T_1830 & _T_1648; // @[MemPrimitives.scala 110:228:@21235.4]
  assign _T_2207 = _T_1836 & _T_1654; // @[MemPrimitives.scala 110:228:@21239.4]
  assign _T_2213 = _T_1842 & _T_1660; // @[MemPrimitives.scala 110:228:@21243.4]
  assign _T_2219 = _T_1848 & _T_1666; // @[MemPrimitives.scala 110:228:@21247.4]
  assign _T_2225 = _T_1854 & _T_1672; // @[MemPrimitives.scala 110:228:@21251.4]
  assign _T_2231 = _T_1860 & _T_1678; // @[MemPrimitives.scala 110:228:@21255.4]
  assign _T_2237 = _T_1866 & _T_1684; // @[MemPrimitives.scala 110:228:@21259.4]
  assign _T_2243 = _T_1872 & _T_1690; // @[MemPrimitives.scala 110:228:@21263.4]
  assign _T_2245 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@21277.4]
  assign _T_2246 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@21278.4]
  assign _T_2247 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@21279.4]
  assign _T_2248 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@21280.4]
  assign _T_2249 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@21281.4]
  assign _T_2250 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@21282.4]
  assign _T_2251 = StickySelects_11_io_outs_6; // @[MemPrimitives.scala 126:35:@21283.4]
  assign _T_2252 = StickySelects_11_io_outs_7; // @[MemPrimitives.scala 126:35:@21284.4]
  assign _T_2253 = StickySelects_11_io_outs_8; // @[MemPrimitives.scala 126:35:@21285.4]
  assign _T_2255 = {_T_2245,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21287.4]
  assign _T_2257 = {_T_2246,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21289.4]
  assign _T_2259 = {_T_2247,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21291.4]
  assign _T_2261 = {_T_2248,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21293.4]
  assign _T_2263 = {_T_2249,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21295.4]
  assign _T_2265 = {_T_2250,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21297.4]
  assign _T_2267 = {_T_2251,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21299.4]
  assign _T_2269 = {_T_2252,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21301.4]
  assign _T_2271 = {_T_2253,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21303.4]
  assign _T_2272 = _T_2252 ? _T_2269 : _T_2271; // @[Mux.scala 31:69:@21304.4]
  assign _T_2273 = _T_2251 ? _T_2267 : _T_2272; // @[Mux.scala 31:69:@21305.4]
  assign _T_2274 = _T_2250 ? _T_2265 : _T_2273; // @[Mux.scala 31:69:@21306.4]
  assign _T_2275 = _T_2249 ? _T_2263 : _T_2274; // @[Mux.scala 31:69:@21307.4]
  assign _T_2276 = _T_2248 ? _T_2261 : _T_2275; // @[Mux.scala 31:69:@21308.4]
  assign _T_2277 = _T_2247 ? _T_2259 : _T_2276; // @[Mux.scala 31:69:@21309.4]
  assign _T_2278 = _T_2246 ? _T_2257 : _T_2277; // @[Mux.scala 31:69:@21310.4]
  assign _T_2279 = _T_2245 ? _T_2255 : _T_2278; // @[Mux.scala 31:69:@21311.4]
  assign _T_2284 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21318.4]
  assign _T_2287 = _T_2284 & _T_1182; // @[MemPrimitives.scala 110:228:@21320.4]
  assign _T_2290 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21322.4]
  assign _T_2293 = _T_2290 & _T_1188; // @[MemPrimitives.scala 110:228:@21324.4]
  assign _T_2296 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21326.4]
  assign _T_2299 = _T_2296 & _T_1194; // @[MemPrimitives.scala 110:228:@21328.4]
  assign _T_2302 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21330.4]
  assign _T_2305 = _T_2302 & _T_1200; // @[MemPrimitives.scala 110:228:@21332.4]
  assign _T_2308 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21334.4]
  assign _T_2311 = _T_2308 & _T_1206; // @[MemPrimitives.scala 110:228:@21336.4]
  assign _T_2314 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21338.4]
  assign _T_2317 = _T_2314 & _T_1212; // @[MemPrimitives.scala 110:228:@21340.4]
  assign _T_2320 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21342.4]
  assign _T_2323 = _T_2320 & _T_1218; // @[MemPrimitives.scala 110:228:@21344.4]
  assign _T_2326 = io_rPort_13_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21346.4]
  assign _T_2329 = _T_2326 & _T_1224; // @[MemPrimitives.scala 110:228:@21348.4]
  assign _T_2332 = io_rPort_16_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21350.4]
  assign _T_2335 = _T_2332 & _T_1230; // @[MemPrimitives.scala 110:228:@21352.4]
  assign _T_2337 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@21366.4]
  assign _T_2338 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@21367.4]
  assign _T_2339 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@21368.4]
  assign _T_2340 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@21369.4]
  assign _T_2341 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 126:35:@21370.4]
  assign _T_2342 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 126:35:@21371.4]
  assign _T_2343 = StickySelects_12_io_outs_6; // @[MemPrimitives.scala 126:35:@21372.4]
  assign _T_2344 = StickySelects_12_io_outs_7; // @[MemPrimitives.scala 126:35:@21373.4]
  assign _T_2345 = StickySelects_12_io_outs_8; // @[MemPrimitives.scala 126:35:@21374.4]
  assign _T_2347 = {_T_2337,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21376.4]
  assign _T_2349 = {_T_2338,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21378.4]
  assign _T_2351 = {_T_2339,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21380.4]
  assign _T_2353 = {_T_2340,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21382.4]
  assign _T_2355 = {_T_2341,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21384.4]
  assign _T_2357 = {_T_2342,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21386.4]
  assign _T_2359 = {_T_2343,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21388.4]
  assign _T_2361 = {_T_2344,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21390.4]
  assign _T_2363 = {_T_2345,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21392.4]
  assign _T_2364 = _T_2344 ? _T_2361 : _T_2363; // @[Mux.scala 31:69:@21393.4]
  assign _T_2365 = _T_2343 ? _T_2359 : _T_2364; // @[Mux.scala 31:69:@21394.4]
  assign _T_2366 = _T_2342 ? _T_2357 : _T_2365; // @[Mux.scala 31:69:@21395.4]
  assign _T_2367 = _T_2341 ? _T_2355 : _T_2366; // @[Mux.scala 31:69:@21396.4]
  assign _T_2368 = _T_2340 ? _T_2353 : _T_2367; // @[Mux.scala 31:69:@21397.4]
  assign _T_2369 = _T_2339 ? _T_2351 : _T_2368; // @[Mux.scala 31:69:@21398.4]
  assign _T_2370 = _T_2338 ? _T_2349 : _T_2369; // @[Mux.scala 31:69:@21399.4]
  assign _T_2371 = _T_2337 ? _T_2347 : _T_2370; // @[Mux.scala 31:69:@21400.4]
  assign _T_2376 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21407.4]
  assign _T_2379 = _T_2376 & _T_1274; // @[MemPrimitives.scala 110:228:@21409.4]
  assign _T_2382 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21411.4]
  assign _T_2385 = _T_2382 & _T_1280; // @[MemPrimitives.scala 110:228:@21413.4]
  assign _T_2388 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21415.4]
  assign _T_2391 = _T_2388 & _T_1286; // @[MemPrimitives.scala 110:228:@21417.4]
  assign _T_2394 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21419.4]
  assign _T_2397 = _T_2394 & _T_1292; // @[MemPrimitives.scala 110:228:@21421.4]
  assign _T_2400 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21423.4]
  assign _T_2403 = _T_2400 & _T_1298; // @[MemPrimitives.scala 110:228:@21425.4]
  assign _T_2406 = io_rPort_12_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21427.4]
  assign _T_2409 = _T_2406 & _T_1304; // @[MemPrimitives.scala 110:228:@21429.4]
  assign _T_2412 = io_rPort_14_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21431.4]
  assign _T_2415 = _T_2412 & _T_1310; // @[MemPrimitives.scala 110:228:@21433.4]
  assign _T_2418 = io_rPort_15_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21435.4]
  assign _T_2421 = _T_2418 & _T_1316; // @[MemPrimitives.scala 110:228:@21437.4]
  assign _T_2424 = io_rPort_17_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@21439.4]
  assign _T_2427 = _T_2424 & _T_1322; // @[MemPrimitives.scala 110:228:@21441.4]
  assign _T_2429 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@21455.4]
  assign _T_2430 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@21456.4]
  assign _T_2431 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@21457.4]
  assign _T_2432 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@21458.4]
  assign _T_2433 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@21459.4]
  assign _T_2434 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@21460.4]
  assign _T_2435 = StickySelects_13_io_outs_6; // @[MemPrimitives.scala 126:35:@21461.4]
  assign _T_2436 = StickySelects_13_io_outs_7; // @[MemPrimitives.scala 126:35:@21462.4]
  assign _T_2437 = StickySelects_13_io_outs_8; // @[MemPrimitives.scala 126:35:@21463.4]
  assign _T_2439 = {_T_2429,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21465.4]
  assign _T_2441 = {_T_2430,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21467.4]
  assign _T_2443 = {_T_2431,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21469.4]
  assign _T_2445 = {_T_2432,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21471.4]
  assign _T_2447 = {_T_2433,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21473.4]
  assign _T_2449 = {_T_2434,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21475.4]
  assign _T_2451 = {_T_2435,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21477.4]
  assign _T_2453 = {_T_2436,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21479.4]
  assign _T_2455 = {_T_2437,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21481.4]
  assign _T_2456 = _T_2436 ? _T_2453 : _T_2455; // @[Mux.scala 31:69:@21482.4]
  assign _T_2457 = _T_2435 ? _T_2451 : _T_2456; // @[Mux.scala 31:69:@21483.4]
  assign _T_2458 = _T_2434 ? _T_2449 : _T_2457; // @[Mux.scala 31:69:@21484.4]
  assign _T_2459 = _T_2433 ? _T_2447 : _T_2458; // @[Mux.scala 31:69:@21485.4]
  assign _T_2460 = _T_2432 ? _T_2445 : _T_2459; // @[Mux.scala 31:69:@21486.4]
  assign _T_2461 = _T_2431 ? _T_2443 : _T_2460; // @[Mux.scala 31:69:@21487.4]
  assign _T_2462 = _T_2430 ? _T_2441 : _T_2461; // @[Mux.scala 31:69:@21488.4]
  assign _T_2463 = _T_2429 ? _T_2439 : _T_2462; // @[Mux.scala 31:69:@21489.4]
  assign _T_2471 = _T_2284 & _T_1366; // @[MemPrimitives.scala 110:228:@21498.4]
  assign _T_2477 = _T_2290 & _T_1372; // @[MemPrimitives.scala 110:228:@21502.4]
  assign _T_2483 = _T_2296 & _T_1378; // @[MemPrimitives.scala 110:228:@21506.4]
  assign _T_2489 = _T_2302 & _T_1384; // @[MemPrimitives.scala 110:228:@21510.4]
  assign _T_2495 = _T_2308 & _T_1390; // @[MemPrimitives.scala 110:228:@21514.4]
  assign _T_2501 = _T_2314 & _T_1396; // @[MemPrimitives.scala 110:228:@21518.4]
  assign _T_2507 = _T_2320 & _T_1402; // @[MemPrimitives.scala 110:228:@21522.4]
  assign _T_2513 = _T_2326 & _T_1408; // @[MemPrimitives.scala 110:228:@21526.4]
  assign _T_2519 = _T_2332 & _T_1414; // @[MemPrimitives.scala 110:228:@21530.4]
  assign _T_2521 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@21544.4]
  assign _T_2522 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@21545.4]
  assign _T_2523 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@21546.4]
  assign _T_2524 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@21547.4]
  assign _T_2525 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 126:35:@21548.4]
  assign _T_2526 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 126:35:@21549.4]
  assign _T_2527 = StickySelects_14_io_outs_6; // @[MemPrimitives.scala 126:35:@21550.4]
  assign _T_2528 = StickySelects_14_io_outs_7; // @[MemPrimitives.scala 126:35:@21551.4]
  assign _T_2529 = StickySelects_14_io_outs_8; // @[MemPrimitives.scala 126:35:@21552.4]
  assign _T_2531 = {_T_2521,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21554.4]
  assign _T_2533 = {_T_2522,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21556.4]
  assign _T_2535 = {_T_2523,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21558.4]
  assign _T_2537 = {_T_2524,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21560.4]
  assign _T_2539 = {_T_2525,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21562.4]
  assign _T_2541 = {_T_2526,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21564.4]
  assign _T_2543 = {_T_2527,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21566.4]
  assign _T_2545 = {_T_2528,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21568.4]
  assign _T_2547 = {_T_2529,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21570.4]
  assign _T_2548 = _T_2528 ? _T_2545 : _T_2547; // @[Mux.scala 31:69:@21571.4]
  assign _T_2549 = _T_2527 ? _T_2543 : _T_2548; // @[Mux.scala 31:69:@21572.4]
  assign _T_2550 = _T_2526 ? _T_2541 : _T_2549; // @[Mux.scala 31:69:@21573.4]
  assign _T_2551 = _T_2525 ? _T_2539 : _T_2550; // @[Mux.scala 31:69:@21574.4]
  assign _T_2552 = _T_2524 ? _T_2537 : _T_2551; // @[Mux.scala 31:69:@21575.4]
  assign _T_2553 = _T_2523 ? _T_2535 : _T_2552; // @[Mux.scala 31:69:@21576.4]
  assign _T_2554 = _T_2522 ? _T_2533 : _T_2553; // @[Mux.scala 31:69:@21577.4]
  assign _T_2555 = _T_2521 ? _T_2531 : _T_2554; // @[Mux.scala 31:69:@21578.4]
  assign _T_2563 = _T_2376 & _T_1458; // @[MemPrimitives.scala 110:228:@21587.4]
  assign _T_2569 = _T_2382 & _T_1464; // @[MemPrimitives.scala 110:228:@21591.4]
  assign _T_2575 = _T_2388 & _T_1470; // @[MemPrimitives.scala 110:228:@21595.4]
  assign _T_2581 = _T_2394 & _T_1476; // @[MemPrimitives.scala 110:228:@21599.4]
  assign _T_2587 = _T_2400 & _T_1482; // @[MemPrimitives.scala 110:228:@21603.4]
  assign _T_2593 = _T_2406 & _T_1488; // @[MemPrimitives.scala 110:228:@21607.4]
  assign _T_2599 = _T_2412 & _T_1494; // @[MemPrimitives.scala 110:228:@21611.4]
  assign _T_2605 = _T_2418 & _T_1500; // @[MemPrimitives.scala 110:228:@21615.4]
  assign _T_2611 = _T_2424 & _T_1506; // @[MemPrimitives.scala 110:228:@21619.4]
  assign _T_2613 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@21633.4]
  assign _T_2614 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@21634.4]
  assign _T_2615 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@21635.4]
  assign _T_2616 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@21636.4]
  assign _T_2617 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@21637.4]
  assign _T_2618 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@21638.4]
  assign _T_2619 = StickySelects_15_io_outs_6; // @[MemPrimitives.scala 126:35:@21639.4]
  assign _T_2620 = StickySelects_15_io_outs_7; // @[MemPrimitives.scala 126:35:@21640.4]
  assign _T_2621 = StickySelects_15_io_outs_8; // @[MemPrimitives.scala 126:35:@21641.4]
  assign _T_2623 = {_T_2613,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21643.4]
  assign _T_2625 = {_T_2614,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21645.4]
  assign _T_2627 = {_T_2615,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21647.4]
  assign _T_2629 = {_T_2616,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21649.4]
  assign _T_2631 = {_T_2617,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21651.4]
  assign _T_2633 = {_T_2618,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21653.4]
  assign _T_2635 = {_T_2619,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21655.4]
  assign _T_2637 = {_T_2620,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21657.4]
  assign _T_2639 = {_T_2621,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21659.4]
  assign _T_2640 = _T_2620 ? _T_2637 : _T_2639; // @[Mux.scala 31:69:@21660.4]
  assign _T_2641 = _T_2619 ? _T_2635 : _T_2640; // @[Mux.scala 31:69:@21661.4]
  assign _T_2642 = _T_2618 ? _T_2633 : _T_2641; // @[Mux.scala 31:69:@21662.4]
  assign _T_2643 = _T_2617 ? _T_2631 : _T_2642; // @[Mux.scala 31:69:@21663.4]
  assign _T_2644 = _T_2616 ? _T_2629 : _T_2643; // @[Mux.scala 31:69:@21664.4]
  assign _T_2645 = _T_2615 ? _T_2627 : _T_2644; // @[Mux.scala 31:69:@21665.4]
  assign _T_2646 = _T_2614 ? _T_2625 : _T_2645; // @[Mux.scala 31:69:@21666.4]
  assign _T_2647 = _T_2613 ? _T_2623 : _T_2646; // @[Mux.scala 31:69:@21667.4]
  assign _T_2655 = _T_2284 & _T_1550; // @[MemPrimitives.scala 110:228:@21676.4]
  assign _T_2661 = _T_2290 & _T_1556; // @[MemPrimitives.scala 110:228:@21680.4]
  assign _T_2667 = _T_2296 & _T_1562; // @[MemPrimitives.scala 110:228:@21684.4]
  assign _T_2673 = _T_2302 & _T_1568; // @[MemPrimitives.scala 110:228:@21688.4]
  assign _T_2679 = _T_2308 & _T_1574; // @[MemPrimitives.scala 110:228:@21692.4]
  assign _T_2685 = _T_2314 & _T_1580; // @[MemPrimitives.scala 110:228:@21696.4]
  assign _T_2691 = _T_2320 & _T_1586; // @[MemPrimitives.scala 110:228:@21700.4]
  assign _T_2697 = _T_2326 & _T_1592; // @[MemPrimitives.scala 110:228:@21704.4]
  assign _T_2703 = _T_2332 & _T_1598; // @[MemPrimitives.scala 110:228:@21708.4]
  assign _T_2705 = StickySelects_16_io_outs_0; // @[MemPrimitives.scala 126:35:@21722.4]
  assign _T_2706 = StickySelects_16_io_outs_1; // @[MemPrimitives.scala 126:35:@21723.4]
  assign _T_2707 = StickySelects_16_io_outs_2; // @[MemPrimitives.scala 126:35:@21724.4]
  assign _T_2708 = StickySelects_16_io_outs_3; // @[MemPrimitives.scala 126:35:@21725.4]
  assign _T_2709 = StickySelects_16_io_outs_4; // @[MemPrimitives.scala 126:35:@21726.4]
  assign _T_2710 = StickySelects_16_io_outs_5; // @[MemPrimitives.scala 126:35:@21727.4]
  assign _T_2711 = StickySelects_16_io_outs_6; // @[MemPrimitives.scala 126:35:@21728.4]
  assign _T_2712 = StickySelects_16_io_outs_7; // @[MemPrimitives.scala 126:35:@21729.4]
  assign _T_2713 = StickySelects_16_io_outs_8; // @[MemPrimitives.scala 126:35:@21730.4]
  assign _T_2715 = {_T_2705,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21732.4]
  assign _T_2717 = {_T_2706,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21734.4]
  assign _T_2719 = {_T_2707,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21736.4]
  assign _T_2721 = {_T_2708,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21738.4]
  assign _T_2723 = {_T_2709,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21740.4]
  assign _T_2725 = {_T_2710,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21742.4]
  assign _T_2727 = {_T_2711,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21744.4]
  assign _T_2729 = {_T_2712,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21746.4]
  assign _T_2731 = {_T_2713,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21748.4]
  assign _T_2732 = _T_2712 ? _T_2729 : _T_2731; // @[Mux.scala 31:69:@21749.4]
  assign _T_2733 = _T_2711 ? _T_2727 : _T_2732; // @[Mux.scala 31:69:@21750.4]
  assign _T_2734 = _T_2710 ? _T_2725 : _T_2733; // @[Mux.scala 31:69:@21751.4]
  assign _T_2735 = _T_2709 ? _T_2723 : _T_2734; // @[Mux.scala 31:69:@21752.4]
  assign _T_2736 = _T_2708 ? _T_2721 : _T_2735; // @[Mux.scala 31:69:@21753.4]
  assign _T_2737 = _T_2707 ? _T_2719 : _T_2736; // @[Mux.scala 31:69:@21754.4]
  assign _T_2738 = _T_2706 ? _T_2717 : _T_2737; // @[Mux.scala 31:69:@21755.4]
  assign _T_2739 = _T_2705 ? _T_2715 : _T_2738; // @[Mux.scala 31:69:@21756.4]
  assign _T_2747 = _T_2376 & _T_1642; // @[MemPrimitives.scala 110:228:@21765.4]
  assign _T_2753 = _T_2382 & _T_1648; // @[MemPrimitives.scala 110:228:@21769.4]
  assign _T_2759 = _T_2388 & _T_1654; // @[MemPrimitives.scala 110:228:@21773.4]
  assign _T_2765 = _T_2394 & _T_1660; // @[MemPrimitives.scala 110:228:@21777.4]
  assign _T_2771 = _T_2400 & _T_1666; // @[MemPrimitives.scala 110:228:@21781.4]
  assign _T_2777 = _T_2406 & _T_1672; // @[MemPrimitives.scala 110:228:@21785.4]
  assign _T_2783 = _T_2412 & _T_1678; // @[MemPrimitives.scala 110:228:@21789.4]
  assign _T_2789 = _T_2418 & _T_1684; // @[MemPrimitives.scala 110:228:@21793.4]
  assign _T_2795 = _T_2424 & _T_1690; // @[MemPrimitives.scala 110:228:@21797.4]
  assign _T_2797 = StickySelects_17_io_outs_0; // @[MemPrimitives.scala 126:35:@21811.4]
  assign _T_2798 = StickySelects_17_io_outs_1; // @[MemPrimitives.scala 126:35:@21812.4]
  assign _T_2799 = StickySelects_17_io_outs_2; // @[MemPrimitives.scala 126:35:@21813.4]
  assign _T_2800 = StickySelects_17_io_outs_3; // @[MemPrimitives.scala 126:35:@21814.4]
  assign _T_2801 = StickySelects_17_io_outs_4; // @[MemPrimitives.scala 126:35:@21815.4]
  assign _T_2802 = StickySelects_17_io_outs_5; // @[MemPrimitives.scala 126:35:@21816.4]
  assign _T_2803 = StickySelects_17_io_outs_6; // @[MemPrimitives.scala 126:35:@21817.4]
  assign _T_2804 = StickySelects_17_io_outs_7; // @[MemPrimitives.scala 126:35:@21818.4]
  assign _T_2805 = StickySelects_17_io_outs_8; // @[MemPrimitives.scala 126:35:@21819.4]
  assign _T_2807 = {_T_2797,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21821.4]
  assign _T_2809 = {_T_2798,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@21823.4]
  assign _T_2811 = {_T_2799,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@21825.4]
  assign _T_2813 = {_T_2800,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@21827.4]
  assign _T_2815 = {_T_2801,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@21829.4]
  assign _T_2817 = {_T_2802,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@21831.4]
  assign _T_2819 = {_T_2803,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@21833.4]
  assign _T_2821 = {_T_2804,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@21835.4]
  assign _T_2823 = {_T_2805,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@21837.4]
  assign _T_2824 = _T_2804 ? _T_2821 : _T_2823; // @[Mux.scala 31:69:@21838.4]
  assign _T_2825 = _T_2803 ? _T_2819 : _T_2824; // @[Mux.scala 31:69:@21839.4]
  assign _T_2826 = _T_2802 ? _T_2817 : _T_2825; // @[Mux.scala 31:69:@21840.4]
  assign _T_2827 = _T_2801 ? _T_2815 : _T_2826; // @[Mux.scala 31:69:@21841.4]
  assign _T_2828 = _T_2800 ? _T_2813 : _T_2827; // @[Mux.scala 31:69:@21842.4]
  assign _T_2829 = _T_2799 ? _T_2811 : _T_2828; // @[Mux.scala 31:69:@21843.4]
  assign _T_2830 = _T_2798 ? _T_2809 : _T_2829; // @[Mux.scala 31:69:@21844.4]
  assign _T_2831 = _T_2797 ? _T_2807 : _T_2830; // @[Mux.scala 31:69:@21845.4]
  assign _T_2836 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21852.4]
  assign _T_2839 = _T_2836 & _T_1182; // @[MemPrimitives.scala 110:228:@21854.4]
  assign _T_2842 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21856.4]
  assign _T_2845 = _T_2842 & _T_1188; // @[MemPrimitives.scala 110:228:@21858.4]
  assign _T_2848 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21860.4]
  assign _T_2851 = _T_2848 & _T_1194; // @[MemPrimitives.scala 110:228:@21862.4]
  assign _T_2854 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21864.4]
  assign _T_2857 = _T_2854 & _T_1200; // @[MemPrimitives.scala 110:228:@21866.4]
  assign _T_2860 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21868.4]
  assign _T_2863 = _T_2860 & _T_1206; // @[MemPrimitives.scala 110:228:@21870.4]
  assign _T_2866 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21872.4]
  assign _T_2869 = _T_2866 & _T_1212; // @[MemPrimitives.scala 110:228:@21874.4]
  assign _T_2872 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21876.4]
  assign _T_2875 = _T_2872 & _T_1218; // @[MemPrimitives.scala 110:228:@21878.4]
  assign _T_2878 = io_rPort_13_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21880.4]
  assign _T_2881 = _T_2878 & _T_1224; // @[MemPrimitives.scala 110:228:@21882.4]
  assign _T_2884 = io_rPort_16_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21884.4]
  assign _T_2887 = _T_2884 & _T_1230; // @[MemPrimitives.scala 110:228:@21886.4]
  assign _T_2889 = StickySelects_18_io_outs_0; // @[MemPrimitives.scala 126:35:@21900.4]
  assign _T_2890 = StickySelects_18_io_outs_1; // @[MemPrimitives.scala 126:35:@21901.4]
  assign _T_2891 = StickySelects_18_io_outs_2; // @[MemPrimitives.scala 126:35:@21902.4]
  assign _T_2892 = StickySelects_18_io_outs_3; // @[MemPrimitives.scala 126:35:@21903.4]
  assign _T_2893 = StickySelects_18_io_outs_4; // @[MemPrimitives.scala 126:35:@21904.4]
  assign _T_2894 = StickySelects_18_io_outs_5; // @[MemPrimitives.scala 126:35:@21905.4]
  assign _T_2895 = StickySelects_18_io_outs_6; // @[MemPrimitives.scala 126:35:@21906.4]
  assign _T_2896 = StickySelects_18_io_outs_7; // @[MemPrimitives.scala 126:35:@21907.4]
  assign _T_2897 = StickySelects_18_io_outs_8; // @[MemPrimitives.scala 126:35:@21908.4]
  assign _T_2899 = {_T_2889,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@21910.4]
  assign _T_2901 = {_T_2890,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@21912.4]
  assign _T_2903 = {_T_2891,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@21914.4]
  assign _T_2905 = {_T_2892,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@21916.4]
  assign _T_2907 = {_T_2893,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@21918.4]
  assign _T_2909 = {_T_2894,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@21920.4]
  assign _T_2911 = {_T_2895,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@21922.4]
  assign _T_2913 = {_T_2896,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@21924.4]
  assign _T_2915 = {_T_2897,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@21926.4]
  assign _T_2916 = _T_2896 ? _T_2913 : _T_2915; // @[Mux.scala 31:69:@21927.4]
  assign _T_2917 = _T_2895 ? _T_2911 : _T_2916; // @[Mux.scala 31:69:@21928.4]
  assign _T_2918 = _T_2894 ? _T_2909 : _T_2917; // @[Mux.scala 31:69:@21929.4]
  assign _T_2919 = _T_2893 ? _T_2907 : _T_2918; // @[Mux.scala 31:69:@21930.4]
  assign _T_2920 = _T_2892 ? _T_2905 : _T_2919; // @[Mux.scala 31:69:@21931.4]
  assign _T_2921 = _T_2891 ? _T_2903 : _T_2920; // @[Mux.scala 31:69:@21932.4]
  assign _T_2922 = _T_2890 ? _T_2901 : _T_2921; // @[Mux.scala 31:69:@21933.4]
  assign _T_2923 = _T_2889 ? _T_2899 : _T_2922; // @[Mux.scala 31:69:@21934.4]
  assign _T_2928 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21941.4]
  assign _T_2931 = _T_2928 & _T_1274; // @[MemPrimitives.scala 110:228:@21943.4]
  assign _T_2934 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21945.4]
  assign _T_2937 = _T_2934 & _T_1280; // @[MemPrimitives.scala 110:228:@21947.4]
  assign _T_2940 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21949.4]
  assign _T_2943 = _T_2940 & _T_1286; // @[MemPrimitives.scala 110:228:@21951.4]
  assign _T_2946 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21953.4]
  assign _T_2949 = _T_2946 & _T_1292; // @[MemPrimitives.scala 110:228:@21955.4]
  assign _T_2952 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21957.4]
  assign _T_2955 = _T_2952 & _T_1298; // @[MemPrimitives.scala 110:228:@21959.4]
  assign _T_2958 = io_rPort_12_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21961.4]
  assign _T_2961 = _T_2958 & _T_1304; // @[MemPrimitives.scala 110:228:@21963.4]
  assign _T_2964 = io_rPort_14_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21965.4]
  assign _T_2967 = _T_2964 & _T_1310; // @[MemPrimitives.scala 110:228:@21967.4]
  assign _T_2970 = io_rPort_15_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21969.4]
  assign _T_2973 = _T_2970 & _T_1316; // @[MemPrimitives.scala 110:228:@21971.4]
  assign _T_2976 = io_rPort_17_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@21973.4]
  assign _T_2979 = _T_2976 & _T_1322; // @[MemPrimitives.scala 110:228:@21975.4]
  assign _T_2981 = StickySelects_19_io_outs_0; // @[MemPrimitives.scala 126:35:@21989.4]
  assign _T_2982 = StickySelects_19_io_outs_1; // @[MemPrimitives.scala 126:35:@21990.4]
  assign _T_2983 = StickySelects_19_io_outs_2; // @[MemPrimitives.scala 126:35:@21991.4]
  assign _T_2984 = StickySelects_19_io_outs_3; // @[MemPrimitives.scala 126:35:@21992.4]
  assign _T_2985 = StickySelects_19_io_outs_4; // @[MemPrimitives.scala 126:35:@21993.4]
  assign _T_2986 = StickySelects_19_io_outs_5; // @[MemPrimitives.scala 126:35:@21994.4]
  assign _T_2987 = StickySelects_19_io_outs_6; // @[MemPrimitives.scala 126:35:@21995.4]
  assign _T_2988 = StickySelects_19_io_outs_7; // @[MemPrimitives.scala 126:35:@21996.4]
  assign _T_2989 = StickySelects_19_io_outs_8; // @[MemPrimitives.scala 126:35:@21997.4]
  assign _T_2991 = {_T_2981,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@21999.4]
  assign _T_2993 = {_T_2982,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22001.4]
  assign _T_2995 = {_T_2983,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22003.4]
  assign _T_2997 = {_T_2984,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22005.4]
  assign _T_2999 = {_T_2985,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22007.4]
  assign _T_3001 = {_T_2986,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22009.4]
  assign _T_3003 = {_T_2987,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22011.4]
  assign _T_3005 = {_T_2988,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22013.4]
  assign _T_3007 = {_T_2989,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22015.4]
  assign _T_3008 = _T_2988 ? _T_3005 : _T_3007; // @[Mux.scala 31:69:@22016.4]
  assign _T_3009 = _T_2987 ? _T_3003 : _T_3008; // @[Mux.scala 31:69:@22017.4]
  assign _T_3010 = _T_2986 ? _T_3001 : _T_3009; // @[Mux.scala 31:69:@22018.4]
  assign _T_3011 = _T_2985 ? _T_2999 : _T_3010; // @[Mux.scala 31:69:@22019.4]
  assign _T_3012 = _T_2984 ? _T_2997 : _T_3011; // @[Mux.scala 31:69:@22020.4]
  assign _T_3013 = _T_2983 ? _T_2995 : _T_3012; // @[Mux.scala 31:69:@22021.4]
  assign _T_3014 = _T_2982 ? _T_2993 : _T_3013; // @[Mux.scala 31:69:@22022.4]
  assign _T_3015 = _T_2981 ? _T_2991 : _T_3014; // @[Mux.scala 31:69:@22023.4]
  assign _T_3023 = _T_2836 & _T_1366; // @[MemPrimitives.scala 110:228:@22032.4]
  assign _T_3029 = _T_2842 & _T_1372; // @[MemPrimitives.scala 110:228:@22036.4]
  assign _T_3035 = _T_2848 & _T_1378; // @[MemPrimitives.scala 110:228:@22040.4]
  assign _T_3041 = _T_2854 & _T_1384; // @[MemPrimitives.scala 110:228:@22044.4]
  assign _T_3047 = _T_2860 & _T_1390; // @[MemPrimitives.scala 110:228:@22048.4]
  assign _T_3053 = _T_2866 & _T_1396; // @[MemPrimitives.scala 110:228:@22052.4]
  assign _T_3059 = _T_2872 & _T_1402; // @[MemPrimitives.scala 110:228:@22056.4]
  assign _T_3065 = _T_2878 & _T_1408; // @[MemPrimitives.scala 110:228:@22060.4]
  assign _T_3071 = _T_2884 & _T_1414; // @[MemPrimitives.scala 110:228:@22064.4]
  assign _T_3073 = StickySelects_20_io_outs_0; // @[MemPrimitives.scala 126:35:@22078.4]
  assign _T_3074 = StickySelects_20_io_outs_1; // @[MemPrimitives.scala 126:35:@22079.4]
  assign _T_3075 = StickySelects_20_io_outs_2; // @[MemPrimitives.scala 126:35:@22080.4]
  assign _T_3076 = StickySelects_20_io_outs_3; // @[MemPrimitives.scala 126:35:@22081.4]
  assign _T_3077 = StickySelects_20_io_outs_4; // @[MemPrimitives.scala 126:35:@22082.4]
  assign _T_3078 = StickySelects_20_io_outs_5; // @[MemPrimitives.scala 126:35:@22083.4]
  assign _T_3079 = StickySelects_20_io_outs_6; // @[MemPrimitives.scala 126:35:@22084.4]
  assign _T_3080 = StickySelects_20_io_outs_7; // @[MemPrimitives.scala 126:35:@22085.4]
  assign _T_3081 = StickySelects_20_io_outs_8; // @[MemPrimitives.scala 126:35:@22086.4]
  assign _T_3083 = {_T_3073,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22088.4]
  assign _T_3085 = {_T_3074,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22090.4]
  assign _T_3087 = {_T_3075,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22092.4]
  assign _T_3089 = {_T_3076,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22094.4]
  assign _T_3091 = {_T_3077,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22096.4]
  assign _T_3093 = {_T_3078,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22098.4]
  assign _T_3095 = {_T_3079,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22100.4]
  assign _T_3097 = {_T_3080,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22102.4]
  assign _T_3099 = {_T_3081,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22104.4]
  assign _T_3100 = _T_3080 ? _T_3097 : _T_3099; // @[Mux.scala 31:69:@22105.4]
  assign _T_3101 = _T_3079 ? _T_3095 : _T_3100; // @[Mux.scala 31:69:@22106.4]
  assign _T_3102 = _T_3078 ? _T_3093 : _T_3101; // @[Mux.scala 31:69:@22107.4]
  assign _T_3103 = _T_3077 ? _T_3091 : _T_3102; // @[Mux.scala 31:69:@22108.4]
  assign _T_3104 = _T_3076 ? _T_3089 : _T_3103; // @[Mux.scala 31:69:@22109.4]
  assign _T_3105 = _T_3075 ? _T_3087 : _T_3104; // @[Mux.scala 31:69:@22110.4]
  assign _T_3106 = _T_3074 ? _T_3085 : _T_3105; // @[Mux.scala 31:69:@22111.4]
  assign _T_3107 = _T_3073 ? _T_3083 : _T_3106; // @[Mux.scala 31:69:@22112.4]
  assign _T_3115 = _T_2928 & _T_1458; // @[MemPrimitives.scala 110:228:@22121.4]
  assign _T_3121 = _T_2934 & _T_1464; // @[MemPrimitives.scala 110:228:@22125.4]
  assign _T_3127 = _T_2940 & _T_1470; // @[MemPrimitives.scala 110:228:@22129.4]
  assign _T_3133 = _T_2946 & _T_1476; // @[MemPrimitives.scala 110:228:@22133.4]
  assign _T_3139 = _T_2952 & _T_1482; // @[MemPrimitives.scala 110:228:@22137.4]
  assign _T_3145 = _T_2958 & _T_1488; // @[MemPrimitives.scala 110:228:@22141.4]
  assign _T_3151 = _T_2964 & _T_1494; // @[MemPrimitives.scala 110:228:@22145.4]
  assign _T_3157 = _T_2970 & _T_1500; // @[MemPrimitives.scala 110:228:@22149.4]
  assign _T_3163 = _T_2976 & _T_1506; // @[MemPrimitives.scala 110:228:@22153.4]
  assign _T_3165 = StickySelects_21_io_outs_0; // @[MemPrimitives.scala 126:35:@22167.4]
  assign _T_3166 = StickySelects_21_io_outs_1; // @[MemPrimitives.scala 126:35:@22168.4]
  assign _T_3167 = StickySelects_21_io_outs_2; // @[MemPrimitives.scala 126:35:@22169.4]
  assign _T_3168 = StickySelects_21_io_outs_3; // @[MemPrimitives.scala 126:35:@22170.4]
  assign _T_3169 = StickySelects_21_io_outs_4; // @[MemPrimitives.scala 126:35:@22171.4]
  assign _T_3170 = StickySelects_21_io_outs_5; // @[MemPrimitives.scala 126:35:@22172.4]
  assign _T_3171 = StickySelects_21_io_outs_6; // @[MemPrimitives.scala 126:35:@22173.4]
  assign _T_3172 = StickySelects_21_io_outs_7; // @[MemPrimitives.scala 126:35:@22174.4]
  assign _T_3173 = StickySelects_21_io_outs_8; // @[MemPrimitives.scala 126:35:@22175.4]
  assign _T_3175 = {_T_3165,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22177.4]
  assign _T_3177 = {_T_3166,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22179.4]
  assign _T_3179 = {_T_3167,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22181.4]
  assign _T_3181 = {_T_3168,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22183.4]
  assign _T_3183 = {_T_3169,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22185.4]
  assign _T_3185 = {_T_3170,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22187.4]
  assign _T_3187 = {_T_3171,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22189.4]
  assign _T_3189 = {_T_3172,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22191.4]
  assign _T_3191 = {_T_3173,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22193.4]
  assign _T_3192 = _T_3172 ? _T_3189 : _T_3191; // @[Mux.scala 31:69:@22194.4]
  assign _T_3193 = _T_3171 ? _T_3187 : _T_3192; // @[Mux.scala 31:69:@22195.4]
  assign _T_3194 = _T_3170 ? _T_3185 : _T_3193; // @[Mux.scala 31:69:@22196.4]
  assign _T_3195 = _T_3169 ? _T_3183 : _T_3194; // @[Mux.scala 31:69:@22197.4]
  assign _T_3196 = _T_3168 ? _T_3181 : _T_3195; // @[Mux.scala 31:69:@22198.4]
  assign _T_3197 = _T_3167 ? _T_3179 : _T_3196; // @[Mux.scala 31:69:@22199.4]
  assign _T_3198 = _T_3166 ? _T_3177 : _T_3197; // @[Mux.scala 31:69:@22200.4]
  assign _T_3199 = _T_3165 ? _T_3175 : _T_3198; // @[Mux.scala 31:69:@22201.4]
  assign _T_3207 = _T_2836 & _T_1550; // @[MemPrimitives.scala 110:228:@22210.4]
  assign _T_3213 = _T_2842 & _T_1556; // @[MemPrimitives.scala 110:228:@22214.4]
  assign _T_3219 = _T_2848 & _T_1562; // @[MemPrimitives.scala 110:228:@22218.4]
  assign _T_3225 = _T_2854 & _T_1568; // @[MemPrimitives.scala 110:228:@22222.4]
  assign _T_3231 = _T_2860 & _T_1574; // @[MemPrimitives.scala 110:228:@22226.4]
  assign _T_3237 = _T_2866 & _T_1580; // @[MemPrimitives.scala 110:228:@22230.4]
  assign _T_3243 = _T_2872 & _T_1586; // @[MemPrimitives.scala 110:228:@22234.4]
  assign _T_3249 = _T_2878 & _T_1592; // @[MemPrimitives.scala 110:228:@22238.4]
  assign _T_3255 = _T_2884 & _T_1598; // @[MemPrimitives.scala 110:228:@22242.4]
  assign _T_3257 = StickySelects_22_io_outs_0; // @[MemPrimitives.scala 126:35:@22256.4]
  assign _T_3258 = StickySelects_22_io_outs_1; // @[MemPrimitives.scala 126:35:@22257.4]
  assign _T_3259 = StickySelects_22_io_outs_2; // @[MemPrimitives.scala 126:35:@22258.4]
  assign _T_3260 = StickySelects_22_io_outs_3; // @[MemPrimitives.scala 126:35:@22259.4]
  assign _T_3261 = StickySelects_22_io_outs_4; // @[MemPrimitives.scala 126:35:@22260.4]
  assign _T_3262 = StickySelects_22_io_outs_5; // @[MemPrimitives.scala 126:35:@22261.4]
  assign _T_3263 = StickySelects_22_io_outs_6; // @[MemPrimitives.scala 126:35:@22262.4]
  assign _T_3264 = StickySelects_22_io_outs_7; // @[MemPrimitives.scala 126:35:@22263.4]
  assign _T_3265 = StickySelects_22_io_outs_8; // @[MemPrimitives.scala 126:35:@22264.4]
  assign _T_3267 = {_T_3257,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@22266.4]
  assign _T_3269 = {_T_3258,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@22268.4]
  assign _T_3271 = {_T_3259,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@22270.4]
  assign _T_3273 = {_T_3260,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@22272.4]
  assign _T_3275 = {_T_3261,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@22274.4]
  assign _T_3277 = {_T_3262,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@22276.4]
  assign _T_3279 = {_T_3263,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@22278.4]
  assign _T_3281 = {_T_3264,io_rPort_13_backpressure,io_rPort_13_ofs_0}; // @[Cat.scala 30:58:@22280.4]
  assign _T_3283 = {_T_3265,io_rPort_16_backpressure,io_rPort_16_ofs_0}; // @[Cat.scala 30:58:@22282.4]
  assign _T_3284 = _T_3264 ? _T_3281 : _T_3283; // @[Mux.scala 31:69:@22283.4]
  assign _T_3285 = _T_3263 ? _T_3279 : _T_3284; // @[Mux.scala 31:69:@22284.4]
  assign _T_3286 = _T_3262 ? _T_3277 : _T_3285; // @[Mux.scala 31:69:@22285.4]
  assign _T_3287 = _T_3261 ? _T_3275 : _T_3286; // @[Mux.scala 31:69:@22286.4]
  assign _T_3288 = _T_3260 ? _T_3273 : _T_3287; // @[Mux.scala 31:69:@22287.4]
  assign _T_3289 = _T_3259 ? _T_3271 : _T_3288; // @[Mux.scala 31:69:@22288.4]
  assign _T_3290 = _T_3258 ? _T_3269 : _T_3289; // @[Mux.scala 31:69:@22289.4]
  assign _T_3291 = _T_3257 ? _T_3267 : _T_3290; // @[Mux.scala 31:69:@22290.4]
  assign _T_3299 = _T_2928 & _T_1642; // @[MemPrimitives.scala 110:228:@22299.4]
  assign _T_3305 = _T_2934 & _T_1648; // @[MemPrimitives.scala 110:228:@22303.4]
  assign _T_3311 = _T_2940 & _T_1654; // @[MemPrimitives.scala 110:228:@22307.4]
  assign _T_3317 = _T_2946 & _T_1660; // @[MemPrimitives.scala 110:228:@22311.4]
  assign _T_3323 = _T_2952 & _T_1666; // @[MemPrimitives.scala 110:228:@22315.4]
  assign _T_3329 = _T_2958 & _T_1672; // @[MemPrimitives.scala 110:228:@22319.4]
  assign _T_3335 = _T_2964 & _T_1678; // @[MemPrimitives.scala 110:228:@22323.4]
  assign _T_3341 = _T_2970 & _T_1684; // @[MemPrimitives.scala 110:228:@22327.4]
  assign _T_3347 = _T_2976 & _T_1690; // @[MemPrimitives.scala 110:228:@22331.4]
  assign _T_3349 = StickySelects_23_io_outs_0; // @[MemPrimitives.scala 126:35:@22345.4]
  assign _T_3350 = StickySelects_23_io_outs_1; // @[MemPrimitives.scala 126:35:@22346.4]
  assign _T_3351 = StickySelects_23_io_outs_2; // @[MemPrimitives.scala 126:35:@22347.4]
  assign _T_3352 = StickySelects_23_io_outs_3; // @[MemPrimitives.scala 126:35:@22348.4]
  assign _T_3353 = StickySelects_23_io_outs_4; // @[MemPrimitives.scala 126:35:@22349.4]
  assign _T_3354 = StickySelects_23_io_outs_5; // @[MemPrimitives.scala 126:35:@22350.4]
  assign _T_3355 = StickySelects_23_io_outs_6; // @[MemPrimitives.scala 126:35:@22351.4]
  assign _T_3356 = StickySelects_23_io_outs_7; // @[MemPrimitives.scala 126:35:@22352.4]
  assign _T_3357 = StickySelects_23_io_outs_8; // @[MemPrimitives.scala 126:35:@22353.4]
  assign _T_3359 = {_T_3349,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@22355.4]
  assign _T_3361 = {_T_3350,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@22357.4]
  assign _T_3363 = {_T_3351,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@22359.4]
  assign _T_3365 = {_T_3352,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@22361.4]
  assign _T_3367 = {_T_3353,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@22363.4]
  assign _T_3369 = {_T_3354,io_rPort_12_backpressure,io_rPort_12_ofs_0}; // @[Cat.scala 30:58:@22365.4]
  assign _T_3371 = {_T_3355,io_rPort_14_backpressure,io_rPort_14_ofs_0}; // @[Cat.scala 30:58:@22367.4]
  assign _T_3373 = {_T_3356,io_rPort_15_backpressure,io_rPort_15_ofs_0}; // @[Cat.scala 30:58:@22369.4]
  assign _T_3375 = {_T_3357,io_rPort_17_backpressure,io_rPort_17_ofs_0}; // @[Cat.scala 30:58:@22371.4]
  assign _T_3376 = _T_3356 ? _T_3373 : _T_3375; // @[Mux.scala 31:69:@22372.4]
  assign _T_3377 = _T_3355 ? _T_3371 : _T_3376; // @[Mux.scala 31:69:@22373.4]
  assign _T_3378 = _T_3354 ? _T_3369 : _T_3377; // @[Mux.scala 31:69:@22374.4]
  assign _T_3379 = _T_3353 ? _T_3367 : _T_3378; // @[Mux.scala 31:69:@22375.4]
  assign _T_3380 = _T_3352 ? _T_3365 : _T_3379; // @[Mux.scala 31:69:@22376.4]
  assign _T_3381 = _T_3351 ? _T_3363 : _T_3380; // @[Mux.scala 31:69:@22377.4]
  assign _T_3382 = _T_3350 ? _T_3361 : _T_3381; // @[Mux.scala 31:69:@22378.4]
  assign _T_3383 = _T_3349 ? _T_3359 : _T_3382; // @[Mux.scala 31:69:@22379.4]
  assign _T_3479 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@22508.4 package.scala 96:25:@22509.4]
  assign _T_3483 = _T_3479 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@22518.4]
  assign _T_3476 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@22500.4 package.scala 96:25:@22501.4]
  assign _T_3484 = _T_3476 ? Mem1D_19_io_output : _T_3483; // @[Mux.scala 31:69:@22519.4]
  assign _T_3473 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@22492.4 package.scala 96:25:@22493.4]
  assign _T_3485 = _T_3473 ? Mem1D_17_io_output : _T_3484; // @[Mux.scala 31:69:@22520.4]
  assign _T_3470 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@22484.4 package.scala 96:25:@22485.4]
  assign _T_3486 = _T_3470 ? Mem1D_15_io_output : _T_3485; // @[Mux.scala 31:69:@22521.4]
  assign _T_3467 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@22476.4 package.scala 96:25:@22477.4]
  assign _T_3487 = _T_3467 ? Mem1D_13_io_output : _T_3486; // @[Mux.scala 31:69:@22522.4]
  assign _T_3464 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@22468.4 package.scala 96:25:@22469.4]
  assign _T_3488 = _T_3464 ? Mem1D_11_io_output : _T_3487; // @[Mux.scala 31:69:@22523.4]
  assign _T_3461 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@22460.4 package.scala 96:25:@22461.4]
  assign _T_3489 = _T_3461 ? Mem1D_9_io_output : _T_3488; // @[Mux.scala 31:69:@22524.4]
  assign _T_3458 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@22452.4 package.scala 96:25:@22453.4]
  assign _T_3490 = _T_3458 ? Mem1D_7_io_output : _T_3489; // @[Mux.scala 31:69:@22525.4]
  assign _T_3455 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@22444.4 package.scala 96:25:@22445.4]
  assign _T_3491 = _T_3455 ? Mem1D_5_io_output : _T_3490; // @[Mux.scala 31:69:@22526.4]
  assign _T_3452 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@22436.4 package.scala 96:25:@22437.4]
  assign _T_3492 = _T_3452 ? Mem1D_3_io_output : _T_3491; // @[Mux.scala 31:69:@22527.4]
  assign _T_3449 = RetimeWrapper_io_out; // @[package.scala 96:25:@22428.4 package.scala 96:25:@22429.4]
  assign _T_3586 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@22652.4 package.scala 96:25:@22653.4]
  assign _T_3590 = _T_3586 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@22662.4]
  assign _T_3583 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@22644.4 package.scala 96:25:@22645.4]
  assign _T_3591 = _T_3583 ? Mem1D_18_io_output : _T_3590; // @[Mux.scala 31:69:@22663.4]
  assign _T_3580 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@22636.4 package.scala 96:25:@22637.4]
  assign _T_3592 = _T_3580 ? Mem1D_16_io_output : _T_3591; // @[Mux.scala 31:69:@22664.4]
  assign _T_3577 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@22628.4 package.scala 96:25:@22629.4]
  assign _T_3593 = _T_3577 ? Mem1D_14_io_output : _T_3592; // @[Mux.scala 31:69:@22665.4]
  assign _T_3574 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@22620.4 package.scala 96:25:@22621.4]
  assign _T_3594 = _T_3574 ? Mem1D_12_io_output : _T_3593; // @[Mux.scala 31:69:@22666.4]
  assign _T_3571 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@22612.4 package.scala 96:25:@22613.4]
  assign _T_3595 = _T_3571 ? Mem1D_10_io_output : _T_3594; // @[Mux.scala 31:69:@22667.4]
  assign _T_3568 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@22604.4 package.scala 96:25:@22605.4]
  assign _T_3596 = _T_3568 ? Mem1D_8_io_output : _T_3595; // @[Mux.scala 31:69:@22668.4]
  assign _T_3565 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@22596.4 package.scala 96:25:@22597.4]
  assign _T_3597 = _T_3565 ? Mem1D_6_io_output : _T_3596; // @[Mux.scala 31:69:@22669.4]
  assign _T_3562 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@22588.4 package.scala 96:25:@22589.4]
  assign _T_3598 = _T_3562 ? Mem1D_4_io_output : _T_3597; // @[Mux.scala 31:69:@22670.4]
  assign _T_3559 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@22580.4 package.scala 96:25:@22581.4]
  assign _T_3599 = _T_3559 ? Mem1D_2_io_output : _T_3598; // @[Mux.scala 31:69:@22671.4]
  assign _T_3556 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@22572.4 package.scala 96:25:@22573.4]
  assign _T_3693 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@22796.4 package.scala 96:25:@22797.4]
  assign _T_3697 = _T_3693 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@22806.4]
  assign _T_3690 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@22788.4 package.scala 96:25:@22789.4]
  assign _T_3698 = _T_3690 ? Mem1D_19_io_output : _T_3697; // @[Mux.scala 31:69:@22807.4]
  assign _T_3687 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@22780.4 package.scala 96:25:@22781.4]
  assign _T_3699 = _T_3687 ? Mem1D_17_io_output : _T_3698; // @[Mux.scala 31:69:@22808.4]
  assign _T_3684 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@22772.4 package.scala 96:25:@22773.4]
  assign _T_3700 = _T_3684 ? Mem1D_15_io_output : _T_3699; // @[Mux.scala 31:69:@22809.4]
  assign _T_3681 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@22764.4 package.scala 96:25:@22765.4]
  assign _T_3701 = _T_3681 ? Mem1D_13_io_output : _T_3700; // @[Mux.scala 31:69:@22810.4]
  assign _T_3678 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@22756.4 package.scala 96:25:@22757.4]
  assign _T_3702 = _T_3678 ? Mem1D_11_io_output : _T_3701; // @[Mux.scala 31:69:@22811.4]
  assign _T_3675 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@22748.4 package.scala 96:25:@22749.4]
  assign _T_3703 = _T_3675 ? Mem1D_9_io_output : _T_3702; // @[Mux.scala 31:69:@22812.4]
  assign _T_3672 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@22740.4 package.scala 96:25:@22741.4]
  assign _T_3704 = _T_3672 ? Mem1D_7_io_output : _T_3703; // @[Mux.scala 31:69:@22813.4]
  assign _T_3669 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@22732.4 package.scala 96:25:@22733.4]
  assign _T_3705 = _T_3669 ? Mem1D_5_io_output : _T_3704; // @[Mux.scala 31:69:@22814.4]
  assign _T_3666 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@22724.4 package.scala 96:25:@22725.4]
  assign _T_3706 = _T_3666 ? Mem1D_3_io_output : _T_3705; // @[Mux.scala 31:69:@22815.4]
  assign _T_3663 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@22716.4 package.scala 96:25:@22717.4]
  assign _T_3800 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@22940.4 package.scala 96:25:@22941.4]
  assign _T_3804 = _T_3800 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@22950.4]
  assign _T_3797 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@22932.4 package.scala 96:25:@22933.4]
  assign _T_3805 = _T_3797 ? Mem1D_19_io_output : _T_3804; // @[Mux.scala 31:69:@22951.4]
  assign _T_3794 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@22924.4 package.scala 96:25:@22925.4]
  assign _T_3806 = _T_3794 ? Mem1D_17_io_output : _T_3805; // @[Mux.scala 31:69:@22952.4]
  assign _T_3791 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@22916.4 package.scala 96:25:@22917.4]
  assign _T_3807 = _T_3791 ? Mem1D_15_io_output : _T_3806; // @[Mux.scala 31:69:@22953.4]
  assign _T_3788 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@22908.4 package.scala 96:25:@22909.4]
  assign _T_3808 = _T_3788 ? Mem1D_13_io_output : _T_3807; // @[Mux.scala 31:69:@22954.4]
  assign _T_3785 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@22900.4 package.scala 96:25:@22901.4]
  assign _T_3809 = _T_3785 ? Mem1D_11_io_output : _T_3808; // @[Mux.scala 31:69:@22955.4]
  assign _T_3782 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@22892.4 package.scala 96:25:@22893.4]
  assign _T_3810 = _T_3782 ? Mem1D_9_io_output : _T_3809; // @[Mux.scala 31:69:@22956.4]
  assign _T_3779 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@22884.4 package.scala 96:25:@22885.4]
  assign _T_3811 = _T_3779 ? Mem1D_7_io_output : _T_3810; // @[Mux.scala 31:69:@22957.4]
  assign _T_3776 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@22876.4 package.scala 96:25:@22877.4]
  assign _T_3812 = _T_3776 ? Mem1D_5_io_output : _T_3811; // @[Mux.scala 31:69:@22958.4]
  assign _T_3773 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@22868.4 package.scala 96:25:@22869.4]
  assign _T_3813 = _T_3773 ? Mem1D_3_io_output : _T_3812; // @[Mux.scala 31:69:@22959.4]
  assign _T_3770 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@22860.4 package.scala 96:25:@22861.4]
  assign _T_3907 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@23084.4 package.scala 96:25:@23085.4]
  assign _T_3911 = _T_3907 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23094.4]
  assign _T_3904 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@23076.4 package.scala 96:25:@23077.4]
  assign _T_3912 = _T_3904 ? Mem1D_18_io_output : _T_3911; // @[Mux.scala 31:69:@23095.4]
  assign _T_3901 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@23068.4 package.scala 96:25:@23069.4]
  assign _T_3913 = _T_3901 ? Mem1D_16_io_output : _T_3912; // @[Mux.scala 31:69:@23096.4]
  assign _T_3898 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@23060.4 package.scala 96:25:@23061.4]
  assign _T_3914 = _T_3898 ? Mem1D_14_io_output : _T_3913; // @[Mux.scala 31:69:@23097.4]
  assign _T_3895 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@23052.4 package.scala 96:25:@23053.4]
  assign _T_3915 = _T_3895 ? Mem1D_12_io_output : _T_3914; // @[Mux.scala 31:69:@23098.4]
  assign _T_3892 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@23044.4 package.scala 96:25:@23045.4]
  assign _T_3916 = _T_3892 ? Mem1D_10_io_output : _T_3915; // @[Mux.scala 31:69:@23099.4]
  assign _T_3889 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@23036.4 package.scala 96:25:@23037.4]
  assign _T_3917 = _T_3889 ? Mem1D_8_io_output : _T_3916; // @[Mux.scala 31:69:@23100.4]
  assign _T_3886 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@23028.4 package.scala 96:25:@23029.4]
  assign _T_3918 = _T_3886 ? Mem1D_6_io_output : _T_3917; // @[Mux.scala 31:69:@23101.4]
  assign _T_3883 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@23020.4 package.scala 96:25:@23021.4]
  assign _T_3919 = _T_3883 ? Mem1D_4_io_output : _T_3918; // @[Mux.scala 31:69:@23102.4]
  assign _T_3880 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@23012.4 package.scala 96:25:@23013.4]
  assign _T_3920 = _T_3880 ? Mem1D_2_io_output : _T_3919; // @[Mux.scala 31:69:@23103.4]
  assign _T_3877 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@23004.4 package.scala 96:25:@23005.4]
  assign _T_4014 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@23228.4 package.scala 96:25:@23229.4]
  assign _T_4018 = _T_4014 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23238.4]
  assign _T_4011 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@23220.4 package.scala 96:25:@23221.4]
  assign _T_4019 = _T_4011 ? Mem1D_18_io_output : _T_4018; // @[Mux.scala 31:69:@23239.4]
  assign _T_4008 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@23212.4 package.scala 96:25:@23213.4]
  assign _T_4020 = _T_4008 ? Mem1D_16_io_output : _T_4019; // @[Mux.scala 31:69:@23240.4]
  assign _T_4005 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@23204.4 package.scala 96:25:@23205.4]
  assign _T_4021 = _T_4005 ? Mem1D_14_io_output : _T_4020; // @[Mux.scala 31:69:@23241.4]
  assign _T_4002 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@23196.4 package.scala 96:25:@23197.4]
  assign _T_4022 = _T_4002 ? Mem1D_12_io_output : _T_4021; // @[Mux.scala 31:69:@23242.4]
  assign _T_3999 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@23188.4 package.scala 96:25:@23189.4]
  assign _T_4023 = _T_3999 ? Mem1D_10_io_output : _T_4022; // @[Mux.scala 31:69:@23243.4]
  assign _T_3996 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@23180.4 package.scala 96:25:@23181.4]
  assign _T_4024 = _T_3996 ? Mem1D_8_io_output : _T_4023; // @[Mux.scala 31:69:@23244.4]
  assign _T_3993 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@23172.4 package.scala 96:25:@23173.4]
  assign _T_4025 = _T_3993 ? Mem1D_6_io_output : _T_4024; // @[Mux.scala 31:69:@23245.4]
  assign _T_3990 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@23164.4 package.scala 96:25:@23165.4]
  assign _T_4026 = _T_3990 ? Mem1D_4_io_output : _T_4025; // @[Mux.scala 31:69:@23246.4]
  assign _T_3987 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@23156.4 package.scala 96:25:@23157.4]
  assign _T_4027 = _T_3987 ? Mem1D_2_io_output : _T_4026; // @[Mux.scala 31:69:@23247.4]
  assign _T_3984 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@23148.4 package.scala 96:25:@23149.4]
  assign _T_4121 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@23372.4 package.scala 96:25:@23373.4]
  assign _T_4125 = _T_4121 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23382.4]
  assign _T_4118 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@23364.4 package.scala 96:25:@23365.4]
  assign _T_4126 = _T_4118 ? Mem1D_19_io_output : _T_4125; // @[Mux.scala 31:69:@23383.4]
  assign _T_4115 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@23356.4 package.scala 96:25:@23357.4]
  assign _T_4127 = _T_4115 ? Mem1D_17_io_output : _T_4126; // @[Mux.scala 31:69:@23384.4]
  assign _T_4112 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@23348.4 package.scala 96:25:@23349.4]
  assign _T_4128 = _T_4112 ? Mem1D_15_io_output : _T_4127; // @[Mux.scala 31:69:@23385.4]
  assign _T_4109 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@23340.4 package.scala 96:25:@23341.4]
  assign _T_4129 = _T_4109 ? Mem1D_13_io_output : _T_4128; // @[Mux.scala 31:69:@23386.4]
  assign _T_4106 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@23332.4 package.scala 96:25:@23333.4]
  assign _T_4130 = _T_4106 ? Mem1D_11_io_output : _T_4129; // @[Mux.scala 31:69:@23387.4]
  assign _T_4103 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@23324.4 package.scala 96:25:@23325.4]
  assign _T_4131 = _T_4103 ? Mem1D_9_io_output : _T_4130; // @[Mux.scala 31:69:@23388.4]
  assign _T_4100 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@23316.4 package.scala 96:25:@23317.4]
  assign _T_4132 = _T_4100 ? Mem1D_7_io_output : _T_4131; // @[Mux.scala 31:69:@23389.4]
  assign _T_4097 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@23308.4 package.scala 96:25:@23309.4]
  assign _T_4133 = _T_4097 ? Mem1D_5_io_output : _T_4132; // @[Mux.scala 31:69:@23390.4]
  assign _T_4094 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@23300.4 package.scala 96:25:@23301.4]
  assign _T_4134 = _T_4094 ? Mem1D_3_io_output : _T_4133; // @[Mux.scala 31:69:@23391.4]
  assign _T_4091 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@23292.4 package.scala 96:25:@23293.4]
  assign _T_4228 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@23516.4 package.scala 96:25:@23517.4]
  assign _T_4232 = _T_4228 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23526.4]
  assign _T_4225 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@23508.4 package.scala 96:25:@23509.4]
  assign _T_4233 = _T_4225 ? Mem1D_18_io_output : _T_4232; // @[Mux.scala 31:69:@23527.4]
  assign _T_4222 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@23500.4 package.scala 96:25:@23501.4]
  assign _T_4234 = _T_4222 ? Mem1D_16_io_output : _T_4233; // @[Mux.scala 31:69:@23528.4]
  assign _T_4219 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@23492.4 package.scala 96:25:@23493.4]
  assign _T_4235 = _T_4219 ? Mem1D_14_io_output : _T_4234; // @[Mux.scala 31:69:@23529.4]
  assign _T_4216 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@23484.4 package.scala 96:25:@23485.4]
  assign _T_4236 = _T_4216 ? Mem1D_12_io_output : _T_4235; // @[Mux.scala 31:69:@23530.4]
  assign _T_4213 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@23476.4 package.scala 96:25:@23477.4]
  assign _T_4237 = _T_4213 ? Mem1D_10_io_output : _T_4236; // @[Mux.scala 31:69:@23531.4]
  assign _T_4210 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@23468.4 package.scala 96:25:@23469.4]
  assign _T_4238 = _T_4210 ? Mem1D_8_io_output : _T_4237; // @[Mux.scala 31:69:@23532.4]
  assign _T_4207 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@23460.4 package.scala 96:25:@23461.4]
  assign _T_4239 = _T_4207 ? Mem1D_6_io_output : _T_4238; // @[Mux.scala 31:69:@23533.4]
  assign _T_4204 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@23452.4 package.scala 96:25:@23453.4]
  assign _T_4240 = _T_4204 ? Mem1D_4_io_output : _T_4239; // @[Mux.scala 31:69:@23534.4]
  assign _T_4201 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@23444.4 package.scala 96:25:@23445.4]
  assign _T_4241 = _T_4201 ? Mem1D_2_io_output : _T_4240; // @[Mux.scala 31:69:@23535.4]
  assign _T_4198 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@23436.4 package.scala 96:25:@23437.4]
  assign _T_4335 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@23660.4 package.scala 96:25:@23661.4]
  assign _T_4339 = _T_4335 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23670.4]
  assign _T_4332 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@23652.4 package.scala 96:25:@23653.4]
  assign _T_4340 = _T_4332 ? Mem1D_18_io_output : _T_4339; // @[Mux.scala 31:69:@23671.4]
  assign _T_4329 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@23644.4 package.scala 96:25:@23645.4]
  assign _T_4341 = _T_4329 ? Mem1D_16_io_output : _T_4340; // @[Mux.scala 31:69:@23672.4]
  assign _T_4326 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@23636.4 package.scala 96:25:@23637.4]
  assign _T_4342 = _T_4326 ? Mem1D_14_io_output : _T_4341; // @[Mux.scala 31:69:@23673.4]
  assign _T_4323 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@23628.4 package.scala 96:25:@23629.4]
  assign _T_4343 = _T_4323 ? Mem1D_12_io_output : _T_4342; // @[Mux.scala 31:69:@23674.4]
  assign _T_4320 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@23620.4 package.scala 96:25:@23621.4]
  assign _T_4344 = _T_4320 ? Mem1D_10_io_output : _T_4343; // @[Mux.scala 31:69:@23675.4]
  assign _T_4317 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@23612.4 package.scala 96:25:@23613.4]
  assign _T_4345 = _T_4317 ? Mem1D_8_io_output : _T_4344; // @[Mux.scala 31:69:@23676.4]
  assign _T_4314 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@23604.4 package.scala 96:25:@23605.4]
  assign _T_4346 = _T_4314 ? Mem1D_6_io_output : _T_4345; // @[Mux.scala 31:69:@23677.4]
  assign _T_4311 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@23596.4 package.scala 96:25:@23597.4]
  assign _T_4347 = _T_4311 ? Mem1D_4_io_output : _T_4346; // @[Mux.scala 31:69:@23678.4]
  assign _T_4308 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@23588.4 package.scala 96:25:@23589.4]
  assign _T_4348 = _T_4308 ? Mem1D_2_io_output : _T_4347; // @[Mux.scala 31:69:@23679.4]
  assign _T_4305 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@23580.4 package.scala 96:25:@23581.4]
  assign _T_4442 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@23804.4 package.scala 96:25:@23805.4]
  assign _T_4446 = _T_4442 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@23814.4]
  assign _T_4439 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@23796.4 package.scala 96:25:@23797.4]
  assign _T_4447 = _T_4439 ? Mem1D_19_io_output : _T_4446; // @[Mux.scala 31:69:@23815.4]
  assign _T_4436 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@23788.4 package.scala 96:25:@23789.4]
  assign _T_4448 = _T_4436 ? Mem1D_17_io_output : _T_4447; // @[Mux.scala 31:69:@23816.4]
  assign _T_4433 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@23780.4 package.scala 96:25:@23781.4]
  assign _T_4449 = _T_4433 ? Mem1D_15_io_output : _T_4448; // @[Mux.scala 31:69:@23817.4]
  assign _T_4430 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@23772.4 package.scala 96:25:@23773.4]
  assign _T_4450 = _T_4430 ? Mem1D_13_io_output : _T_4449; // @[Mux.scala 31:69:@23818.4]
  assign _T_4427 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@23764.4 package.scala 96:25:@23765.4]
  assign _T_4451 = _T_4427 ? Mem1D_11_io_output : _T_4450; // @[Mux.scala 31:69:@23819.4]
  assign _T_4424 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@23756.4 package.scala 96:25:@23757.4]
  assign _T_4452 = _T_4424 ? Mem1D_9_io_output : _T_4451; // @[Mux.scala 31:69:@23820.4]
  assign _T_4421 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@23748.4 package.scala 96:25:@23749.4]
  assign _T_4453 = _T_4421 ? Mem1D_7_io_output : _T_4452; // @[Mux.scala 31:69:@23821.4]
  assign _T_4418 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@23740.4 package.scala 96:25:@23741.4]
  assign _T_4454 = _T_4418 ? Mem1D_5_io_output : _T_4453; // @[Mux.scala 31:69:@23822.4]
  assign _T_4415 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@23732.4 package.scala 96:25:@23733.4]
  assign _T_4455 = _T_4415 ? Mem1D_3_io_output : _T_4454; // @[Mux.scala 31:69:@23823.4]
  assign _T_4412 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@23724.4 package.scala 96:25:@23725.4]
  assign _T_4549 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@23948.4 package.scala 96:25:@23949.4]
  assign _T_4553 = _T_4549 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@23958.4]
  assign _T_4546 = RetimeWrapper_129_io_out; // @[package.scala 96:25:@23940.4 package.scala 96:25:@23941.4]
  assign _T_4554 = _T_4546 ? Mem1D_18_io_output : _T_4553; // @[Mux.scala 31:69:@23959.4]
  assign _T_4543 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@23932.4 package.scala 96:25:@23933.4]
  assign _T_4555 = _T_4543 ? Mem1D_16_io_output : _T_4554; // @[Mux.scala 31:69:@23960.4]
  assign _T_4540 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@23924.4 package.scala 96:25:@23925.4]
  assign _T_4556 = _T_4540 ? Mem1D_14_io_output : _T_4555; // @[Mux.scala 31:69:@23961.4]
  assign _T_4537 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@23916.4 package.scala 96:25:@23917.4]
  assign _T_4557 = _T_4537 ? Mem1D_12_io_output : _T_4556; // @[Mux.scala 31:69:@23962.4]
  assign _T_4534 = RetimeWrapper_125_io_out; // @[package.scala 96:25:@23908.4 package.scala 96:25:@23909.4]
  assign _T_4558 = _T_4534 ? Mem1D_10_io_output : _T_4557; // @[Mux.scala 31:69:@23963.4]
  assign _T_4531 = RetimeWrapper_124_io_out; // @[package.scala 96:25:@23900.4 package.scala 96:25:@23901.4]
  assign _T_4559 = _T_4531 ? Mem1D_8_io_output : _T_4558; // @[Mux.scala 31:69:@23964.4]
  assign _T_4528 = RetimeWrapper_123_io_out; // @[package.scala 96:25:@23892.4 package.scala 96:25:@23893.4]
  assign _T_4560 = _T_4528 ? Mem1D_6_io_output : _T_4559; // @[Mux.scala 31:69:@23965.4]
  assign _T_4525 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@23884.4 package.scala 96:25:@23885.4]
  assign _T_4561 = _T_4525 ? Mem1D_4_io_output : _T_4560; // @[Mux.scala 31:69:@23966.4]
  assign _T_4522 = RetimeWrapper_121_io_out; // @[package.scala 96:25:@23876.4 package.scala 96:25:@23877.4]
  assign _T_4562 = _T_4522 ? Mem1D_2_io_output : _T_4561; // @[Mux.scala 31:69:@23967.4]
  assign _T_4519 = RetimeWrapper_120_io_out; // @[package.scala 96:25:@23868.4 package.scala 96:25:@23869.4]
  assign _T_4656 = RetimeWrapper_142_io_out; // @[package.scala 96:25:@24092.4 package.scala 96:25:@24093.4]
  assign _T_4660 = _T_4656 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24102.4]
  assign _T_4653 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@24084.4 package.scala 96:25:@24085.4]
  assign _T_4661 = _T_4653 ? Mem1D_18_io_output : _T_4660; // @[Mux.scala 31:69:@24103.4]
  assign _T_4650 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@24076.4 package.scala 96:25:@24077.4]
  assign _T_4662 = _T_4650 ? Mem1D_16_io_output : _T_4661; // @[Mux.scala 31:69:@24104.4]
  assign _T_4647 = RetimeWrapper_139_io_out; // @[package.scala 96:25:@24068.4 package.scala 96:25:@24069.4]
  assign _T_4663 = _T_4647 ? Mem1D_14_io_output : _T_4662; // @[Mux.scala 31:69:@24105.4]
  assign _T_4644 = RetimeWrapper_138_io_out; // @[package.scala 96:25:@24060.4 package.scala 96:25:@24061.4]
  assign _T_4664 = _T_4644 ? Mem1D_12_io_output : _T_4663; // @[Mux.scala 31:69:@24106.4]
  assign _T_4641 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@24052.4 package.scala 96:25:@24053.4]
  assign _T_4665 = _T_4641 ? Mem1D_10_io_output : _T_4664; // @[Mux.scala 31:69:@24107.4]
  assign _T_4638 = RetimeWrapper_136_io_out; // @[package.scala 96:25:@24044.4 package.scala 96:25:@24045.4]
  assign _T_4666 = _T_4638 ? Mem1D_8_io_output : _T_4665; // @[Mux.scala 31:69:@24108.4]
  assign _T_4635 = RetimeWrapper_135_io_out; // @[package.scala 96:25:@24036.4 package.scala 96:25:@24037.4]
  assign _T_4667 = _T_4635 ? Mem1D_6_io_output : _T_4666; // @[Mux.scala 31:69:@24109.4]
  assign _T_4632 = RetimeWrapper_134_io_out; // @[package.scala 96:25:@24028.4 package.scala 96:25:@24029.4]
  assign _T_4668 = _T_4632 ? Mem1D_4_io_output : _T_4667; // @[Mux.scala 31:69:@24110.4]
  assign _T_4629 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@24020.4 package.scala 96:25:@24021.4]
  assign _T_4669 = _T_4629 ? Mem1D_2_io_output : _T_4668; // @[Mux.scala 31:69:@24111.4]
  assign _T_4626 = RetimeWrapper_132_io_out; // @[package.scala 96:25:@24012.4 package.scala 96:25:@24013.4]
  assign _T_4763 = RetimeWrapper_154_io_out; // @[package.scala 96:25:@24236.4 package.scala 96:25:@24237.4]
  assign _T_4767 = _T_4763 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24246.4]
  assign _T_4760 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@24228.4 package.scala 96:25:@24229.4]
  assign _T_4768 = _T_4760 ? Mem1D_19_io_output : _T_4767; // @[Mux.scala 31:69:@24247.4]
  assign _T_4757 = RetimeWrapper_152_io_out; // @[package.scala 96:25:@24220.4 package.scala 96:25:@24221.4]
  assign _T_4769 = _T_4757 ? Mem1D_17_io_output : _T_4768; // @[Mux.scala 31:69:@24248.4]
  assign _T_4754 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@24212.4 package.scala 96:25:@24213.4]
  assign _T_4770 = _T_4754 ? Mem1D_15_io_output : _T_4769; // @[Mux.scala 31:69:@24249.4]
  assign _T_4751 = RetimeWrapper_150_io_out; // @[package.scala 96:25:@24204.4 package.scala 96:25:@24205.4]
  assign _T_4771 = _T_4751 ? Mem1D_13_io_output : _T_4770; // @[Mux.scala 31:69:@24250.4]
  assign _T_4748 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@24196.4 package.scala 96:25:@24197.4]
  assign _T_4772 = _T_4748 ? Mem1D_11_io_output : _T_4771; // @[Mux.scala 31:69:@24251.4]
  assign _T_4745 = RetimeWrapper_148_io_out; // @[package.scala 96:25:@24188.4 package.scala 96:25:@24189.4]
  assign _T_4773 = _T_4745 ? Mem1D_9_io_output : _T_4772; // @[Mux.scala 31:69:@24252.4]
  assign _T_4742 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@24180.4 package.scala 96:25:@24181.4]
  assign _T_4774 = _T_4742 ? Mem1D_7_io_output : _T_4773; // @[Mux.scala 31:69:@24253.4]
  assign _T_4739 = RetimeWrapper_146_io_out; // @[package.scala 96:25:@24172.4 package.scala 96:25:@24173.4]
  assign _T_4775 = _T_4739 ? Mem1D_5_io_output : _T_4774; // @[Mux.scala 31:69:@24254.4]
  assign _T_4736 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@24164.4 package.scala 96:25:@24165.4]
  assign _T_4776 = _T_4736 ? Mem1D_3_io_output : _T_4775; // @[Mux.scala 31:69:@24255.4]
  assign _T_4733 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@24156.4 package.scala 96:25:@24157.4]
  assign _T_4870 = RetimeWrapper_166_io_out; // @[package.scala 96:25:@24380.4 package.scala 96:25:@24381.4]
  assign _T_4874 = _T_4870 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24390.4]
  assign _T_4867 = RetimeWrapper_165_io_out; // @[package.scala 96:25:@24372.4 package.scala 96:25:@24373.4]
  assign _T_4875 = _T_4867 ? Mem1D_18_io_output : _T_4874; // @[Mux.scala 31:69:@24391.4]
  assign _T_4864 = RetimeWrapper_164_io_out; // @[package.scala 96:25:@24364.4 package.scala 96:25:@24365.4]
  assign _T_4876 = _T_4864 ? Mem1D_16_io_output : _T_4875; // @[Mux.scala 31:69:@24392.4]
  assign _T_4861 = RetimeWrapper_163_io_out; // @[package.scala 96:25:@24356.4 package.scala 96:25:@24357.4]
  assign _T_4877 = _T_4861 ? Mem1D_14_io_output : _T_4876; // @[Mux.scala 31:69:@24393.4]
  assign _T_4858 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@24348.4 package.scala 96:25:@24349.4]
  assign _T_4878 = _T_4858 ? Mem1D_12_io_output : _T_4877; // @[Mux.scala 31:69:@24394.4]
  assign _T_4855 = RetimeWrapper_161_io_out; // @[package.scala 96:25:@24340.4 package.scala 96:25:@24341.4]
  assign _T_4879 = _T_4855 ? Mem1D_10_io_output : _T_4878; // @[Mux.scala 31:69:@24395.4]
  assign _T_4852 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@24332.4 package.scala 96:25:@24333.4]
  assign _T_4880 = _T_4852 ? Mem1D_8_io_output : _T_4879; // @[Mux.scala 31:69:@24396.4]
  assign _T_4849 = RetimeWrapper_159_io_out; // @[package.scala 96:25:@24324.4 package.scala 96:25:@24325.4]
  assign _T_4881 = _T_4849 ? Mem1D_6_io_output : _T_4880; // @[Mux.scala 31:69:@24397.4]
  assign _T_4846 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@24316.4 package.scala 96:25:@24317.4]
  assign _T_4882 = _T_4846 ? Mem1D_4_io_output : _T_4881; // @[Mux.scala 31:69:@24398.4]
  assign _T_4843 = RetimeWrapper_157_io_out; // @[package.scala 96:25:@24308.4 package.scala 96:25:@24309.4]
  assign _T_4883 = _T_4843 ? Mem1D_2_io_output : _T_4882; // @[Mux.scala 31:69:@24399.4]
  assign _T_4840 = RetimeWrapper_156_io_out; // @[package.scala 96:25:@24300.4 package.scala 96:25:@24301.4]
  assign _T_4977 = RetimeWrapper_178_io_out; // @[package.scala 96:25:@24524.4 package.scala 96:25:@24525.4]
  assign _T_4981 = _T_4977 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24534.4]
  assign _T_4974 = RetimeWrapper_177_io_out; // @[package.scala 96:25:@24516.4 package.scala 96:25:@24517.4]
  assign _T_4982 = _T_4974 ? Mem1D_19_io_output : _T_4981; // @[Mux.scala 31:69:@24535.4]
  assign _T_4971 = RetimeWrapper_176_io_out; // @[package.scala 96:25:@24508.4 package.scala 96:25:@24509.4]
  assign _T_4983 = _T_4971 ? Mem1D_17_io_output : _T_4982; // @[Mux.scala 31:69:@24536.4]
  assign _T_4968 = RetimeWrapper_175_io_out; // @[package.scala 96:25:@24500.4 package.scala 96:25:@24501.4]
  assign _T_4984 = _T_4968 ? Mem1D_15_io_output : _T_4983; // @[Mux.scala 31:69:@24537.4]
  assign _T_4965 = RetimeWrapper_174_io_out; // @[package.scala 96:25:@24492.4 package.scala 96:25:@24493.4]
  assign _T_4985 = _T_4965 ? Mem1D_13_io_output : _T_4984; // @[Mux.scala 31:69:@24538.4]
  assign _T_4962 = RetimeWrapper_173_io_out; // @[package.scala 96:25:@24484.4 package.scala 96:25:@24485.4]
  assign _T_4986 = _T_4962 ? Mem1D_11_io_output : _T_4985; // @[Mux.scala 31:69:@24539.4]
  assign _T_4959 = RetimeWrapper_172_io_out; // @[package.scala 96:25:@24476.4 package.scala 96:25:@24477.4]
  assign _T_4987 = _T_4959 ? Mem1D_9_io_output : _T_4986; // @[Mux.scala 31:69:@24540.4]
  assign _T_4956 = RetimeWrapper_171_io_out; // @[package.scala 96:25:@24468.4 package.scala 96:25:@24469.4]
  assign _T_4988 = _T_4956 ? Mem1D_7_io_output : _T_4987; // @[Mux.scala 31:69:@24541.4]
  assign _T_4953 = RetimeWrapper_170_io_out; // @[package.scala 96:25:@24460.4 package.scala 96:25:@24461.4]
  assign _T_4989 = _T_4953 ? Mem1D_5_io_output : _T_4988; // @[Mux.scala 31:69:@24542.4]
  assign _T_4950 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@24452.4 package.scala 96:25:@24453.4]
  assign _T_4990 = _T_4950 ? Mem1D_3_io_output : _T_4989; // @[Mux.scala 31:69:@24543.4]
  assign _T_4947 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@24444.4 package.scala 96:25:@24445.4]
  assign _T_5084 = RetimeWrapper_190_io_out; // @[package.scala 96:25:@24668.4 package.scala 96:25:@24669.4]
  assign _T_5088 = _T_5084 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24678.4]
  assign _T_5081 = RetimeWrapper_189_io_out; // @[package.scala 96:25:@24660.4 package.scala 96:25:@24661.4]
  assign _T_5089 = _T_5081 ? Mem1D_19_io_output : _T_5088; // @[Mux.scala 31:69:@24679.4]
  assign _T_5078 = RetimeWrapper_188_io_out; // @[package.scala 96:25:@24652.4 package.scala 96:25:@24653.4]
  assign _T_5090 = _T_5078 ? Mem1D_17_io_output : _T_5089; // @[Mux.scala 31:69:@24680.4]
  assign _T_5075 = RetimeWrapper_187_io_out; // @[package.scala 96:25:@24644.4 package.scala 96:25:@24645.4]
  assign _T_5091 = _T_5075 ? Mem1D_15_io_output : _T_5090; // @[Mux.scala 31:69:@24681.4]
  assign _T_5072 = RetimeWrapper_186_io_out; // @[package.scala 96:25:@24636.4 package.scala 96:25:@24637.4]
  assign _T_5092 = _T_5072 ? Mem1D_13_io_output : _T_5091; // @[Mux.scala 31:69:@24682.4]
  assign _T_5069 = RetimeWrapper_185_io_out; // @[package.scala 96:25:@24628.4 package.scala 96:25:@24629.4]
  assign _T_5093 = _T_5069 ? Mem1D_11_io_output : _T_5092; // @[Mux.scala 31:69:@24683.4]
  assign _T_5066 = RetimeWrapper_184_io_out; // @[package.scala 96:25:@24620.4 package.scala 96:25:@24621.4]
  assign _T_5094 = _T_5066 ? Mem1D_9_io_output : _T_5093; // @[Mux.scala 31:69:@24684.4]
  assign _T_5063 = RetimeWrapper_183_io_out; // @[package.scala 96:25:@24612.4 package.scala 96:25:@24613.4]
  assign _T_5095 = _T_5063 ? Mem1D_7_io_output : _T_5094; // @[Mux.scala 31:69:@24685.4]
  assign _T_5060 = RetimeWrapper_182_io_out; // @[package.scala 96:25:@24604.4 package.scala 96:25:@24605.4]
  assign _T_5096 = _T_5060 ? Mem1D_5_io_output : _T_5095; // @[Mux.scala 31:69:@24686.4]
  assign _T_5057 = RetimeWrapper_181_io_out; // @[package.scala 96:25:@24596.4 package.scala 96:25:@24597.4]
  assign _T_5097 = _T_5057 ? Mem1D_3_io_output : _T_5096; // @[Mux.scala 31:69:@24687.4]
  assign _T_5054 = RetimeWrapper_180_io_out; // @[package.scala 96:25:@24588.4 package.scala 96:25:@24589.4]
  assign _T_5191 = RetimeWrapper_202_io_out; // @[package.scala 96:25:@24812.4 package.scala 96:25:@24813.4]
  assign _T_5195 = _T_5191 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@24822.4]
  assign _T_5188 = RetimeWrapper_201_io_out; // @[package.scala 96:25:@24804.4 package.scala 96:25:@24805.4]
  assign _T_5196 = _T_5188 ? Mem1D_18_io_output : _T_5195; // @[Mux.scala 31:69:@24823.4]
  assign _T_5185 = RetimeWrapper_200_io_out; // @[package.scala 96:25:@24796.4 package.scala 96:25:@24797.4]
  assign _T_5197 = _T_5185 ? Mem1D_16_io_output : _T_5196; // @[Mux.scala 31:69:@24824.4]
  assign _T_5182 = RetimeWrapper_199_io_out; // @[package.scala 96:25:@24788.4 package.scala 96:25:@24789.4]
  assign _T_5198 = _T_5182 ? Mem1D_14_io_output : _T_5197; // @[Mux.scala 31:69:@24825.4]
  assign _T_5179 = RetimeWrapper_198_io_out; // @[package.scala 96:25:@24780.4 package.scala 96:25:@24781.4]
  assign _T_5199 = _T_5179 ? Mem1D_12_io_output : _T_5198; // @[Mux.scala 31:69:@24826.4]
  assign _T_5176 = RetimeWrapper_197_io_out; // @[package.scala 96:25:@24772.4 package.scala 96:25:@24773.4]
  assign _T_5200 = _T_5176 ? Mem1D_10_io_output : _T_5199; // @[Mux.scala 31:69:@24827.4]
  assign _T_5173 = RetimeWrapper_196_io_out; // @[package.scala 96:25:@24764.4 package.scala 96:25:@24765.4]
  assign _T_5201 = _T_5173 ? Mem1D_8_io_output : _T_5200; // @[Mux.scala 31:69:@24828.4]
  assign _T_5170 = RetimeWrapper_195_io_out; // @[package.scala 96:25:@24756.4 package.scala 96:25:@24757.4]
  assign _T_5202 = _T_5170 ? Mem1D_6_io_output : _T_5201; // @[Mux.scala 31:69:@24829.4]
  assign _T_5167 = RetimeWrapper_194_io_out; // @[package.scala 96:25:@24748.4 package.scala 96:25:@24749.4]
  assign _T_5203 = _T_5167 ? Mem1D_4_io_output : _T_5202; // @[Mux.scala 31:69:@24830.4]
  assign _T_5164 = RetimeWrapper_193_io_out; // @[package.scala 96:25:@24740.4 package.scala 96:25:@24741.4]
  assign _T_5204 = _T_5164 ? Mem1D_2_io_output : _T_5203; // @[Mux.scala 31:69:@24831.4]
  assign _T_5161 = RetimeWrapper_192_io_out; // @[package.scala 96:25:@24732.4 package.scala 96:25:@24733.4]
  assign _T_5298 = RetimeWrapper_214_io_out; // @[package.scala 96:25:@24956.4 package.scala 96:25:@24957.4]
  assign _T_5302 = _T_5298 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@24966.4]
  assign _T_5295 = RetimeWrapper_213_io_out; // @[package.scala 96:25:@24948.4 package.scala 96:25:@24949.4]
  assign _T_5303 = _T_5295 ? Mem1D_19_io_output : _T_5302; // @[Mux.scala 31:69:@24967.4]
  assign _T_5292 = RetimeWrapper_212_io_out; // @[package.scala 96:25:@24940.4 package.scala 96:25:@24941.4]
  assign _T_5304 = _T_5292 ? Mem1D_17_io_output : _T_5303; // @[Mux.scala 31:69:@24968.4]
  assign _T_5289 = RetimeWrapper_211_io_out; // @[package.scala 96:25:@24932.4 package.scala 96:25:@24933.4]
  assign _T_5305 = _T_5289 ? Mem1D_15_io_output : _T_5304; // @[Mux.scala 31:69:@24969.4]
  assign _T_5286 = RetimeWrapper_210_io_out; // @[package.scala 96:25:@24924.4 package.scala 96:25:@24925.4]
  assign _T_5306 = _T_5286 ? Mem1D_13_io_output : _T_5305; // @[Mux.scala 31:69:@24970.4]
  assign _T_5283 = RetimeWrapper_209_io_out; // @[package.scala 96:25:@24916.4 package.scala 96:25:@24917.4]
  assign _T_5307 = _T_5283 ? Mem1D_11_io_output : _T_5306; // @[Mux.scala 31:69:@24971.4]
  assign _T_5280 = RetimeWrapper_208_io_out; // @[package.scala 96:25:@24908.4 package.scala 96:25:@24909.4]
  assign _T_5308 = _T_5280 ? Mem1D_9_io_output : _T_5307; // @[Mux.scala 31:69:@24972.4]
  assign _T_5277 = RetimeWrapper_207_io_out; // @[package.scala 96:25:@24900.4 package.scala 96:25:@24901.4]
  assign _T_5309 = _T_5277 ? Mem1D_7_io_output : _T_5308; // @[Mux.scala 31:69:@24973.4]
  assign _T_5274 = RetimeWrapper_206_io_out; // @[package.scala 96:25:@24892.4 package.scala 96:25:@24893.4]
  assign _T_5310 = _T_5274 ? Mem1D_5_io_output : _T_5309; // @[Mux.scala 31:69:@24974.4]
  assign _T_5271 = RetimeWrapper_205_io_out; // @[package.scala 96:25:@24884.4 package.scala 96:25:@24885.4]
  assign _T_5311 = _T_5271 ? Mem1D_3_io_output : _T_5310; // @[Mux.scala 31:69:@24975.4]
  assign _T_5268 = RetimeWrapper_204_io_out; // @[package.scala 96:25:@24876.4 package.scala 96:25:@24877.4]
  assign io_rPort_17_output_0 = _T_5268 ? Mem1D_1_io_output : _T_5311; // @[MemPrimitives.scala 152:13:@24977.4]
  assign io_rPort_16_output_0 = _T_5161 ? Mem1D_io_output : _T_5204; // @[MemPrimitives.scala 152:13:@24833.4]
  assign io_rPort_15_output_0 = _T_5054 ? Mem1D_1_io_output : _T_5097; // @[MemPrimitives.scala 152:13:@24689.4]
  assign io_rPort_14_output_0 = _T_4947 ? Mem1D_1_io_output : _T_4990; // @[MemPrimitives.scala 152:13:@24545.4]
  assign io_rPort_13_output_0 = _T_4840 ? Mem1D_io_output : _T_4883; // @[MemPrimitives.scala 152:13:@24401.4]
  assign io_rPort_12_output_0 = _T_4733 ? Mem1D_1_io_output : _T_4776; // @[MemPrimitives.scala 152:13:@24257.4]
  assign io_rPort_11_output_0 = _T_4626 ? Mem1D_io_output : _T_4669; // @[MemPrimitives.scala 152:13:@24113.4]
  assign io_rPort_10_output_0 = _T_4519 ? Mem1D_io_output : _T_4562; // @[MemPrimitives.scala 152:13:@23969.4]
  assign io_rPort_9_output_0 = _T_4412 ? Mem1D_1_io_output : _T_4455; // @[MemPrimitives.scala 152:13:@23825.4]
  assign io_rPort_8_output_0 = _T_4305 ? Mem1D_io_output : _T_4348; // @[MemPrimitives.scala 152:13:@23681.4]
  assign io_rPort_7_output_0 = _T_4198 ? Mem1D_io_output : _T_4241; // @[MemPrimitives.scala 152:13:@23537.4]
  assign io_rPort_6_output_0 = _T_4091 ? Mem1D_1_io_output : _T_4134; // @[MemPrimitives.scala 152:13:@23393.4]
  assign io_rPort_5_output_0 = _T_3984 ? Mem1D_io_output : _T_4027; // @[MemPrimitives.scala 152:13:@23249.4]
  assign io_rPort_4_output_0 = _T_3877 ? Mem1D_io_output : _T_3920; // @[MemPrimitives.scala 152:13:@23105.4]
  assign io_rPort_3_output_0 = _T_3770 ? Mem1D_1_io_output : _T_3813; // @[MemPrimitives.scala 152:13:@22961.4]
  assign io_rPort_2_output_0 = _T_3663 ? Mem1D_1_io_output : _T_3706; // @[MemPrimitives.scala 152:13:@22817.4]
  assign io_rPort_1_output_0 = _T_3556 ? Mem1D_io_output : _T_3599; // @[MemPrimitives.scala 152:13:@22673.4]
  assign io_rPort_0_output_0 = _T_3449 ? Mem1D_1_io_output : _T_3492; // @[MemPrimitives.scala 152:13:@22529.4]
  assign Mem1D_clock = clock; // @[:@19411.4]
  assign Mem1D_reset = reset; // @[:@19412.4]
  assign Mem1D_io_r_ofs_0 = _T_1267[8:0]; // @[MemPrimitives.scala 131:28:@20336.4]
  assign Mem1D_io_r_backpressure = _T_1267[9]; // @[MemPrimitives.scala 132:32:@20337.4]
  assign Mem1D_io_w_ofs_0 = _T_715[8:0]; // @[MemPrimitives.scala 94:28:@19810.4]
  assign Mem1D_io_w_data_0 = _T_715[40:9]; // @[MemPrimitives.scala 95:29:@19811.4]
  assign Mem1D_io_w_en_0 = _T_715[41]; // @[MemPrimitives.scala 96:27:@19812.4]
  assign Mem1D_1_clock = clock; // @[:@19427.4]
  assign Mem1D_1_reset = reset; // @[:@19428.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 131:28:@20425.4]
  assign Mem1D_1_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 132:32:@20426.4]
  assign Mem1D_1_io_w_ofs_0 = _T_735[8:0]; // @[MemPrimitives.scala 94:28:@19829.4]
  assign Mem1D_1_io_w_data_0 = _T_735[40:9]; // @[MemPrimitives.scala 95:29:@19830.4]
  assign Mem1D_1_io_w_en_0 = _T_735[41]; // @[MemPrimitives.scala 96:27:@19831.4]
  assign Mem1D_2_clock = clock; // @[:@19443.4]
  assign Mem1D_2_reset = reset; // @[:@19444.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1451[8:0]; // @[MemPrimitives.scala 131:28:@20514.4]
  assign Mem1D_2_io_r_backpressure = _T_1451[9]; // @[MemPrimitives.scala 132:32:@20515.4]
  assign Mem1D_2_io_w_ofs_0 = _T_755[8:0]; // @[MemPrimitives.scala 94:28:@19848.4]
  assign Mem1D_2_io_w_data_0 = _T_755[40:9]; // @[MemPrimitives.scala 95:29:@19849.4]
  assign Mem1D_2_io_w_en_0 = _T_755[41]; // @[MemPrimitives.scala 96:27:@19850.4]
  assign Mem1D_3_clock = clock; // @[:@19459.4]
  assign Mem1D_3_reset = reset; // @[:@19460.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1543[8:0]; // @[MemPrimitives.scala 131:28:@20603.4]
  assign Mem1D_3_io_r_backpressure = _T_1543[9]; // @[MemPrimitives.scala 132:32:@20604.4]
  assign Mem1D_3_io_w_ofs_0 = _T_775[8:0]; // @[MemPrimitives.scala 94:28:@19867.4]
  assign Mem1D_3_io_w_data_0 = _T_775[40:9]; // @[MemPrimitives.scala 95:29:@19868.4]
  assign Mem1D_3_io_w_en_0 = _T_775[41]; // @[MemPrimitives.scala 96:27:@19869.4]
  assign Mem1D_4_clock = clock; // @[:@19475.4]
  assign Mem1D_4_reset = reset; // @[:@19476.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1635[8:0]; // @[MemPrimitives.scala 131:28:@20692.4]
  assign Mem1D_4_io_r_backpressure = _T_1635[9]; // @[MemPrimitives.scala 132:32:@20693.4]
  assign Mem1D_4_io_w_ofs_0 = _T_795[8:0]; // @[MemPrimitives.scala 94:28:@19886.4]
  assign Mem1D_4_io_w_data_0 = _T_795[40:9]; // @[MemPrimitives.scala 95:29:@19887.4]
  assign Mem1D_4_io_w_en_0 = _T_795[41]; // @[MemPrimitives.scala 96:27:@19888.4]
  assign Mem1D_5_clock = clock; // @[:@19491.4]
  assign Mem1D_5_reset = reset; // @[:@19492.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1727[8:0]; // @[MemPrimitives.scala 131:28:@20781.4]
  assign Mem1D_5_io_r_backpressure = _T_1727[9]; // @[MemPrimitives.scala 132:32:@20782.4]
  assign Mem1D_5_io_w_ofs_0 = _T_815[8:0]; // @[MemPrimitives.scala 94:28:@19905.4]
  assign Mem1D_5_io_w_data_0 = _T_815[40:9]; // @[MemPrimitives.scala 95:29:@19906.4]
  assign Mem1D_5_io_w_en_0 = _T_815[41]; // @[MemPrimitives.scala 96:27:@19907.4]
  assign Mem1D_6_clock = clock; // @[:@19507.4]
  assign Mem1D_6_reset = reset; // @[:@19508.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1819[8:0]; // @[MemPrimitives.scala 131:28:@20870.4]
  assign Mem1D_6_io_r_backpressure = _T_1819[9]; // @[MemPrimitives.scala 132:32:@20871.4]
  assign Mem1D_6_io_w_ofs_0 = _T_835[8:0]; // @[MemPrimitives.scala 94:28:@19924.4]
  assign Mem1D_6_io_w_data_0 = _T_835[40:9]; // @[MemPrimitives.scala 95:29:@19925.4]
  assign Mem1D_6_io_w_en_0 = _T_835[41]; // @[MemPrimitives.scala 96:27:@19926.4]
  assign Mem1D_7_clock = clock; // @[:@19523.4]
  assign Mem1D_7_reset = reset; // @[:@19524.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1911[8:0]; // @[MemPrimitives.scala 131:28:@20959.4]
  assign Mem1D_7_io_r_backpressure = _T_1911[9]; // @[MemPrimitives.scala 132:32:@20960.4]
  assign Mem1D_7_io_w_ofs_0 = _T_855[8:0]; // @[MemPrimitives.scala 94:28:@19943.4]
  assign Mem1D_7_io_w_data_0 = _T_855[40:9]; // @[MemPrimitives.scala 95:29:@19944.4]
  assign Mem1D_7_io_w_en_0 = _T_855[41]; // @[MemPrimitives.scala 96:27:@19945.4]
  assign Mem1D_8_clock = clock; // @[:@19539.4]
  assign Mem1D_8_reset = reset; // @[:@19540.4]
  assign Mem1D_8_io_r_ofs_0 = _T_2003[8:0]; // @[MemPrimitives.scala 131:28:@21048.4]
  assign Mem1D_8_io_r_backpressure = _T_2003[9]; // @[MemPrimitives.scala 132:32:@21049.4]
  assign Mem1D_8_io_w_ofs_0 = _T_875[8:0]; // @[MemPrimitives.scala 94:28:@19962.4]
  assign Mem1D_8_io_w_data_0 = _T_875[40:9]; // @[MemPrimitives.scala 95:29:@19963.4]
  assign Mem1D_8_io_w_en_0 = _T_875[41]; // @[MemPrimitives.scala 96:27:@19964.4]
  assign Mem1D_9_clock = clock; // @[:@19555.4]
  assign Mem1D_9_reset = reset; // @[:@19556.4]
  assign Mem1D_9_io_r_ofs_0 = _T_2095[8:0]; // @[MemPrimitives.scala 131:28:@21137.4]
  assign Mem1D_9_io_r_backpressure = _T_2095[9]; // @[MemPrimitives.scala 132:32:@21138.4]
  assign Mem1D_9_io_w_ofs_0 = _T_895[8:0]; // @[MemPrimitives.scala 94:28:@19981.4]
  assign Mem1D_9_io_w_data_0 = _T_895[40:9]; // @[MemPrimitives.scala 95:29:@19982.4]
  assign Mem1D_9_io_w_en_0 = _T_895[41]; // @[MemPrimitives.scala 96:27:@19983.4]
  assign Mem1D_10_clock = clock; // @[:@19571.4]
  assign Mem1D_10_reset = reset; // @[:@19572.4]
  assign Mem1D_10_io_r_ofs_0 = _T_2187[8:0]; // @[MemPrimitives.scala 131:28:@21226.4]
  assign Mem1D_10_io_r_backpressure = _T_2187[9]; // @[MemPrimitives.scala 132:32:@21227.4]
  assign Mem1D_10_io_w_ofs_0 = _T_915[8:0]; // @[MemPrimitives.scala 94:28:@20000.4]
  assign Mem1D_10_io_w_data_0 = _T_915[40:9]; // @[MemPrimitives.scala 95:29:@20001.4]
  assign Mem1D_10_io_w_en_0 = _T_915[41]; // @[MemPrimitives.scala 96:27:@20002.4]
  assign Mem1D_11_clock = clock; // @[:@19587.4]
  assign Mem1D_11_reset = reset; // @[:@19588.4]
  assign Mem1D_11_io_r_ofs_0 = _T_2279[8:0]; // @[MemPrimitives.scala 131:28:@21315.4]
  assign Mem1D_11_io_r_backpressure = _T_2279[9]; // @[MemPrimitives.scala 132:32:@21316.4]
  assign Mem1D_11_io_w_ofs_0 = _T_935[8:0]; // @[MemPrimitives.scala 94:28:@20019.4]
  assign Mem1D_11_io_w_data_0 = _T_935[40:9]; // @[MemPrimitives.scala 95:29:@20020.4]
  assign Mem1D_11_io_w_en_0 = _T_935[41]; // @[MemPrimitives.scala 96:27:@20021.4]
  assign Mem1D_12_clock = clock; // @[:@19603.4]
  assign Mem1D_12_reset = reset; // @[:@19604.4]
  assign Mem1D_12_io_r_ofs_0 = _T_2371[8:0]; // @[MemPrimitives.scala 131:28:@21404.4]
  assign Mem1D_12_io_r_backpressure = _T_2371[9]; // @[MemPrimitives.scala 132:32:@21405.4]
  assign Mem1D_12_io_w_ofs_0 = _T_955[8:0]; // @[MemPrimitives.scala 94:28:@20038.4]
  assign Mem1D_12_io_w_data_0 = _T_955[40:9]; // @[MemPrimitives.scala 95:29:@20039.4]
  assign Mem1D_12_io_w_en_0 = _T_955[41]; // @[MemPrimitives.scala 96:27:@20040.4]
  assign Mem1D_13_clock = clock; // @[:@19619.4]
  assign Mem1D_13_reset = reset; // @[:@19620.4]
  assign Mem1D_13_io_r_ofs_0 = _T_2463[8:0]; // @[MemPrimitives.scala 131:28:@21493.4]
  assign Mem1D_13_io_r_backpressure = _T_2463[9]; // @[MemPrimitives.scala 132:32:@21494.4]
  assign Mem1D_13_io_w_ofs_0 = _T_975[8:0]; // @[MemPrimitives.scala 94:28:@20057.4]
  assign Mem1D_13_io_w_data_0 = _T_975[40:9]; // @[MemPrimitives.scala 95:29:@20058.4]
  assign Mem1D_13_io_w_en_0 = _T_975[41]; // @[MemPrimitives.scala 96:27:@20059.4]
  assign Mem1D_14_clock = clock; // @[:@19635.4]
  assign Mem1D_14_reset = reset; // @[:@19636.4]
  assign Mem1D_14_io_r_ofs_0 = _T_2555[8:0]; // @[MemPrimitives.scala 131:28:@21582.4]
  assign Mem1D_14_io_r_backpressure = _T_2555[9]; // @[MemPrimitives.scala 132:32:@21583.4]
  assign Mem1D_14_io_w_ofs_0 = _T_995[8:0]; // @[MemPrimitives.scala 94:28:@20076.4]
  assign Mem1D_14_io_w_data_0 = _T_995[40:9]; // @[MemPrimitives.scala 95:29:@20077.4]
  assign Mem1D_14_io_w_en_0 = _T_995[41]; // @[MemPrimitives.scala 96:27:@20078.4]
  assign Mem1D_15_clock = clock; // @[:@19651.4]
  assign Mem1D_15_reset = reset; // @[:@19652.4]
  assign Mem1D_15_io_r_ofs_0 = _T_2647[8:0]; // @[MemPrimitives.scala 131:28:@21671.4]
  assign Mem1D_15_io_r_backpressure = _T_2647[9]; // @[MemPrimitives.scala 132:32:@21672.4]
  assign Mem1D_15_io_w_ofs_0 = _T_1015[8:0]; // @[MemPrimitives.scala 94:28:@20095.4]
  assign Mem1D_15_io_w_data_0 = _T_1015[40:9]; // @[MemPrimitives.scala 95:29:@20096.4]
  assign Mem1D_15_io_w_en_0 = _T_1015[41]; // @[MemPrimitives.scala 96:27:@20097.4]
  assign Mem1D_16_clock = clock; // @[:@19667.4]
  assign Mem1D_16_reset = reset; // @[:@19668.4]
  assign Mem1D_16_io_r_ofs_0 = _T_2739[8:0]; // @[MemPrimitives.scala 131:28:@21760.4]
  assign Mem1D_16_io_r_backpressure = _T_2739[9]; // @[MemPrimitives.scala 132:32:@21761.4]
  assign Mem1D_16_io_w_ofs_0 = _T_1035[8:0]; // @[MemPrimitives.scala 94:28:@20114.4]
  assign Mem1D_16_io_w_data_0 = _T_1035[40:9]; // @[MemPrimitives.scala 95:29:@20115.4]
  assign Mem1D_16_io_w_en_0 = _T_1035[41]; // @[MemPrimitives.scala 96:27:@20116.4]
  assign Mem1D_17_clock = clock; // @[:@19683.4]
  assign Mem1D_17_reset = reset; // @[:@19684.4]
  assign Mem1D_17_io_r_ofs_0 = _T_2831[8:0]; // @[MemPrimitives.scala 131:28:@21849.4]
  assign Mem1D_17_io_r_backpressure = _T_2831[9]; // @[MemPrimitives.scala 132:32:@21850.4]
  assign Mem1D_17_io_w_ofs_0 = _T_1055[8:0]; // @[MemPrimitives.scala 94:28:@20133.4]
  assign Mem1D_17_io_w_data_0 = _T_1055[40:9]; // @[MemPrimitives.scala 95:29:@20134.4]
  assign Mem1D_17_io_w_en_0 = _T_1055[41]; // @[MemPrimitives.scala 96:27:@20135.4]
  assign Mem1D_18_clock = clock; // @[:@19699.4]
  assign Mem1D_18_reset = reset; // @[:@19700.4]
  assign Mem1D_18_io_r_ofs_0 = _T_2923[8:0]; // @[MemPrimitives.scala 131:28:@21938.4]
  assign Mem1D_18_io_r_backpressure = _T_2923[9]; // @[MemPrimitives.scala 132:32:@21939.4]
  assign Mem1D_18_io_w_ofs_0 = _T_1075[8:0]; // @[MemPrimitives.scala 94:28:@20152.4]
  assign Mem1D_18_io_w_data_0 = _T_1075[40:9]; // @[MemPrimitives.scala 95:29:@20153.4]
  assign Mem1D_18_io_w_en_0 = _T_1075[41]; // @[MemPrimitives.scala 96:27:@20154.4]
  assign Mem1D_19_clock = clock; // @[:@19715.4]
  assign Mem1D_19_reset = reset; // @[:@19716.4]
  assign Mem1D_19_io_r_ofs_0 = _T_3015[8:0]; // @[MemPrimitives.scala 131:28:@22027.4]
  assign Mem1D_19_io_r_backpressure = _T_3015[9]; // @[MemPrimitives.scala 132:32:@22028.4]
  assign Mem1D_19_io_w_ofs_0 = _T_1095[8:0]; // @[MemPrimitives.scala 94:28:@20171.4]
  assign Mem1D_19_io_w_data_0 = _T_1095[40:9]; // @[MemPrimitives.scala 95:29:@20172.4]
  assign Mem1D_19_io_w_en_0 = _T_1095[41]; // @[MemPrimitives.scala 96:27:@20173.4]
  assign Mem1D_20_clock = clock; // @[:@19731.4]
  assign Mem1D_20_reset = reset; // @[:@19732.4]
  assign Mem1D_20_io_r_ofs_0 = _T_3107[8:0]; // @[MemPrimitives.scala 131:28:@22116.4]
  assign Mem1D_20_io_r_backpressure = _T_3107[9]; // @[MemPrimitives.scala 132:32:@22117.4]
  assign Mem1D_20_io_w_ofs_0 = _T_1115[8:0]; // @[MemPrimitives.scala 94:28:@20190.4]
  assign Mem1D_20_io_w_data_0 = _T_1115[40:9]; // @[MemPrimitives.scala 95:29:@20191.4]
  assign Mem1D_20_io_w_en_0 = _T_1115[41]; // @[MemPrimitives.scala 96:27:@20192.4]
  assign Mem1D_21_clock = clock; // @[:@19747.4]
  assign Mem1D_21_reset = reset; // @[:@19748.4]
  assign Mem1D_21_io_r_ofs_0 = _T_3199[8:0]; // @[MemPrimitives.scala 131:28:@22205.4]
  assign Mem1D_21_io_r_backpressure = _T_3199[9]; // @[MemPrimitives.scala 132:32:@22206.4]
  assign Mem1D_21_io_w_ofs_0 = _T_1135[8:0]; // @[MemPrimitives.scala 94:28:@20209.4]
  assign Mem1D_21_io_w_data_0 = _T_1135[40:9]; // @[MemPrimitives.scala 95:29:@20210.4]
  assign Mem1D_21_io_w_en_0 = _T_1135[41]; // @[MemPrimitives.scala 96:27:@20211.4]
  assign Mem1D_22_clock = clock; // @[:@19763.4]
  assign Mem1D_22_reset = reset; // @[:@19764.4]
  assign Mem1D_22_io_r_ofs_0 = _T_3291[8:0]; // @[MemPrimitives.scala 131:28:@22294.4]
  assign Mem1D_22_io_r_backpressure = _T_3291[9]; // @[MemPrimitives.scala 132:32:@22295.4]
  assign Mem1D_22_io_w_ofs_0 = _T_1155[8:0]; // @[MemPrimitives.scala 94:28:@20228.4]
  assign Mem1D_22_io_w_data_0 = _T_1155[40:9]; // @[MemPrimitives.scala 95:29:@20229.4]
  assign Mem1D_22_io_w_en_0 = _T_1155[41]; // @[MemPrimitives.scala 96:27:@20230.4]
  assign Mem1D_23_clock = clock; // @[:@19779.4]
  assign Mem1D_23_reset = reset; // @[:@19780.4]
  assign Mem1D_23_io_r_ofs_0 = _T_3383[8:0]; // @[MemPrimitives.scala 131:28:@22383.4]
  assign Mem1D_23_io_r_backpressure = _T_3383[9]; // @[MemPrimitives.scala 132:32:@22384.4]
  assign Mem1D_23_io_w_ofs_0 = _T_1175[8:0]; // @[MemPrimitives.scala 94:28:@20247.4]
  assign Mem1D_23_io_w_data_0 = _T_1175[40:9]; // @[MemPrimitives.scala 95:29:@20248.4]
  assign Mem1D_23_io_w_en_0 = _T_1175[41]; // @[MemPrimitives.scala 96:27:@20249.4]
  assign StickySelects_clock = clock; // @[:@20287.4]
  assign StickySelects_reset = reset; // @[:@20288.4]
  assign StickySelects_io_ins_0 = io_rPort_1_en_0 & _T_1183; // @[MemPrimitives.scala 125:64:@20289.4]
  assign StickySelects_io_ins_1 = io_rPort_4_en_0 & _T_1189; // @[MemPrimitives.scala 125:64:@20290.4]
  assign StickySelects_io_ins_2 = io_rPort_5_en_0 & _T_1195; // @[MemPrimitives.scala 125:64:@20291.4]
  assign StickySelects_io_ins_3 = io_rPort_7_en_0 & _T_1201; // @[MemPrimitives.scala 125:64:@20292.4]
  assign StickySelects_io_ins_4 = io_rPort_8_en_0 & _T_1207; // @[MemPrimitives.scala 125:64:@20293.4]
  assign StickySelects_io_ins_5 = io_rPort_10_en_0 & _T_1213; // @[MemPrimitives.scala 125:64:@20294.4]
  assign StickySelects_io_ins_6 = io_rPort_11_en_0 & _T_1219; // @[MemPrimitives.scala 125:64:@20295.4]
  assign StickySelects_io_ins_7 = io_rPort_13_en_0 & _T_1225; // @[MemPrimitives.scala 125:64:@20296.4]
  assign StickySelects_io_ins_8 = io_rPort_16_en_0 & _T_1231; // @[MemPrimitives.scala 125:64:@20297.4]
  assign StickySelects_1_clock = clock; // @[:@20376.4]
  assign StickySelects_1_reset = reset; // @[:@20377.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_1275; // @[MemPrimitives.scala 125:64:@20378.4]
  assign StickySelects_1_io_ins_1 = io_rPort_2_en_0 & _T_1281; // @[MemPrimitives.scala 125:64:@20379.4]
  assign StickySelects_1_io_ins_2 = io_rPort_3_en_0 & _T_1287; // @[MemPrimitives.scala 125:64:@20380.4]
  assign StickySelects_1_io_ins_3 = io_rPort_6_en_0 & _T_1293; // @[MemPrimitives.scala 125:64:@20381.4]
  assign StickySelects_1_io_ins_4 = io_rPort_9_en_0 & _T_1299; // @[MemPrimitives.scala 125:64:@20382.4]
  assign StickySelects_1_io_ins_5 = io_rPort_12_en_0 & _T_1305; // @[MemPrimitives.scala 125:64:@20383.4]
  assign StickySelects_1_io_ins_6 = io_rPort_14_en_0 & _T_1311; // @[MemPrimitives.scala 125:64:@20384.4]
  assign StickySelects_1_io_ins_7 = io_rPort_15_en_0 & _T_1317; // @[MemPrimitives.scala 125:64:@20385.4]
  assign StickySelects_1_io_ins_8 = io_rPort_17_en_0 & _T_1323; // @[MemPrimitives.scala 125:64:@20386.4]
  assign StickySelects_2_clock = clock; // @[:@20465.4]
  assign StickySelects_2_reset = reset; // @[:@20466.4]
  assign StickySelects_2_io_ins_0 = io_rPort_1_en_0 & _T_1367; // @[MemPrimitives.scala 125:64:@20467.4]
  assign StickySelects_2_io_ins_1 = io_rPort_4_en_0 & _T_1373; // @[MemPrimitives.scala 125:64:@20468.4]
  assign StickySelects_2_io_ins_2 = io_rPort_5_en_0 & _T_1379; // @[MemPrimitives.scala 125:64:@20469.4]
  assign StickySelects_2_io_ins_3 = io_rPort_7_en_0 & _T_1385; // @[MemPrimitives.scala 125:64:@20470.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_1391; // @[MemPrimitives.scala 125:64:@20471.4]
  assign StickySelects_2_io_ins_5 = io_rPort_10_en_0 & _T_1397; // @[MemPrimitives.scala 125:64:@20472.4]
  assign StickySelects_2_io_ins_6 = io_rPort_11_en_0 & _T_1403; // @[MemPrimitives.scala 125:64:@20473.4]
  assign StickySelects_2_io_ins_7 = io_rPort_13_en_0 & _T_1409; // @[MemPrimitives.scala 125:64:@20474.4]
  assign StickySelects_2_io_ins_8 = io_rPort_16_en_0 & _T_1415; // @[MemPrimitives.scala 125:64:@20475.4]
  assign StickySelects_3_clock = clock; // @[:@20554.4]
  assign StickySelects_3_reset = reset; // @[:@20555.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_1459; // @[MemPrimitives.scala 125:64:@20556.4]
  assign StickySelects_3_io_ins_1 = io_rPort_2_en_0 & _T_1465; // @[MemPrimitives.scala 125:64:@20557.4]
  assign StickySelects_3_io_ins_2 = io_rPort_3_en_0 & _T_1471; // @[MemPrimitives.scala 125:64:@20558.4]
  assign StickySelects_3_io_ins_3 = io_rPort_6_en_0 & _T_1477; // @[MemPrimitives.scala 125:64:@20559.4]
  assign StickySelects_3_io_ins_4 = io_rPort_9_en_0 & _T_1483; // @[MemPrimitives.scala 125:64:@20560.4]
  assign StickySelects_3_io_ins_5 = io_rPort_12_en_0 & _T_1489; // @[MemPrimitives.scala 125:64:@20561.4]
  assign StickySelects_3_io_ins_6 = io_rPort_14_en_0 & _T_1495; // @[MemPrimitives.scala 125:64:@20562.4]
  assign StickySelects_3_io_ins_7 = io_rPort_15_en_0 & _T_1501; // @[MemPrimitives.scala 125:64:@20563.4]
  assign StickySelects_3_io_ins_8 = io_rPort_17_en_0 & _T_1507; // @[MemPrimitives.scala 125:64:@20564.4]
  assign StickySelects_4_clock = clock; // @[:@20643.4]
  assign StickySelects_4_reset = reset; // @[:@20644.4]
  assign StickySelects_4_io_ins_0 = io_rPort_1_en_0 & _T_1551; // @[MemPrimitives.scala 125:64:@20645.4]
  assign StickySelects_4_io_ins_1 = io_rPort_4_en_0 & _T_1557; // @[MemPrimitives.scala 125:64:@20646.4]
  assign StickySelects_4_io_ins_2 = io_rPort_5_en_0 & _T_1563; // @[MemPrimitives.scala 125:64:@20647.4]
  assign StickySelects_4_io_ins_3 = io_rPort_7_en_0 & _T_1569; // @[MemPrimitives.scala 125:64:@20648.4]
  assign StickySelects_4_io_ins_4 = io_rPort_8_en_0 & _T_1575; // @[MemPrimitives.scala 125:64:@20649.4]
  assign StickySelects_4_io_ins_5 = io_rPort_10_en_0 & _T_1581; // @[MemPrimitives.scala 125:64:@20650.4]
  assign StickySelects_4_io_ins_6 = io_rPort_11_en_0 & _T_1587; // @[MemPrimitives.scala 125:64:@20651.4]
  assign StickySelects_4_io_ins_7 = io_rPort_13_en_0 & _T_1593; // @[MemPrimitives.scala 125:64:@20652.4]
  assign StickySelects_4_io_ins_8 = io_rPort_16_en_0 & _T_1599; // @[MemPrimitives.scala 125:64:@20653.4]
  assign StickySelects_5_clock = clock; // @[:@20732.4]
  assign StickySelects_5_reset = reset; // @[:@20733.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_1643; // @[MemPrimitives.scala 125:64:@20734.4]
  assign StickySelects_5_io_ins_1 = io_rPort_2_en_0 & _T_1649; // @[MemPrimitives.scala 125:64:@20735.4]
  assign StickySelects_5_io_ins_2 = io_rPort_3_en_0 & _T_1655; // @[MemPrimitives.scala 125:64:@20736.4]
  assign StickySelects_5_io_ins_3 = io_rPort_6_en_0 & _T_1661; // @[MemPrimitives.scala 125:64:@20737.4]
  assign StickySelects_5_io_ins_4 = io_rPort_9_en_0 & _T_1667; // @[MemPrimitives.scala 125:64:@20738.4]
  assign StickySelects_5_io_ins_5 = io_rPort_12_en_0 & _T_1673; // @[MemPrimitives.scala 125:64:@20739.4]
  assign StickySelects_5_io_ins_6 = io_rPort_14_en_0 & _T_1679; // @[MemPrimitives.scala 125:64:@20740.4]
  assign StickySelects_5_io_ins_7 = io_rPort_15_en_0 & _T_1685; // @[MemPrimitives.scala 125:64:@20741.4]
  assign StickySelects_5_io_ins_8 = io_rPort_17_en_0 & _T_1691; // @[MemPrimitives.scala 125:64:@20742.4]
  assign StickySelects_6_clock = clock; // @[:@20821.4]
  assign StickySelects_6_reset = reset; // @[:@20822.4]
  assign StickySelects_6_io_ins_0 = io_rPort_1_en_0 & _T_1735; // @[MemPrimitives.scala 125:64:@20823.4]
  assign StickySelects_6_io_ins_1 = io_rPort_4_en_0 & _T_1741; // @[MemPrimitives.scala 125:64:@20824.4]
  assign StickySelects_6_io_ins_2 = io_rPort_5_en_0 & _T_1747; // @[MemPrimitives.scala 125:64:@20825.4]
  assign StickySelects_6_io_ins_3 = io_rPort_7_en_0 & _T_1753; // @[MemPrimitives.scala 125:64:@20826.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1759; // @[MemPrimitives.scala 125:64:@20827.4]
  assign StickySelects_6_io_ins_5 = io_rPort_10_en_0 & _T_1765; // @[MemPrimitives.scala 125:64:@20828.4]
  assign StickySelects_6_io_ins_6 = io_rPort_11_en_0 & _T_1771; // @[MemPrimitives.scala 125:64:@20829.4]
  assign StickySelects_6_io_ins_7 = io_rPort_13_en_0 & _T_1777; // @[MemPrimitives.scala 125:64:@20830.4]
  assign StickySelects_6_io_ins_8 = io_rPort_16_en_0 & _T_1783; // @[MemPrimitives.scala 125:64:@20831.4]
  assign StickySelects_7_clock = clock; // @[:@20910.4]
  assign StickySelects_7_reset = reset; // @[:@20911.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1827; // @[MemPrimitives.scala 125:64:@20912.4]
  assign StickySelects_7_io_ins_1 = io_rPort_2_en_0 & _T_1833; // @[MemPrimitives.scala 125:64:@20913.4]
  assign StickySelects_7_io_ins_2 = io_rPort_3_en_0 & _T_1839; // @[MemPrimitives.scala 125:64:@20914.4]
  assign StickySelects_7_io_ins_3 = io_rPort_6_en_0 & _T_1845; // @[MemPrimitives.scala 125:64:@20915.4]
  assign StickySelects_7_io_ins_4 = io_rPort_9_en_0 & _T_1851; // @[MemPrimitives.scala 125:64:@20916.4]
  assign StickySelects_7_io_ins_5 = io_rPort_12_en_0 & _T_1857; // @[MemPrimitives.scala 125:64:@20917.4]
  assign StickySelects_7_io_ins_6 = io_rPort_14_en_0 & _T_1863; // @[MemPrimitives.scala 125:64:@20918.4]
  assign StickySelects_7_io_ins_7 = io_rPort_15_en_0 & _T_1869; // @[MemPrimitives.scala 125:64:@20919.4]
  assign StickySelects_7_io_ins_8 = io_rPort_17_en_0 & _T_1875; // @[MemPrimitives.scala 125:64:@20920.4]
  assign StickySelects_8_clock = clock; // @[:@20999.4]
  assign StickySelects_8_reset = reset; // @[:@21000.4]
  assign StickySelects_8_io_ins_0 = io_rPort_1_en_0 & _T_1919; // @[MemPrimitives.scala 125:64:@21001.4]
  assign StickySelects_8_io_ins_1 = io_rPort_4_en_0 & _T_1925; // @[MemPrimitives.scala 125:64:@21002.4]
  assign StickySelects_8_io_ins_2 = io_rPort_5_en_0 & _T_1931; // @[MemPrimitives.scala 125:64:@21003.4]
  assign StickySelects_8_io_ins_3 = io_rPort_7_en_0 & _T_1937; // @[MemPrimitives.scala 125:64:@21004.4]
  assign StickySelects_8_io_ins_4 = io_rPort_8_en_0 & _T_1943; // @[MemPrimitives.scala 125:64:@21005.4]
  assign StickySelects_8_io_ins_5 = io_rPort_10_en_0 & _T_1949; // @[MemPrimitives.scala 125:64:@21006.4]
  assign StickySelects_8_io_ins_6 = io_rPort_11_en_0 & _T_1955; // @[MemPrimitives.scala 125:64:@21007.4]
  assign StickySelects_8_io_ins_7 = io_rPort_13_en_0 & _T_1961; // @[MemPrimitives.scala 125:64:@21008.4]
  assign StickySelects_8_io_ins_8 = io_rPort_16_en_0 & _T_1967; // @[MemPrimitives.scala 125:64:@21009.4]
  assign StickySelects_9_clock = clock; // @[:@21088.4]
  assign StickySelects_9_reset = reset; // @[:@21089.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_2011; // @[MemPrimitives.scala 125:64:@21090.4]
  assign StickySelects_9_io_ins_1 = io_rPort_2_en_0 & _T_2017; // @[MemPrimitives.scala 125:64:@21091.4]
  assign StickySelects_9_io_ins_2 = io_rPort_3_en_0 & _T_2023; // @[MemPrimitives.scala 125:64:@21092.4]
  assign StickySelects_9_io_ins_3 = io_rPort_6_en_0 & _T_2029; // @[MemPrimitives.scala 125:64:@21093.4]
  assign StickySelects_9_io_ins_4 = io_rPort_9_en_0 & _T_2035; // @[MemPrimitives.scala 125:64:@21094.4]
  assign StickySelects_9_io_ins_5 = io_rPort_12_en_0 & _T_2041; // @[MemPrimitives.scala 125:64:@21095.4]
  assign StickySelects_9_io_ins_6 = io_rPort_14_en_0 & _T_2047; // @[MemPrimitives.scala 125:64:@21096.4]
  assign StickySelects_9_io_ins_7 = io_rPort_15_en_0 & _T_2053; // @[MemPrimitives.scala 125:64:@21097.4]
  assign StickySelects_9_io_ins_8 = io_rPort_17_en_0 & _T_2059; // @[MemPrimitives.scala 125:64:@21098.4]
  assign StickySelects_10_clock = clock; // @[:@21177.4]
  assign StickySelects_10_reset = reset; // @[:@21178.4]
  assign StickySelects_10_io_ins_0 = io_rPort_1_en_0 & _T_2103; // @[MemPrimitives.scala 125:64:@21179.4]
  assign StickySelects_10_io_ins_1 = io_rPort_4_en_0 & _T_2109; // @[MemPrimitives.scala 125:64:@21180.4]
  assign StickySelects_10_io_ins_2 = io_rPort_5_en_0 & _T_2115; // @[MemPrimitives.scala 125:64:@21181.4]
  assign StickySelects_10_io_ins_3 = io_rPort_7_en_0 & _T_2121; // @[MemPrimitives.scala 125:64:@21182.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_2127; // @[MemPrimitives.scala 125:64:@21183.4]
  assign StickySelects_10_io_ins_5 = io_rPort_10_en_0 & _T_2133; // @[MemPrimitives.scala 125:64:@21184.4]
  assign StickySelects_10_io_ins_6 = io_rPort_11_en_0 & _T_2139; // @[MemPrimitives.scala 125:64:@21185.4]
  assign StickySelects_10_io_ins_7 = io_rPort_13_en_0 & _T_2145; // @[MemPrimitives.scala 125:64:@21186.4]
  assign StickySelects_10_io_ins_8 = io_rPort_16_en_0 & _T_2151; // @[MemPrimitives.scala 125:64:@21187.4]
  assign StickySelects_11_clock = clock; // @[:@21266.4]
  assign StickySelects_11_reset = reset; // @[:@21267.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_2195; // @[MemPrimitives.scala 125:64:@21268.4]
  assign StickySelects_11_io_ins_1 = io_rPort_2_en_0 & _T_2201; // @[MemPrimitives.scala 125:64:@21269.4]
  assign StickySelects_11_io_ins_2 = io_rPort_3_en_0 & _T_2207; // @[MemPrimitives.scala 125:64:@21270.4]
  assign StickySelects_11_io_ins_3 = io_rPort_6_en_0 & _T_2213; // @[MemPrimitives.scala 125:64:@21271.4]
  assign StickySelects_11_io_ins_4 = io_rPort_9_en_0 & _T_2219; // @[MemPrimitives.scala 125:64:@21272.4]
  assign StickySelects_11_io_ins_5 = io_rPort_12_en_0 & _T_2225; // @[MemPrimitives.scala 125:64:@21273.4]
  assign StickySelects_11_io_ins_6 = io_rPort_14_en_0 & _T_2231; // @[MemPrimitives.scala 125:64:@21274.4]
  assign StickySelects_11_io_ins_7 = io_rPort_15_en_0 & _T_2237; // @[MemPrimitives.scala 125:64:@21275.4]
  assign StickySelects_11_io_ins_8 = io_rPort_17_en_0 & _T_2243; // @[MemPrimitives.scala 125:64:@21276.4]
  assign StickySelects_12_clock = clock; // @[:@21355.4]
  assign StickySelects_12_reset = reset; // @[:@21356.4]
  assign StickySelects_12_io_ins_0 = io_rPort_1_en_0 & _T_2287; // @[MemPrimitives.scala 125:64:@21357.4]
  assign StickySelects_12_io_ins_1 = io_rPort_4_en_0 & _T_2293; // @[MemPrimitives.scala 125:64:@21358.4]
  assign StickySelects_12_io_ins_2 = io_rPort_5_en_0 & _T_2299; // @[MemPrimitives.scala 125:64:@21359.4]
  assign StickySelects_12_io_ins_3 = io_rPort_7_en_0 & _T_2305; // @[MemPrimitives.scala 125:64:@21360.4]
  assign StickySelects_12_io_ins_4 = io_rPort_8_en_0 & _T_2311; // @[MemPrimitives.scala 125:64:@21361.4]
  assign StickySelects_12_io_ins_5 = io_rPort_10_en_0 & _T_2317; // @[MemPrimitives.scala 125:64:@21362.4]
  assign StickySelects_12_io_ins_6 = io_rPort_11_en_0 & _T_2323; // @[MemPrimitives.scala 125:64:@21363.4]
  assign StickySelects_12_io_ins_7 = io_rPort_13_en_0 & _T_2329; // @[MemPrimitives.scala 125:64:@21364.4]
  assign StickySelects_12_io_ins_8 = io_rPort_16_en_0 & _T_2335; // @[MemPrimitives.scala 125:64:@21365.4]
  assign StickySelects_13_clock = clock; // @[:@21444.4]
  assign StickySelects_13_reset = reset; // @[:@21445.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_2379; // @[MemPrimitives.scala 125:64:@21446.4]
  assign StickySelects_13_io_ins_1 = io_rPort_2_en_0 & _T_2385; // @[MemPrimitives.scala 125:64:@21447.4]
  assign StickySelects_13_io_ins_2 = io_rPort_3_en_0 & _T_2391; // @[MemPrimitives.scala 125:64:@21448.4]
  assign StickySelects_13_io_ins_3 = io_rPort_6_en_0 & _T_2397; // @[MemPrimitives.scala 125:64:@21449.4]
  assign StickySelects_13_io_ins_4 = io_rPort_9_en_0 & _T_2403; // @[MemPrimitives.scala 125:64:@21450.4]
  assign StickySelects_13_io_ins_5 = io_rPort_12_en_0 & _T_2409; // @[MemPrimitives.scala 125:64:@21451.4]
  assign StickySelects_13_io_ins_6 = io_rPort_14_en_0 & _T_2415; // @[MemPrimitives.scala 125:64:@21452.4]
  assign StickySelects_13_io_ins_7 = io_rPort_15_en_0 & _T_2421; // @[MemPrimitives.scala 125:64:@21453.4]
  assign StickySelects_13_io_ins_8 = io_rPort_17_en_0 & _T_2427; // @[MemPrimitives.scala 125:64:@21454.4]
  assign StickySelects_14_clock = clock; // @[:@21533.4]
  assign StickySelects_14_reset = reset; // @[:@21534.4]
  assign StickySelects_14_io_ins_0 = io_rPort_1_en_0 & _T_2471; // @[MemPrimitives.scala 125:64:@21535.4]
  assign StickySelects_14_io_ins_1 = io_rPort_4_en_0 & _T_2477; // @[MemPrimitives.scala 125:64:@21536.4]
  assign StickySelects_14_io_ins_2 = io_rPort_5_en_0 & _T_2483; // @[MemPrimitives.scala 125:64:@21537.4]
  assign StickySelects_14_io_ins_3 = io_rPort_7_en_0 & _T_2489; // @[MemPrimitives.scala 125:64:@21538.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_2495; // @[MemPrimitives.scala 125:64:@21539.4]
  assign StickySelects_14_io_ins_5 = io_rPort_10_en_0 & _T_2501; // @[MemPrimitives.scala 125:64:@21540.4]
  assign StickySelects_14_io_ins_6 = io_rPort_11_en_0 & _T_2507; // @[MemPrimitives.scala 125:64:@21541.4]
  assign StickySelects_14_io_ins_7 = io_rPort_13_en_0 & _T_2513; // @[MemPrimitives.scala 125:64:@21542.4]
  assign StickySelects_14_io_ins_8 = io_rPort_16_en_0 & _T_2519; // @[MemPrimitives.scala 125:64:@21543.4]
  assign StickySelects_15_clock = clock; // @[:@21622.4]
  assign StickySelects_15_reset = reset; // @[:@21623.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_2563; // @[MemPrimitives.scala 125:64:@21624.4]
  assign StickySelects_15_io_ins_1 = io_rPort_2_en_0 & _T_2569; // @[MemPrimitives.scala 125:64:@21625.4]
  assign StickySelects_15_io_ins_2 = io_rPort_3_en_0 & _T_2575; // @[MemPrimitives.scala 125:64:@21626.4]
  assign StickySelects_15_io_ins_3 = io_rPort_6_en_0 & _T_2581; // @[MemPrimitives.scala 125:64:@21627.4]
  assign StickySelects_15_io_ins_4 = io_rPort_9_en_0 & _T_2587; // @[MemPrimitives.scala 125:64:@21628.4]
  assign StickySelects_15_io_ins_5 = io_rPort_12_en_0 & _T_2593; // @[MemPrimitives.scala 125:64:@21629.4]
  assign StickySelects_15_io_ins_6 = io_rPort_14_en_0 & _T_2599; // @[MemPrimitives.scala 125:64:@21630.4]
  assign StickySelects_15_io_ins_7 = io_rPort_15_en_0 & _T_2605; // @[MemPrimitives.scala 125:64:@21631.4]
  assign StickySelects_15_io_ins_8 = io_rPort_17_en_0 & _T_2611; // @[MemPrimitives.scala 125:64:@21632.4]
  assign StickySelects_16_clock = clock; // @[:@21711.4]
  assign StickySelects_16_reset = reset; // @[:@21712.4]
  assign StickySelects_16_io_ins_0 = io_rPort_1_en_0 & _T_2655; // @[MemPrimitives.scala 125:64:@21713.4]
  assign StickySelects_16_io_ins_1 = io_rPort_4_en_0 & _T_2661; // @[MemPrimitives.scala 125:64:@21714.4]
  assign StickySelects_16_io_ins_2 = io_rPort_5_en_0 & _T_2667; // @[MemPrimitives.scala 125:64:@21715.4]
  assign StickySelects_16_io_ins_3 = io_rPort_7_en_0 & _T_2673; // @[MemPrimitives.scala 125:64:@21716.4]
  assign StickySelects_16_io_ins_4 = io_rPort_8_en_0 & _T_2679; // @[MemPrimitives.scala 125:64:@21717.4]
  assign StickySelects_16_io_ins_5 = io_rPort_10_en_0 & _T_2685; // @[MemPrimitives.scala 125:64:@21718.4]
  assign StickySelects_16_io_ins_6 = io_rPort_11_en_0 & _T_2691; // @[MemPrimitives.scala 125:64:@21719.4]
  assign StickySelects_16_io_ins_7 = io_rPort_13_en_0 & _T_2697; // @[MemPrimitives.scala 125:64:@21720.4]
  assign StickySelects_16_io_ins_8 = io_rPort_16_en_0 & _T_2703; // @[MemPrimitives.scala 125:64:@21721.4]
  assign StickySelects_17_clock = clock; // @[:@21800.4]
  assign StickySelects_17_reset = reset; // @[:@21801.4]
  assign StickySelects_17_io_ins_0 = io_rPort_0_en_0 & _T_2747; // @[MemPrimitives.scala 125:64:@21802.4]
  assign StickySelects_17_io_ins_1 = io_rPort_2_en_0 & _T_2753; // @[MemPrimitives.scala 125:64:@21803.4]
  assign StickySelects_17_io_ins_2 = io_rPort_3_en_0 & _T_2759; // @[MemPrimitives.scala 125:64:@21804.4]
  assign StickySelects_17_io_ins_3 = io_rPort_6_en_0 & _T_2765; // @[MemPrimitives.scala 125:64:@21805.4]
  assign StickySelects_17_io_ins_4 = io_rPort_9_en_0 & _T_2771; // @[MemPrimitives.scala 125:64:@21806.4]
  assign StickySelects_17_io_ins_5 = io_rPort_12_en_0 & _T_2777; // @[MemPrimitives.scala 125:64:@21807.4]
  assign StickySelects_17_io_ins_6 = io_rPort_14_en_0 & _T_2783; // @[MemPrimitives.scala 125:64:@21808.4]
  assign StickySelects_17_io_ins_7 = io_rPort_15_en_0 & _T_2789; // @[MemPrimitives.scala 125:64:@21809.4]
  assign StickySelects_17_io_ins_8 = io_rPort_17_en_0 & _T_2795; // @[MemPrimitives.scala 125:64:@21810.4]
  assign StickySelects_18_clock = clock; // @[:@21889.4]
  assign StickySelects_18_reset = reset; // @[:@21890.4]
  assign StickySelects_18_io_ins_0 = io_rPort_1_en_0 & _T_2839; // @[MemPrimitives.scala 125:64:@21891.4]
  assign StickySelects_18_io_ins_1 = io_rPort_4_en_0 & _T_2845; // @[MemPrimitives.scala 125:64:@21892.4]
  assign StickySelects_18_io_ins_2 = io_rPort_5_en_0 & _T_2851; // @[MemPrimitives.scala 125:64:@21893.4]
  assign StickySelects_18_io_ins_3 = io_rPort_7_en_0 & _T_2857; // @[MemPrimitives.scala 125:64:@21894.4]
  assign StickySelects_18_io_ins_4 = io_rPort_8_en_0 & _T_2863; // @[MemPrimitives.scala 125:64:@21895.4]
  assign StickySelects_18_io_ins_5 = io_rPort_10_en_0 & _T_2869; // @[MemPrimitives.scala 125:64:@21896.4]
  assign StickySelects_18_io_ins_6 = io_rPort_11_en_0 & _T_2875; // @[MemPrimitives.scala 125:64:@21897.4]
  assign StickySelects_18_io_ins_7 = io_rPort_13_en_0 & _T_2881; // @[MemPrimitives.scala 125:64:@21898.4]
  assign StickySelects_18_io_ins_8 = io_rPort_16_en_0 & _T_2887; // @[MemPrimitives.scala 125:64:@21899.4]
  assign StickySelects_19_clock = clock; // @[:@21978.4]
  assign StickySelects_19_reset = reset; // @[:@21979.4]
  assign StickySelects_19_io_ins_0 = io_rPort_0_en_0 & _T_2931; // @[MemPrimitives.scala 125:64:@21980.4]
  assign StickySelects_19_io_ins_1 = io_rPort_2_en_0 & _T_2937; // @[MemPrimitives.scala 125:64:@21981.4]
  assign StickySelects_19_io_ins_2 = io_rPort_3_en_0 & _T_2943; // @[MemPrimitives.scala 125:64:@21982.4]
  assign StickySelects_19_io_ins_3 = io_rPort_6_en_0 & _T_2949; // @[MemPrimitives.scala 125:64:@21983.4]
  assign StickySelects_19_io_ins_4 = io_rPort_9_en_0 & _T_2955; // @[MemPrimitives.scala 125:64:@21984.4]
  assign StickySelects_19_io_ins_5 = io_rPort_12_en_0 & _T_2961; // @[MemPrimitives.scala 125:64:@21985.4]
  assign StickySelects_19_io_ins_6 = io_rPort_14_en_0 & _T_2967; // @[MemPrimitives.scala 125:64:@21986.4]
  assign StickySelects_19_io_ins_7 = io_rPort_15_en_0 & _T_2973; // @[MemPrimitives.scala 125:64:@21987.4]
  assign StickySelects_19_io_ins_8 = io_rPort_17_en_0 & _T_2979; // @[MemPrimitives.scala 125:64:@21988.4]
  assign StickySelects_20_clock = clock; // @[:@22067.4]
  assign StickySelects_20_reset = reset; // @[:@22068.4]
  assign StickySelects_20_io_ins_0 = io_rPort_1_en_0 & _T_3023; // @[MemPrimitives.scala 125:64:@22069.4]
  assign StickySelects_20_io_ins_1 = io_rPort_4_en_0 & _T_3029; // @[MemPrimitives.scala 125:64:@22070.4]
  assign StickySelects_20_io_ins_2 = io_rPort_5_en_0 & _T_3035; // @[MemPrimitives.scala 125:64:@22071.4]
  assign StickySelects_20_io_ins_3 = io_rPort_7_en_0 & _T_3041; // @[MemPrimitives.scala 125:64:@22072.4]
  assign StickySelects_20_io_ins_4 = io_rPort_8_en_0 & _T_3047; // @[MemPrimitives.scala 125:64:@22073.4]
  assign StickySelects_20_io_ins_5 = io_rPort_10_en_0 & _T_3053; // @[MemPrimitives.scala 125:64:@22074.4]
  assign StickySelects_20_io_ins_6 = io_rPort_11_en_0 & _T_3059; // @[MemPrimitives.scala 125:64:@22075.4]
  assign StickySelects_20_io_ins_7 = io_rPort_13_en_0 & _T_3065; // @[MemPrimitives.scala 125:64:@22076.4]
  assign StickySelects_20_io_ins_8 = io_rPort_16_en_0 & _T_3071; // @[MemPrimitives.scala 125:64:@22077.4]
  assign StickySelects_21_clock = clock; // @[:@22156.4]
  assign StickySelects_21_reset = reset; // @[:@22157.4]
  assign StickySelects_21_io_ins_0 = io_rPort_0_en_0 & _T_3115; // @[MemPrimitives.scala 125:64:@22158.4]
  assign StickySelects_21_io_ins_1 = io_rPort_2_en_0 & _T_3121; // @[MemPrimitives.scala 125:64:@22159.4]
  assign StickySelects_21_io_ins_2 = io_rPort_3_en_0 & _T_3127; // @[MemPrimitives.scala 125:64:@22160.4]
  assign StickySelects_21_io_ins_3 = io_rPort_6_en_0 & _T_3133; // @[MemPrimitives.scala 125:64:@22161.4]
  assign StickySelects_21_io_ins_4 = io_rPort_9_en_0 & _T_3139; // @[MemPrimitives.scala 125:64:@22162.4]
  assign StickySelects_21_io_ins_5 = io_rPort_12_en_0 & _T_3145; // @[MemPrimitives.scala 125:64:@22163.4]
  assign StickySelects_21_io_ins_6 = io_rPort_14_en_0 & _T_3151; // @[MemPrimitives.scala 125:64:@22164.4]
  assign StickySelects_21_io_ins_7 = io_rPort_15_en_0 & _T_3157; // @[MemPrimitives.scala 125:64:@22165.4]
  assign StickySelects_21_io_ins_8 = io_rPort_17_en_0 & _T_3163; // @[MemPrimitives.scala 125:64:@22166.4]
  assign StickySelects_22_clock = clock; // @[:@22245.4]
  assign StickySelects_22_reset = reset; // @[:@22246.4]
  assign StickySelects_22_io_ins_0 = io_rPort_1_en_0 & _T_3207; // @[MemPrimitives.scala 125:64:@22247.4]
  assign StickySelects_22_io_ins_1 = io_rPort_4_en_0 & _T_3213; // @[MemPrimitives.scala 125:64:@22248.4]
  assign StickySelects_22_io_ins_2 = io_rPort_5_en_0 & _T_3219; // @[MemPrimitives.scala 125:64:@22249.4]
  assign StickySelects_22_io_ins_3 = io_rPort_7_en_0 & _T_3225; // @[MemPrimitives.scala 125:64:@22250.4]
  assign StickySelects_22_io_ins_4 = io_rPort_8_en_0 & _T_3231; // @[MemPrimitives.scala 125:64:@22251.4]
  assign StickySelects_22_io_ins_5 = io_rPort_10_en_0 & _T_3237; // @[MemPrimitives.scala 125:64:@22252.4]
  assign StickySelects_22_io_ins_6 = io_rPort_11_en_0 & _T_3243; // @[MemPrimitives.scala 125:64:@22253.4]
  assign StickySelects_22_io_ins_7 = io_rPort_13_en_0 & _T_3249; // @[MemPrimitives.scala 125:64:@22254.4]
  assign StickySelects_22_io_ins_8 = io_rPort_16_en_0 & _T_3255; // @[MemPrimitives.scala 125:64:@22255.4]
  assign StickySelects_23_clock = clock; // @[:@22334.4]
  assign StickySelects_23_reset = reset; // @[:@22335.4]
  assign StickySelects_23_io_ins_0 = io_rPort_0_en_0 & _T_3299; // @[MemPrimitives.scala 125:64:@22336.4]
  assign StickySelects_23_io_ins_1 = io_rPort_2_en_0 & _T_3305; // @[MemPrimitives.scala 125:64:@22337.4]
  assign StickySelects_23_io_ins_2 = io_rPort_3_en_0 & _T_3311; // @[MemPrimitives.scala 125:64:@22338.4]
  assign StickySelects_23_io_ins_3 = io_rPort_6_en_0 & _T_3317; // @[MemPrimitives.scala 125:64:@22339.4]
  assign StickySelects_23_io_ins_4 = io_rPort_9_en_0 & _T_3323; // @[MemPrimitives.scala 125:64:@22340.4]
  assign StickySelects_23_io_ins_5 = io_rPort_12_en_0 & _T_3329; // @[MemPrimitives.scala 125:64:@22341.4]
  assign StickySelects_23_io_ins_6 = io_rPort_14_en_0 & _T_3335; // @[MemPrimitives.scala 125:64:@22342.4]
  assign StickySelects_23_io_ins_7 = io_rPort_15_en_0 & _T_3341; // @[MemPrimitives.scala 125:64:@22343.4]
  assign StickySelects_23_io_ins_8 = io_rPort_17_en_0 & _T_3347; // @[MemPrimitives.scala 125:64:@22344.4]
  assign RetimeWrapper_clock = clock; // @[:@22424.4]
  assign RetimeWrapper_reset = reset; // @[:@22425.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22427.4]
  assign RetimeWrapper_io_in = _T_1275 & io_rPort_0_en_0; // @[package.scala 94:16:@22426.4]
  assign RetimeWrapper_1_clock = clock; // @[:@22432.4]
  assign RetimeWrapper_1_reset = reset; // @[:@22433.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22435.4]
  assign RetimeWrapper_1_io_in = _T_1459 & io_rPort_0_en_0; // @[package.scala 94:16:@22434.4]
  assign RetimeWrapper_2_clock = clock; // @[:@22440.4]
  assign RetimeWrapper_2_reset = reset; // @[:@22441.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22443.4]
  assign RetimeWrapper_2_io_in = _T_1643 & io_rPort_0_en_0; // @[package.scala 94:16:@22442.4]
  assign RetimeWrapper_3_clock = clock; // @[:@22448.4]
  assign RetimeWrapper_3_reset = reset; // @[:@22449.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22451.4]
  assign RetimeWrapper_3_io_in = _T_1827 & io_rPort_0_en_0; // @[package.scala 94:16:@22450.4]
  assign RetimeWrapper_4_clock = clock; // @[:@22456.4]
  assign RetimeWrapper_4_reset = reset; // @[:@22457.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22459.4]
  assign RetimeWrapper_4_io_in = _T_2011 & io_rPort_0_en_0; // @[package.scala 94:16:@22458.4]
  assign RetimeWrapper_5_clock = clock; // @[:@22464.4]
  assign RetimeWrapper_5_reset = reset; // @[:@22465.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22467.4]
  assign RetimeWrapper_5_io_in = _T_2195 & io_rPort_0_en_0; // @[package.scala 94:16:@22466.4]
  assign RetimeWrapper_6_clock = clock; // @[:@22472.4]
  assign RetimeWrapper_6_reset = reset; // @[:@22473.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22475.4]
  assign RetimeWrapper_6_io_in = _T_2379 & io_rPort_0_en_0; // @[package.scala 94:16:@22474.4]
  assign RetimeWrapper_7_clock = clock; // @[:@22480.4]
  assign RetimeWrapper_7_reset = reset; // @[:@22481.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22483.4]
  assign RetimeWrapper_7_io_in = _T_2563 & io_rPort_0_en_0; // @[package.scala 94:16:@22482.4]
  assign RetimeWrapper_8_clock = clock; // @[:@22488.4]
  assign RetimeWrapper_8_reset = reset; // @[:@22489.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22491.4]
  assign RetimeWrapper_8_io_in = _T_2747 & io_rPort_0_en_0; // @[package.scala 94:16:@22490.4]
  assign RetimeWrapper_9_clock = clock; // @[:@22496.4]
  assign RetimeWrapper_9_reset = reset; // @[:@22497.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22499.4]
  assign RetimeWrapper_9_io_in = _T_2931 & io_rPort_0_en_0; // @[package.scala 94:16:@22498.4]
  assign RetimeWrapper_10_clock = clock; // @[:@22504.4]
  assign RetimeWrapper_10_reset = reset; // @[:@22505.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22507.4]
  assign RetimeWrapper_10_io_in = _T_3115 & io_rPort_0_en_0; // @[package.scala 94:16:@22506.4]
  assign RetimeWrapper_11_clock = clock; // @[:@22512.4]
  assign RetimeWrapper_11_reset = reset; // @[:@22513.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@22515.4]
  assign RetimeWrapper_11_io_in = _T_3299 & io_rPort_0_en_0; // @[package.scala 94:16:@22514.4]
  assign RetimeWrapper_12_clock = clock; // @[:@22568.4]
  assign RetimeWrapper_12_reset = reset; // @[:@22569.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22571.4]
  assign RetimeWrapper_12_io_in = _T_1183 & io_rPort_1_en_0; // @[package.scala 94:16:@22570.4]
  assign RetimeWrapper_13_clock = clock; // @[:@22576.4]
  assign RetimeWrapper_13_reset = reset; // @[:@22577.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22579.4]
  assign RetimeWrapper_13_io_in = _T_1367 & io_rPort_1_en_0; // @[package.scala 94:16:@22578.4]
  assign RetimeWrapper_14_clock = clock; // @[:@22584.4]
  assign RetimeWrapper_14_reset = reset; // @[:@22585.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22587.4]
  assign RetimeWrapper_14_io_in = _T_1551 & io_rPort_1_en_0; // @[package.scala 94:16:@22586.4]
  assign RetimeWrapper_15_clock = clock; // @[:@22592.4]
  assign RetimeWrapper_15_reset = reset; // @[:@22593.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22595.4]
  assign RetimeWrapper_15_io_in = _T_1735 & io_rPort_1_en_0; // @[package.scala 94:16:@22594.4]
  assign RetimeWrapper_16_clock = clock; // @[:@22600.4]
  assign RetimeWrapper_16_reset = reset; // @[:@22601.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22603.4]
  assign RetimeWrapper_16_io_in = _T_1919 & io_rPort_1_en_0; // @[package.scala 94:16:@22602.4]
  assign RetimeWrapper_17_clock = clock; // @[:@22608.4]
  assign RetimeWrapper_17_reset = reset; // @[:@22609.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22611.4]
  assign RetimeWrapper_17_io_in = _T_2103 & io_rPort_1_en_0; // @[package.scala 94:16:@22610.4]
  assign RetimeWrapper_18_clock = clock; // @[:@22616.4]
  assign RetimeWrapper_18_reset = reset; // @[:@22617.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22619.4]
  assign RetimeWrapper_18_io_in = _T_2287 & io_rPort_1_en_0; // @[package.scala 94:16:@22618.4]
  assign RetimeWrapper_19_clock = clock; // @[:@22624.4]
  assign RetimeWrapper_19_reset = reset; // @[:@22625.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22627.4]
  assign RetimeWrapper_19_io_in = _T_2471 & io_rPort_1_en_0; // @[package.scala 94:16:@22626.4]
  assign RetimeWrapper_20_clock = clock; // @[:@22632.4]
  assign RetimeWrapper_20_reset = reset; // @[:@22633.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22635.4]
  assign RetimeWrapper_20_io_in = _T_2655 & io_rPort_1_en_0; // @[package.scala 94:16:@22634.4]
  assign RetimeWrapper_21_clock = clock; // @[:@22640.4]
  assign RetimeWrapper_21_reset = reset; // @[:@22641.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22643.4]
  assign RetimeWrapper_21_io_in = _T_2839 & io_rPort_1_en_0; // @[package.scala 94:16:@22642.4]
  assign RetimeWrapper_22_clock = clock; // @[:@22648.4]
  assign RetimeWrapper_22_reset = reset; // @[:@22649.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22651.4]
  assign RetimeWrapper_22_io_in = _T_3023 & io_rPort_1_en_0; // @[package.scala 94:16:@22650.4]
  assign RetimeWrapper_23_clock = clock; // @[:@22656.4]
  assign RetimeWrapper_23_reset = reset; // @[:@22657.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@22659.4]
  assign RetimeWrapper_23_io_in = _T_3207 & io_rPort_1_en_0; // @[package.scala 94:16:@22658.4]
  assign RetimeWrapper_24_clock = clock; // @[:@22712.4]
  assign RetimeWrapper_24_reset = reset; // @[:@22713.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22715.4]
  assign RetimeWrapper_24_io_in = _T_1281 & io_rPort_2_en_0; // @[package.scala 94:16:@22714.4]
  assign RetimeWrapper_25_clock = clock; // @[:@22720.4]
  assign RetimeWrapper_25_reset = reset; // @[:@22721.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22723.4]
  assign RetimeWrapper_25_io_in = _T_1465 & io_rPort_2_en_0; // @[package.scala 94:16:@22722.4]
  assign RetimeWrapper_26_clock = clock; // @[:@22728.4]
  assign RetimeWrapper_26_reset = reset; // @[:@22729.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22731.4]
  assign RetimeWrapper_26_io_in = _T_1649 & io_rPort_2_en_0; // @[package.scala 94:16:@22730.4]
  assign RetimeWrapper_27_clock = clock; // @[:@22736.4]
  assign RetimeWrapper_27_reset = reset; // @[:@22737.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22739.4]
  assign RetimeWrapper_27_io_in = _T_1833 & io_rPort_2_en_0; // @[package.scala 94:16:@22738.4]
  assign RetimeWrapper_28_clock = clock; // @[:@22744.4]
  assign RetimeWrapper_28_reset = reset; // @[:@22745.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22747.4]
  assign RetimeWrapper_28_io_in = _T_2017 & io_rPort_2_en_0; // @[package.scala 94:16:@22746.4]
  assign RetimeWrapper_29_clock = clock; // @[:@22752.4]
  assign RetimeWrapper_29_reset = reset; // @[:@22753.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22755.4]
  assign RetimeWrapper_29_io_in = _T_2201 & io_rPort_2_en_0; // @[package.scala 94:16:@22754.4]
  assign RetimeWrapper_30_clock = clock; // @[:@22760.4]
  assign RetimeWrapper_30_reset = reset; // @[:@22761.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22763.4]
  assign RetimeWrapper_30_io_in = _T_2385 & io_rPort_2_en_0; // @[package.scala 94:16:@22762.4]
  assign RetimeWrapper_31_clock = clock; // @[:@22768.4]
  assign RetimeWrapper_31_reset = reset; // @[:@22769.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22771.4]
  assign RetimeWrapper_31_io_in = _T_2569 & io_rPort_2_en_0; // @[package.scala 94:16:@22770.4]
  assign RetimeWrapper_32_clock = clock; // @[:@22776.4]
  assign RetimeWrapper_32_reset = reset; // @[:@22777.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22779.4]
  assign RetimeWrapper_32_io_in = _T_2753 & io_rPort_2_en_0; // @[package.scala 94:16:@22778.4]
  assign RetimeWrapper_33_clock = clock; // @[:@22784.4]
  assign RetimeWrapper_33_reset = reset; // @[:@22785.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22787.4]
  assign RetimeWrapper_33_io_in = _T_2937 & io_rPort_2_en_0; // @[package.scala 94:16:@22786.4]
  assign RetimeWrapper_34_clock = clock; // @[:@22792.4]
  assign RetimeWrapper_34_reset = reset; // @[:@22793.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22795.4]
  assign RetimeWrapper_34_io_in = _T_3121 & io_rPort_2_en_0; // @[package.scala 94:16:@22794.4]
  assign RetimeWrapper_35_clock = clock; // @[:@22800.4]
  assign RetimeWrapper_35_reset = reset; // @[:@22801.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@22803.4]
  assign RetimeWrapper_35_io_in = _T_3305 & io_rPort_2_en_0; // @[package.scala 94:16:@22802.4]
  assign RetimeWrapper_36_clock = clock; // @[:@22856.4]
  assign RetimeWrapper_36_reset = reset; // @[:@22857.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22859.4]
  assign RetimeWrapper_36_io_in = _T_1287 & io_rPort_3_en_0; // @[package.scala 94:16:@22858.4]
  assign RetimeWrapper_37_clock = clock; // @[:@22864.4]
  assign RetimeWrapper_37_reset = reset; // @[:@22865.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22867.4]
  assign RetimeWrapper_37_io_in = _T_1471 & io_rPort_3_en_0; // @[package.scala 94:16:@22866.4]
  assign RetimeWrapper_38_clock = clock; // @[:@22872.4]
  assign RetimeWrapper_38_reset = reset; // @[:@22873.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22875.4]
  assign RetimeWrapper_38_io_in = _T_1655 & io_rPort_3_en_0; // @[package.scala 94:16:@22874.4]
  assign RetimeWrapper_39_clock = clock; // @[:@22880.4]
  assign RetimeWrapper_39_reset = reset; // @[:@22881.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22883.4]
  assign RetimeWrapper_39_io_in = _T_1839 & io_rPort_3_en_0; // @[package.scala 94:16:@22882.4]
  assign RetimeWrapper_40_clock = clock; // @[:@22888.4]
  assign RetimeWrapper_40_reset = reset; // @[:@22889.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22891.4]
  assign RetimeWrapper_40_io_in = _T_2023 & io_rPort_3_en_0; // @[package.scala 94:16:@22890.4]
  assign RetimeWrapper_41_clock = clock; // @[:@22896.4]
  assign RetimeWrapper_41_reset = reset; // @[:@22897.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22899.4]
  assign RetimeWrapper_41_io_in = _T_2207 & io_rPort_3_en_0; // @[package.scala 94:16:@22898.4]
  assign RetimeWrapper_42_clock = clock; // @[:@22904.4]
  assign RetimeWrapper_42_reset = reset; // @[:@22905.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22907.4]
  assign RetimeWrapper_42_io_in = _T_2391 & io_rPort_3_en_0; // @[package.scala 94:16:@22906.4]
  assign RetimeWrapper_43_clock = clock; // @[:@22912.4]
  assign RetimeWrapper_43_reset = reset; // @[:@22913.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22915.4]
  assign RetimeWrapper_43_io_in = _T_2575 & io_rPort_3_en_0; // @[package.scala 94:16:@22914.4]
  assign RetimeWrapper_44_clock = clock; // @[:@22920.4]
  assign RetimeWrapper_44_reset = reset; // @[:@22921.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22923.4]
  assign RetimeWrapper_44_io_in = _T_2759 & io_rPort_3_en_0; // @[package.scala 94:16:@22922.4]
  assign RetimeWrapper_45_clock = clock; // @[:@22928.4]
  assign RetimeWrapper_45_reset = reset; // @[:@22929.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22931.4]
  assign RetimeWrapper_45_io_in = _T_2943 & io_rPort_3_en_0; // @[package.scala 94:16:@22930.4]
  assign RetimeWrapper_46_clock = clock; // @[:@22936.4]
  assign RetimeWrapper_46_reset = reset; // @[:@22937.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22939.4]
  assign RetimeWrapper_46_io_in = _T_3127 & io_rPort_3_en_0; // @[package.scala 94:16:@22938.4]
  assign RetimeWrapper_47_clock = clock; // @[:@22944.4]
  assign RetimeWrapper_47_reset = reset; // @[:@22945.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@22947.4]
  assign RetimeWrapper_47_io_in = _T_3311 & io_rPort_3_en_0; // @[package.scala 94:16:@22946.4]
  assign RetimeWrapper_48_clock = clock; // @[:@23000.4]
  assign RetimeWrapper_48_reset = reset; // @[:@23001.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23003.4]
  assign RetimeWrapper_48_io_in = _T_1189 & io_rPort_4_en_0; // @[package.scala 94:16:@23002.4]
  assign RetimeWrapper_49_clock = clock; // @[:@23008.4]
  assign RetimeWrapper_49_reset = reset; // @[:@23009.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23011.4]
  assign RetimeWrapper_49_io_in = _T_1373 & io_rPort_4_en_0; // @[package.scala 94:16:@23010.4]
  assign RetimeWrapper_50_clock = clock; // @[:@23016.4]
  assign RetimeWrapper_50_reset = reset; // @[:@23017.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23019.4]
  assign RetimeWrapper_50_io_in = _T_1557 & io_rPort_4_en_0; // @[package.scala 94:16:@23018.4]
  assign RetimeWrapper_51_clock = clock; // @[:@23024.4]
  assign RetimeWrapper_51_reset = reset; // @[:@23025.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23027.4]
  assign RetimeWrapper_51_io_in = _T_1741 & io_rPort_4_en_0; // @[package.scala 94:16:@23026.4]
  assign RetimeWrapper_52_clock = clock; // @[:@23032.4]
  assign RetimeWrapper_52_reset = reset; // @[:@23033.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23035.4]
  assign RetimeWrapper_52_io_in = _T_1925 & io_rPort_4_en_0; // @[package.scala 94:16:@23034.4]
  assign RetimeWrapper_53_clock = clock; // @[:@23040.4]
  assign RetimeWrapper_53_reset = reset; // @[:@23041.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23043.4]
  assign RetimeWrapper_53_io_in = _T_2109 & io_rPort_4_en_0; // @[package.scala 94:16:@23042.4]
  assign RetimeWrapper_54_clock = clock; // @[:@23048.4]
  assign RetimeWrapper_54_reset = reset; // @[:@23049.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23051.4]
  assign RetimeWrapper_54_io_in = _T_2293 & io_rPort_4_en_0; // @[package.scala 94:16:@23050.4]
  assign RetimeWrapper_55_clock = clock; // @[:@23056.4]
  assign RetimeWrapper_55_reset = reset; // @[:@23057.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23059.4]
  assign RetimeWrapper_55_io_in = _T_2477 & io_rPort_4_en_0; // @[package.scala 94:16:@23058.4]
  assign RetimeWrapper_56_clock = clock; // @[:@23064.4]
  assign RetimeWrapper_56_reset = reset; // @[:@23065.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23067.4]
  assign RetimeWrapper_56_io_in = _T_2661 & io_rPort_4_en_0; // @[package.scala 94:16:@23066.4]
  assign RetimeWrapper_57_clock = clock; // @[:@23072.4]
  assign RetimeWrapper_57_reset = reset; // @[:@23073.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23075.4]
  assign RetimeWrapper_57_io_in = _T_2845 & io_rPort_4_en_0; // @[package.scala 94:16:@23074.4]
  assign RetimeWrapper_58_clock = clock; // @[:@23080.4]
  assign RetimeWrapper_58_reset = reset; // @[:@23081.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23083.4]
  assign RetimeWrapper_58_io_in = _T_3029 & io_rPort_4_en_0; // @[package.scala 94:16:@23082.4]
  assign RetimeWrapper_59_clock = clock; // @[:@23088.4]
  assign RetimeWrapper_59_reset = reset; // @[:@23089.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@23091.4]
  assign RetimeWrapper_59_io_in = _T_3213 & io_rPort_4_en_0; // @[package.scala 94:16:@23090.4]
  assign RetimeWrapper_60_clock = clock; // @[:@23144.4]
  assign RetimeWrapper_60_reset = reset; // @[:@23145.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23147.4]
  assign RetimeWrapper_60_io_in = _T_1195 & io_rPort_5_en_0; // @[package.scala 94:16:@23146.4]
  assign RetimeWrapper_61_clock = clock; // @[:@23152.4]
  assign RetimeWrapper_61_reset = reset; // @[:@23153.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23155.4]
  assign RetimeWrapper_61_io_in = _T_1379 & io_rPort_5_en_0; // @[package.scala 94:16:@23154.4]
  assign RetimeWrapper_62_clock = clock; // @[:@23160.4]
  assign RetimeWrapper_62_reset = reset; // @[:@23161.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23163.4]
  assign RetimeWrapper_62_io_in = _T_1563 & io_rPort_5_en_0; // @[package.scala 94:16:@23162.4]
  assign RetimeWrapper_63_clock = clock; // @[:@23168.4]
  assign RetimeWrapper_63_reset = reset; // @[:@23169.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23171.4]
  assign RetimeWrapper_63_io_in = _T_1747 & io_rPort_5_en_0; // @[package.scala 94:16:@23170.4]
  assign RetimeWrapper_64_clock = clock; // @[:@23176.4]
  assign RetimeWrapper_64_reset = reset; // @[:@23177.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23179.4]
  assign RetimeWrapper_64_io_in = _T_1931 & io_rPort_5_en_0; // @[package.scala 94:16:@23178.4]
  assign RetimeWrapper_65_clock = clock; // @[:@23184.4]
  assign RetimeWrapper_65_reset = reset; // @[:@23185.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23187.4]
  assign RetimeWrapper_65_io_in = _T_2115 & io_rPort_5_en_0; // @[package.scala 94:16:@23186.4]
  assign RetimeWrapper_66_clock = clock; // @[:@23192.4]
  assign RetimeWrapper_66_reset = reset; // @[:@23193.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23195.4]
  assign RetimeWrapper_66_io_in = _T_2299 & io_rPort_5_en_0; // @[package.scala 94:16:@23194.4]
  assign RetimeWrapper_67_clock = clock; // @[:@23200.4]
  assign RetimeWrapper_67_reset = reset; // @[:@23201.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23203.4]
  assign RetimeWrapper_67_io_in = _T_2483 & io_rPort_5_en_0; // @[package.scala 94:16:@23202.4]
  assign RetimeWrapper_68_clock = clock; // @[:@23208.4]
  assign RetimeWrapper_68_reset = reset; // @[:@23209.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23211.4]
  assign RetimeWrapper_68_io_in = _T_2667 & io_rPort_5_en_0; // @[package.scala 94:16:@23210.4]
  assign RetimeWrapper_69_clock = clock; // @[:@23216.4]
  assign RetimeWrapper_69_reset = reset; // @[:@23217.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23219.4]
  assign RetimeWrapper_69_io_in = _T_2851 & io_rPort_5_en_0; // @[package.scala 94:16:@23218.4]
  assign RetimeWrapper_70_clock = clock; // @[:@23224.4]
  assign RetimeWrapper_70_reset = reset; // @[:@23225.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23227.4]
  assign RetimeWrapper_70_io_in = _T_3035 & io_rPort_5_en_0; // @[package.scala 94:16:@23226.4]
  assign RetimeWrapper_71_clock = clock; // @[:@23232.4]
  assign RetimeWrapper_71_reset = reset; // @[:@23233.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@23235.4]
  assign RetimeWrapper_71_io_in = _T_3219 & io_rPort_5_en_0; // @[package.scala 94:16:@23234.4]
  assign RetimeWrapper_72_clock = clock; // @[:@23288.4]
  assign RetimeWrapper_72_reset = reset; // @[:@23289.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23291.4]
  assign RetimeWrapper_72_io_in = _T_1293 & io_rPort_6_en_0; // @[package.scala 94:16:@23290.4]
  assign RetimeWrapper_73_clock = clock; // @[:@23296.4]
  assign RetimeWrapper_73_reset = reset; // @[:@23297.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23299.4]
  assign RetimeWrapper_73_io_in = _T_1477 & io_rPort_6_en_0; // @[package.scala 94:16:@23298.4]
  assign RetimeWrapper_74_clock = clock; // @[:@23304.4]
  assign RetimeWrapper_74_reset = reset; // @[:@23305.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23307.4]
  assign RetimeWrapper_74_io_in = _T_1661 & io_rPort_6_en_0; // @[package.scala 94:16:@23306.4]
  assign RetimeWrapper_75_clock = clock; // @[:@23312.4]
  assign RetimeWrapper_75_reset = reset; // @[:@23313.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23315.4]
  assign RetimeWrapper_75_io_in = _T_1845 & io_rPort_6_en_0; // @[package.scala 94:16:@23314.4]
  assign RetimeWrapper_76_clock = clock; // @[:@23320.4]
  assign RetimeWrapper_76_reset = reset; // @[:@23321.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23323.4]
  assign RetimeWrapper_76_io_in = _T_2029 & io_rPort_6_en_0; // @[package.scala 94:16:@23322.4]
  assign RetimeWrapper_77_clock = clock; // @[:@23328.4]
  assign RetimeWrapper_77_reset = reset; // @[:@23329.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23331.4]
  assign RetimeWrapper_77_io_in = _T_2213 & io_rPort_6_en_0; // @[package.scala 94:16:@23330.4]
  assign RetimeWrapper_78_clock = clock; // @[:@23336.4]
  assign RetimeWrapper_78_reset = reset; // @[:@23337.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23339.4]
  assign RetimeWrapper_78_io_in = _T_2397 & io_rPort_6_en_0; // @[package.scala 94:16:@23338.4]
  assign RetimeWrapper_79_clock = clock; // @[:@23344.4]
  assign RetimeWrapper_79_reset = reset; // @[:@23345.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23347.4]
  assign RetimeWrapper_79_io_in = _T_2581 & io_rPort_6_en_0; // @[package.scala 94:16:@23346.4]
  assign RetimeWrapper_80_clock = clock; // @[:@23352.4]
  assign RetimeWrapper_80_reset = reset; // @[:@23353.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23355.4]
  assign RetimeWrapper_80_io_in = _T_2765 & io_rPort_6_en_0; // @[package.scala 94:16:@23354.4]
  assign RetimeWrapper_81_clock = clock; // @[:@23360.4]
  assign RetimeWrapper_81_reset = reset; // @[:@23361.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23363.4]
  assign RetimeWrapper_81_io_in = _T_2949 & io_rPort_6_en_0; // @[package.scala 94:16:@23362.4]
  assign RetimeWrapper_82_clock = clock; // @[:@23368.4]
  assign RetimeWrapper_82_reset = reset; // @[:@23369.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23371.4]
  assign RetimeWrapper_82_io_in = _T_3133 & io_rPort_6_en_0; // @[package.scala 94:16:@23370.4]
  assign RetimeWrapper_83_clock = clock; // @[:@23376.4]
  assign RetimeWrapper_83_reset = reset; // @[:@23377.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@23379.4]
  assign RetimeWrapper_83_io_in = _T_3317 & io_rPort_6_en_0; // @[package.scala 94:16:@23378.4]
  assign RetimeWrapper_84_clock = clock; // @[:@23432.4]
  assign RetimeWrapper_84_reset = reset; // @[:@23433.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23435.4]
  assign RetimeWrapper_84_io_in = _T_1201 & io_rPort_7_en_0; // @[package.scala 94:16:@23434.4]
  assign RetimeWrapper_85_clock = clock; // @[:@23440.4]
  assign RetimeWrapper_85_reset = reset; // @[:@23441.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23443.4]
  assign RetimeWrapper_85_io_in = _T_1385 & io_rPort_7_en_0; // @[package.scala 94:16:@23442.4]
  assign RetimeWrapper_86_clock = clock; // @[:@23448.4]
  assign RetimeWrapper_86_reset = reset; // @[:@23449.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23451.4]
  assign RetimeWrapper_86_io_in = _T_1569 & io_rPort_7_en_0; // @[package.scala 94:16:@23450.4]
  assign RetimeWrapper_87_clock = clock; // @[:@23456.4]
  assign RetimeWrapper_87_reset = reset; // @[:@23457.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23459.4]
  assign RetimeWrapper_87_io_in = _T_1753 & io_rPort_7_en_0; // @[package.scala 94:16:@23458.4]
  assign RetimeWrapper_88_clock = clock; // @[:@23464.4]
  assign RetimeWrapper_88_reset = reset; // @[:@23465.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23467.4]
  assign RetimeWrapper_88_io_in = _T_1937 & io_rPort_7_en_0; // @[package.scala 94:16:@23466.4]
  assign RetimeWrapper_89_clock = clock; // @[:@23472.4]
  assign RetimeWrapper_89_reset = reset; // @[:@23473.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23475.4]
  assign RetimeWrapper_89_io_in = _T_2121 & io_rPort_7_en_0; // @[package.scala 94:16:@23474.4]
  assign RetimeWrapper_90_clock = clock; // @[:@23480.4]
  assign RetimeWrapper_90_reset = reset; // @[:@23481.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23483.4]
  assign RetimeWrapper_90_io_in = _T_2305 & io_rPort_7_en_0; // @[package.scala 94:16:@23482.4]
  assign RetimeWrapper_91_clock = clock; // @[:@23488.4]
  assign RetimeWrapper_91_reset = reset; // @[:@23489.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23491.4]
  assign RetimeWrapper_91_io_in = _T_2489 & io_rPort_7_en_0; // @[package.scala 94:16:@23490.4]
  assign RetimeWrapper_92_clock = clock; // @[:@23496.4]
  assign RetimeWrapper_92_reset = reset; // @[:@23497.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23499.4]
  assign RetimeWrapper_92_io_in = _T_2673 & io_rPort_7_en_0; // @[package.scala 94:16:@23498.4]
  assign RetimeWrapper_93_clock = clock; // @[:@23504.4]
  assign RetimeWrapper_93_reset = reset; // @[:@23505.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23507.4]
  assign RetimeWrapper_93_io_in = _T_2857 & io_rPort_7_en_0; // @[package.scala 94:16:@23506.4]
  assign RetimeWrapper_94_clock = clock; // @[:@23512.4]
  assign RetimeWrapper_94_reset = reset; // @[:@23513.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23515.4]
  assign RetimeWrapper_94_io_in = _T_3041 & io_rPort_7_en_0; // @[package.scala 94:16:@23514.4]
  assign RetimeWrapper_95_clock = clock; // @[:@23520.4]
  assign RetimeWrapper_95_reset = reset; // @[:@23521.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@23523.4]
  assign RetimeWrapper_95_io_in = _T_3225 & io_rPort_7_en_0; // @[package.scala 94:16:@23522.4]
  assign RetimeWrapper_96_clock = clock; // @[:@23576.4]
  assign RetimeWrapper_96_reset = reset; // @[:@23577.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23579.4]
  assign RetimeWrapper_96_io_in = _T_1207 & io_rPort_8_en_0; // @[package.scala 94:16:@23578.4]
  assign RetimeWrapper_97_clock = clock; // @[:@23584.4]
  assign RetimeWrapper_97_reset = reset; // @[:@23585.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23587.4]
  assign RetimeWrapper_97_io_in = _T_1391 & io_rPort_8_en_0; // @[package.scala 94:16:@23586.4]
  assign RetimeWrapper_98_clock = clock; // @[:@23592.4]
  assign RetimeWrapper_98_reset = reset; // @[:@23593.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23595.4]
  assign RetimeWrapper_98_io_in = _T_1575 & io_rPort_8_en_0; // @[package.scala 94:16:@23594.4]
  assign RetimeWrapper_99_clock = clock; // @[:@23600.4]
  assign RetimeWrapper_99_reset = reset; // @[:@23601.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23603.4]
  assign RetimeWrapper_99_io_in = _T_1759 & io_rPort_8_en_0; // @[package.scala 94:16:@23602.4]
  assign RetimeWrapper_100_clock = clock; // @[:@23608.4]
  assign RetimeWrapper_100_reset = reset; // @[:@23609.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23611.4]
  assign RetimeWrapper_100_io_in = _T_1943 & io_rPort_8_en_0; // @[package.scala 94:16:@23610.4]
  assign RetimeWrapper_101_clock = clock; // @[:@23616.4]
  assign RetimeWrapper_101_reset = reset; // @[:@23617.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23619.4]
  assign RetimeWrapper_101_io_in = _T_2127 & io_rPort_8_en_0; // @[package.scala 94:16:@23618.4]
  assign RetimeWrapper_102_clock = clock; // @[:@23624.4]
  assign RetimeWrapper_102_reset = reset; // @[:@23625.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23627.4]
  assign RetimeWrapper_102_io_in = _T_2311 & io_rPort_8_en_0; // @[package.scala 94:16:@23626.4]
  assign RetimeWrapper_103_clock = clock; // @[:@23632.4]
  assign RetimeWrapper_103_reset = reset; // @[:@23633.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23635.4]
  assign RetimeWrapper_103_io_in = _T_2495 & io_rPort_8_en_0; // @[package.scala 94:16:@23634.4]
  assign RetimeWrapper_104_clock = clock; // @[:@23640.4]
  assign RetimeWrapper_104_reset = reset; // @[:@23641.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23643.4]
  assign RetimeWrapper_104_io_in = _T_2679 & io_rPort_8_en_0; // @[package.scala 94:16:@23642.4]
  assign RetimeWrapper_105_clock = clock; // @[:@23648.4]
  assign RetimeWrapper_105_reset = reset; // @[:@23649.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23651.4]
  assign RetimeWrapper_105_io_in = _T_2863 & io_rPort_8_en_0; // @[package.scala 94:16:@23650.4]
  assign RetimeWrapper_106_clock = clock; // @[:@23656.4]
  assign RetimeWrapper_106_reset = reset; // @[:@23657.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23659.4]
  assign RetimeWrapper_106_io_in = _T_3047 & io_rPort_8_en_0; // @[package.scala 94:16:@23658.4]
  assign RetimeWrapper_107_clock = clock; // @[:@23664.4]
  assign RetimeWrapper_107_reset = reset; // @[:@23665.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@23667.4]
  assign RetimeWrapper_107_io_in = _T_3231 & io_rPort_8_en_0; // @[package.scala 94:16:@23666.4]
  assign RetimeWrapper_108_clock = clock; // @[:@23720.4]
  assign RetimeWrapper_108_reset = reset; // @[:@23721.4]
  assign RetimeWrapper_108_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23723.4]
  assign RetimeWrapper_108_io_in = _T_1299 & io_rPort_9_en_0; // @[package.scala 94:16:@23722.4]
  assign RetimeWrapper_109_clock = clock; // @[:@23728.4]
  assign RetimeWrapper_109_reset = reset; // @[:@23729.4]
  assign RetimeWrapper_109_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23731.4]
  assign RetimeWrapper_109_io_in = _T_1483 & io_rPort_9_en_0; // @[package.scala 94:16:@23730.4]
  assign RetimeWrapper_110_clock = clock; // @[:@23736.4]
  assign RetimeWrapper_110_reset = reset; // @[:@23737.4]
  assign RetimeWrapper_110_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23739.4]
  assign RetimeWrapper_110_io_in = _T_1667 & io_rPort_9_en_0; // @[package.scala 94:16:@23738.4]
  assign RetimeWrapper_111_clock = clock; // @[:@23744.4]
  assign RetimeWrapper_111_reset = reset; // @[:@23745.4]
  assign RetimeWrapper_111_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23747.4]
  assign RetimeWrapper_111_io_in = _T_1851 & io_rPort_9_en_0; // @[package.scala 94:16:@23746.4]
  assign RetimeWrapper_112_clock = clock; // @[:@23752.4]
  assign RetimeWrapper_112_reset = reset; // @[:@23753.4]
  assign RetimeWrapper_112_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23755.4]
  assign RetimeWrapper_112_io_in = _T_2035 & io_rPort_9_en_0; // @[package.scala 94:16:@23754.4]
  assign RetimeWrapper_113_clock = clock; // @[:@23760.4]
  assign RetimeWrapper_113_reset = reset; // @[:@23761.4]
  assign RetimeWrapper_113_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23763.4]
  assign RetimeWrapper_113_io_in = _T_2219 & io_rPort_9_en_0; // @[package.scala 94:16:@23762.4]
  assign RetimeWrapper_114_clock = clock; // @[:@23768.4]
  assign RetimeWrapper_114_reset = reset; // @[:@23769.4]
  assign RetimeWrapper_114_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23771.4]
  assign RetimeWrapper_114_io_in = _T_2403 & io_rPort_9_en_0; // @[package.scala 94:16:@23770.4]
  assign RetimeWrapper_115_clock = clock; // @[:@23776.4]
  assign RetimeWrapper_115_reset = reset; // @[:@23777.4]
  assign RetimeWrapper_115_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23779.4]
  assign RetimeWrapper_115_io_in = _T_2587 & io_rPort_9_en_0; // @[package.scala 94:16:@23778.4]
  assign RetimeWrapper_116_clock = clock; // @[:@23784.4]
  assign RetimeWrapper_116_reset = reset; // @[:@23785.4]
  assign RetimeWrapper_116_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23787.4]
  assign RetimeWrapper_116_io_in = _T_2771 & io_rPort_9_en_0; // @[package.scala 94:16:@23786.4]
  assign RetimeWrapper_117_clock = clock; // @[:@23792.4]
  assign RetimeWrapper_117_reset = reset; // @[:@23793.4]
  assign RetimeWrapper_117_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23795.4]
  assign RetimeWrapper_117_io_in = _T_2955 & io_rPort_9_en_0; // @[package.scala 94:16:@23794.4]
  assign RetimeWrapper_118_clock = clock; // @[:@23800.4]
  assign RetimeWrapper_118_reset = reset; // @[:@23801.4]
  assign RetimeWrapper_118_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23803.4]
  assign RetimeWrapper_118_io_in = _T_3139 & io_rPort_9_en_0; // @[package.scala 94:16:@23802.4]
  assign RetimeWrapper_119_clock = clock; // @[:@23808.4]
  assign RetimeWrapper_119_reset = reset; // @[:@23809.4]
  assign RetimeWrapper_119_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@23811.4]
  assign RetimeWrapper_119_io_in = _T_3323 & io_rPort_9_en_0; // @[package.scala 94:16:@23810.4]
  assign RetimeWrapper_120_clock = clock; // @[:@23864.4]
  assign RetimeWrapper_120_reset = reset; // @[:@23865.4]
  assign RetimeWrapper_120_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23867.4]
  assign RetimeWrapper_120_io_in = _T_1213 & io_rPort_10_en_0; // @[package.scala 94:16:@23866.4]
  assign RetimeWrapper_121_clock = clock; // @[:@23872.4]
  assign RetimeWrapper_121_reset = reset; // @[:@23873.4]
  assign RetimeWrapper_121_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23875.4]
  assign RetimeWrapper_121_io_in = _T_1397 & io_rPort_10_en_0; // @[package.scala 94:16:@23874.4]
  assign RetimeWrapper_122_clock = clock; // @[:@23880.4]
  assign RetimeWrapper_122_reset = reset; // @[:@23881.4]
  assign RetimeWrapper_122_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23883.4]
  assign RetimeWrapper_122_io_in = _T_1581 & io_rPort_10_en_0; // @[package.scala 94:16:@23882.4]
  assign RetimeWrapper_123_clock = clock; // @[:@23888.4]
  assign RetimeWrapper_123_reset = reset; // @[:@23889.4]
  assign RetimeWrapper_123_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23891.4]
  assign RetimeWrapper_123_io_in = _T_1765 & io_rPort_10_en_0; // @[package.scala 94:16:@23890.4]
  assign RetimeWrapper_124_clock = clock; // @[:@23896.4]
  assign RetimeWrapper_124_reset = reset; // @[:@23897.4]
  assign RetimeWrapper_124_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23899.4]
  assign RetimeWrapper_124_io_in = _T_1949 & io_rPort_10_en_0; // @[package.scala 94:16:@23898.4]
  assign RetimeWrapper_125_clock = clock; // @[:@23904.4]
  assign RetimeWrapper_125_reset = reset; // @[:@23905.4]
  assign RetimeWrapper_125_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23907.4]
  assign RetimeWrapper_125_io_in = _T_2133 & io_rPort_10_en_0; // @[package.scala 94:16:@23906.4]
  assign RetimeWrapper_126_clock = clock; // @[:@23912.4]
  assign RetimeWrapper_126_reset = reset; // @[:@23913.4]
  assign RetimeWrapper_126_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23915.4]
  assign RetimeWrapper_126_io_in = _T_2317 & io_rPort_10_en_0; // @[package.scala 94:16:@23914.4]
  assign RetimeWrapper_127_clock = clock; // @[:@23920.4]
  assign RetimeWrapper_127_reset = reset; // @[:@23921.4]
  assign RetimeWrapper_127_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23923.4]
  assign RetimeWrapper_127_io_in = _T_2501 & io_rPort_10_en_0; // @[package.scala 94:16:@23922.4]
  assign RetimeWrapper_128_clock = clock; // @[:@23928.4]
  assign RetimeWrapper_128_reset = reset; // @[:@23929.4]
  assign RetimeWrapper_128_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23931.4]
  assign RetimeWrapper_128_io_in = _T_2685 & io_rPort_10_en_0; // @[package.scala 94:16:@23930.4]
  assign RetimeWrapper_129_clock = clock; // @[:@23936.4]
  assign RetimeWrapper_129_reset = reset; // @[:@23937.4]
  assign RetimeWrapper_129_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23939.4]
  assign RetimeWrapper_129_io_in = _T_2869 & io_rPort_10_en_0; // @[package.scala 94:16:@23938.4]
  assign RetimeWrapper_130_clock = clock; // @[:@23944.4]
  assign RetimeWrapper_130_reset = reset; // @[:@23945.4]
  assign RetimeWrapper_130_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23947.4]
  assign RetimeWrapper_130_io_in = _T_3053 & io_rPort_10_en_0; // @[package.scala 94:16:@23946.4]
  assign RetimeWrapper_131_clock = clock; // @[:@23952.4]
  assign RetimeWrapper_131_reset = reset; // @[:@23953.4]
  assign RetimeWrapper_131_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@23955.4]
  assign RetimeWrapper_131_io_in = _T_3237 & io_rPort_10_en_0; // @[package.scala 94:16:@23954.4]
  assign RetimeWrapper_132_clock = clock; // @[:@24008.4]
  assign RetimeWrapper_132_reset = reset; // @[:@24009.4]
  assign RetimeWrapper_132_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24011.4]
  assign RetimeWrapper_132_io_in = _T_1219 & io_rPort_11_en_0; // @[package.scala 94:16:@24010.4]
  assign RetimeWrapper_133_clock = clock; // @[:@24016.4]
  assign RetimeWrapper_133_reset = reset; // @[:@24017.4]
  assign RetimeWrapper_133_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24019.4]
  assign RetimeWrapper_133_io_in = _T_1403 & io_rPort_11_en_0; // @[package.scala 94:16:@24018.4]
  assign RetimeWrapper_134_clock = clock; // @[:@24024.4]
  assign RetimeWrapper_134_reset = reset; // @[:@24025.4]
  assign RetimeWrapper_134_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24027.4]
  assign RetimeWrapper_134_io_in = _T_1587 & io_rPort_11_en_0; // @[package.scala 94:16:@24026.4]
  assign RetimeWrapper_135_clock = clock; // @[:@24032.4]
  assign RetimeWrapper_135_reset = reset; // @[:@24033.4]
  assign RetimeWrapper_135_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24035.4]
  assign RetimeWrapper_135_io_in = _T_1771 & io_rPort_11_en_0; // @[package.scala 94:16:@24034.4]
  assign RetimeWrapper_136_clock = clock; // @[:@24040.4]
  assign RetimeWrapper_136_reset = reset; // @[:@24041.4]
  assign RetimeWrapper_136_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24043.4]
  assign RetimeWrapper_136_io_in = _T_1955 & io_rPort_11_en_0; // @[package.scala 94:16:@24042.4]
  assign RetimeWrapper_137_clock = clock; // @[:@24048.4]
  assign RetimeWrapper_137_reset = reset; // @[:@24049.4]
  assign RetimeWrapper_137_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24051.4]
  assign RetimeWrapper_137_io_in = _T_2139 & io_rPort_11_en_0; // @[package.scala 94:16:@24050.4]
  assign RetimeWrapper_138_clock = clock; // @[:@24056.4]
  assign RetimeWrapper_138_reset = reset; // @[:@24057.4]
  assign RetimeWrapper_138_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24059.4]
  assign RetimeWrapper_138_io_in = _T_2323 & io_rPort_11_en_0; // @[package.scala 94:16:@24058.4]
  assign RetimeWrapper_139_clock = clock; // @[:@24064.4]
  assign RetimeWrapper_139_reset = reset; // @[:@24065.4]
  assign RetimeWrapper_139_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24067.4]
  assign RetimeWrapper_139_io_in = _T_2507 & io_rPort_11_en_0; // @[package.scala 94:16:@24066.4]
  assign RetimeWrapper_140_clock = clock; // @[:@24072.4]
  assign RetimeWrapper_140_reset = reset; // @[:@24073.4]
  assign RetimeWrapper_140_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24075.4]
  assign RetimeWrapper_140_io_in = _T_2691 & io_rPort_11_en_0; // @[package.scala 94:16:@24074.4]
  assign RetimeWrapper_141_clock = clock; // @[:@24080.4]
  assign RetimeWrapper_141_reset = reset; // @[:@24081.4]
  assign RetimeWrapper_141_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24083.4]
  assign RetimeWrapper_141_io_in = _T_2875 & io_rPort_11_en_0; // @[package.scala 94:16:@24082.4]
  assign RetimeWrapper_142_clock = clock; // @[:@24088.4]
  assign RetimeWrapper_142_reset = reset; // @[:@24089.4]
  assign RetimeWrapper_142_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24091.4]
  assign RetimeWrapper_142_io_in = _T_3059 & io_rPort_11_en_0; // @[package.scala 94:16:@24090.4]
  assign RetimeWrapper_143_clock = clock; // @[:@24096.4]
  assign RetimeWrapper_143_reset = reset; // @[:@24097.4]
  assign RetimeWrapper_143_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@24099.4]
  assign RetimeWrapper_143_io_in = _T_3243 & io_rPort_11_en_0; // @[package.scala 94:16:@24098.4]
  assign RetimeWrapper_144_clock = clock; // @[:@24152.4]
  assign RetimeWrapper_144_reset = reset; // @[:@24153.4]
  assign RetimeWrapper_144_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24155.4]
  assign RetimeWrapper_144_io_in = _T_1305 & io_rPort_12_en_0; // @[package.scala 94:16:@24154.4]
  assign RetimeWrapper_145_clock = clock; // @[:@24160.4]
  assign RetimeWrapper_145_reset = reset; // @[:@24161.4]
  assign RetimeWrapper_145_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24163.4]
  assign RetimeWrapper_145_io_in = _T_1489 & io_rPort_12_en_0; // @[package.scala 94:16:@24162.4]
  assign RetimeWrapper_146_clock = clock; // @[:@24168.4]
  assign RetimeWrapper_146_reset = reset; // @[:@24169.4]
  assign RetimeWrapper_146_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24171.4]
  assign RetimeWrapper_146_io_in = _T_1673 & io_rPort_12_en_0; // @[package.scala 94:16:@24170.4]
  assign RetimeWrapper_147_clock = clock; // @[:@24176.4]
  assign RetimeWrapper_147_reset = reset; // @[:@24177.4]
  assign RetimeWrapper_147_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24179.4]
  assign RetimeWrapper_147_io_in = _T_1857 & io_rPort_12_en_0; // @[package.scala 94:16:@24178.4]
  assign RetimeWrapper_148_clock = clock; // @[:@24184.4]
  assign RetimeWrapper_148_reset = reset; // @[:@24185.4]
  assign RetimeWrapper_148_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24187.4]
  assign RetimeWrapper_148_io_in = _T_2041 & io_rPort_12_en_0; // @[package.scala 94:16:@24186.4]
  assign RetimeWrapper_149_clock = clock; // @[:@24192.4]
  assign RetimeWrapper_149_reset = reset; // @[:@24193.4]
  assign RetimeWrapper_149_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24195.4]
  assign RetimeWrapper_149_io_in = _T_2225 & io_rPort_12_en_0; // @[package.scala 94:16:@24194.4]
  assign RetimeWrapper_150_clock = clock; // @[:@24200.4]
  assign RetimeWrapper_150_reset = reset; // @[:@24201.4]
  assign RetimeWrapper_150_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24203.4]
  assign RetimeWrapper_150_io_in = _T_2409 & io_rPort_12_en_0; // @[package.scala 94:16:@24202.4]
  assign RetimeWrapper_151_clock = clock; // @[:@24208.4]
  assign RetimeWrapper_151_reset = reset; // @[:@24209.4]
  assign RetimeWrapper_151_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24211.4]
  assign RetimeWrapper_151_io_in = _T_2593 & io_rPort_12_en_0; // @[package.scala 94:16:@24210.4]
  assign RetimeWrapper_152_clock = clock; // @[:@24216.4]
  assign RetimeWrapper_152_reset = reset; // @[:@24217.4]
  assign RetimeWrapper_152_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24219.4]
  assign RetimeWrapper_152_io_in = _T_2777 & io_rPort_12_en_0; // @[package.scala 94:16:@24218.4]
  assign RetimeWrapper_153_clock = clock; // @[:@24224.4]
  assign RetimeWrapper_153_reset = reset; // @[:@24225.4]
  assign RetimeWrapper_153_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24227.4]
  assign RetimeWrapper_153_io_in = _T_2961 & io_rPort_12_en_0; // @[package.scala 94:16:@24226.4]
  assign RetimeWrapper_154_clock = clock; // @[:@24232.4]
  assign RetimeWrapper_154_reset = reset; // @[:@24233.4]
  assign RetimeWrapper_154_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24235.4]
  assign RetimeWrapper_154_io_in = _T_3145 & io_rPort_12_en_0; // @[package.scala 94:16:@24234.4]
  assign RetimeWrapper_155_clock = clock; // @[:@24240.4]
  assign RetimeWrapper_155_reset = reset; // @[:@24241.4]
  assign RetimeWrapper_155_io_flow = io_rPort_12_backpressure; // @[package.scala 95:18:@24243.4]
  assign RetimeWrapper_155_io_in = _T_3329 & io_rPort_12_en_0; // @[package.scala 94:16:@24242.4]
  assign RetimeWrapper_156_clock = clock; // @[:@24296.4]
  assign RetimeWrapper_156_reset = reset; // @[:@24297.4]
  assign RetimeWrapper_156_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24299.4]
  assign RetimeWrapper_156_io_in = _T_1225 & io_rPort_13_en_0; // @[package.scala 94:16:@24298.4]
  assign RetimeWrapper_157_clock = clock; // @[:@24304.4]
  assign RetimeWrapper_157_reset = reset; // @[:@24305.4]
  assign RetimeWrapper_157_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24307.4]
  assign RetimeWrapper_157_io_in = _T_1409 & io_rPort_13_en_0; // @[package.scala 94:16:@24306.4]
  assign RetimeWrapper_158_clock = clock; // @[:@24312.4]
  assign RetimeWrapper_158_reset = reset; // @[:@24313.4]
  assign RetimeWrapper_158_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24315.4]
  assign RetimeWrapper_158_io_in = _T_1593 & io_rPort_13_en_0; // @[package.scala 94:16:@24314.4]
  assign RetimeWrapper_159_clock = clock; // @[:@24320.4]
  assign RetimeWrapper_159_reset = reset; // @[:@24321.4]
  assign RetimeWrapper_159_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24323.4]
  assign RetimeWrapper_159_io_in = _T_1777 & io_rPort_13_en_0; // @[package.scala 94:16:@24322.4]
  assign RetimeWrapper_160_clock = clock; // @[:@24328.4]
  assign RetimeWrapper_160_reset = reset; // @[:@24329.4]
  assign RetimeWrapper_160_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24331.4]
  assign RetimeWrapper_160_io_in = _T_1961 & io_rPort_13_en_0; // @[package.scala 94:16:@24330.4]
  assign RetimeWrapper_161_clock = clock; // @[:@24336.4]
  assign RetimeWrapper_161_reset = reset; // @[:@24337.4]
  assign RetimeWrapper_161_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24339.4]
  assign RetimeWrapper_161_io_in = _T_2145 & io_rPort_13_en_0; // @[package.scala 94:16:@24338.4]
  assign RetimeWrapper_162_clock = clock; // @[:@24344.4]
  assign RetimeWrapper_162_reset = reset; // @[:@24345.4]
  assign RetimeWrapper_162_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24347.4]
  assign RetimeWrapper_162_io_in = _T_2329 & io_rPort_13_en_0; // @[package.scala 94:16:@24346.4]
  assign RetimeWrapper_163_clock = clock; // @[:@24352.4]
  assign RetimeWrapper_163_reset = reset; // @[:@24353.4]
  assign RetimeWrapper_163_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24355.4]
  assign RetimeWrapper_163_io_in = _T_2513 & io_rPort_13_en_0; // @[package.scala 94:16:@24354.4]
  assign RetimeWrapper_164_clock = clock; // @[:@24360.4]
  assign RetimeWrapper_164_reset = reset; // @[:@24361.4]
  assign RetimeWrapper_164_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24363.4]
  assign RetimeWrapper_164_io_in = _T_2697 & io_rPort_13_en_0; // @[package.scala 94:16:@24362.4]
  assign RetimeWrapper_165_clock = clock; // @[:@24368.4]
  assign RetimeWrapper_165_reset = reset; // @[:@24369.4]
  assign RetimeWrapper_165_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24371.4]
  assign RetimeWrapper_165_io_in = _T_2881 & io_rPort_13_en_0; // @[package.scala 94:16:@24370.4]
  assign RetimeWrapper_166_clock = clock; // @[:@24376.4]
  assign RetimeWrapper_166_reset = reset; // @[:@24377.4]
  assign RetimeWrapper_166_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24379.4]
  assign RetimeWrapper_166_io_in = _T_3065 & io_rPort_13_en_0; // @[package.scala 94:16:@24378.4]
  assign RetimeWrapper_167_clock = clock; // @[:@24384.4]
  assign RetimeWrapper_167_reset = reset; // @[:@24385.4]
  assign RetimeWrapper_167_io_flow = io_rPort_13_backpressure; // @[package.scala 95:18:@24387.4]
  assign RetimeWrapper_167_io_in = _T_3249 & io_rPort_13_en_0; // @[package.scala 94:16:@24386.4]
  assign RetimeWrapper_168_clock = clock; // @[:@24440.4]
  assign RetimeWrapper_168_reset = reset; // @[:@24441.4]
  assign RetimeWrapper_168_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24443.4]
  assign RetimeWrapper_168_io_in = _T_1311 & io_rPort_14_en_0; // @[package.scala 94:16:@24442.4]
  assign RetimeWrapper_169_clock = clock; // @[:@24448.4]
  assign RetimeWrapper_169_reset = reset; // @[:@24449.4]
  assign RetimeWrapper_169_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24451.4]
  assign RetimeWrapper_169_io_in = _T_1495 & io_rPort_14_en_0; // @[package.scala 94:16:@24450.4]
  assign RetimeWrapper_170_clock = clock; // @[:@24456.4]
  assign RetimeWrapper_170_reset = reset; // @[:@24457.4]
  assign RetimeWrapper_170_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24459.4]
  assign RetimeWrapper_170_io_in = _T_1679 & io_rPort_14_en_0; // @[package.scala 94:16:@24458.4]
  assign RetimeWrapper_171_clock = clock; // @[:@24464.4]
  assign RetimeWrapper_171_reset = reset; // @[:@24465.4]
  assign RetimeWrapper_171_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24467.4]
  assign RetimeWrapper_171_io_in = _T_1863 & io_rPort_14_en_0; // @[package.scala 94:16:@24466.4]
  assign RetimeWrapper_172_clock = clock; // @[:@24472.4]
  assign RetimeWrapper_172_reset = reset; // @[:@24473.4]
  assign RetimeWrapper_172_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24475.4]
  assign RetimeWrapper_172_io_in = _T_2047 & io_rPort_14_en_0; // @[package.scala 94:16:@24474.4]
  assign RetimeWrapper_173_clock = clock; // @[:@24480.4]
  assign RetimeWrapper_173_reset = reset; // @[:@24481.4]
  assign RetimeWrapper_173_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24483.4]
  assign RetimeWrapper_173_io_in = _T_2231 & io_rPort_14_en_0; // @[package.scala 94:16:@24482.4]
  assign RetimeWrapper_174_clock = clock; // @[:@24488.4]
  assign RetimeWrapper_174_reset = reset; // @[:@24489.4]
  assign RetimeWrapper_174_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24491.4]
  assign RetimeWrapper_174_io_in = _T_2415 & io_rPort_14_en_0; // @[package.scala 94:16:@24490.4]
  assign RetimeWrapper_175_clock = clock; // @[:@24496.4]
  assign RetimeWrapper_175_reset = reset; // @[:@24497.4]
  assign RetimeWrapper_175_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24499.4]
  assign RetimeWrapper_175_io_in = _T_2599 & io_rPort_14_en_0; // @[package.scala 94:16:@24498.4]
  assign RetimeWrapper_176_clock = clock; // @[:@24504.4]
  assign RetimeWrapper_176_reset = reset; // @[:@24505.4]
  assign RetimeWrapper_176_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24507.4]
  assign RetimeWrapper_176_io_in = _T_2783 & io_rPort_14_en_0; // @[package.scala 94:16:@24506.4]
  assign RetimeWrapper_177_clock = clock; // @[:@24512.4]
  assign RetimeWrapper_177_reset = reset; // @[:@24513.4]
  assign RetimeWrapper_177_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24515.4]
  assign RetimeWrapper_177_io_in = _T_2967 & io_rPort_14_en_0; // @[package.scala 94:16:@24514.4]
  assign RetimeWrapper_178_clock = clock; // @[:@24520.4]
  assign RetimeWrapper_178_reset = reset; // @[:@24521.4]
  assign RetimeWrapper_178_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24523.4]
  assign RetimeWrapper_178_io_in = _T_3151 & io_rPort_14_en_0; // @[package.scala 94:16:@24522.4]
  assign RetimeWrapper_179_clock = clock; // @[:@24528.4]
  assign RetimeWrapper_179_reset = reset; // @[:@24529.4]
  assign RetimeWrapper_179_io_flow = io_rPort_14_backpressure; // @[package.scala 95:18:@24531.4]
  assign RetimeWrapper_179_io_in = _T_3335 & io_rPort_14_en_0; // @[package.scala 94:16:@24530.4]
  assign RetimeWrapper_180_clock = clock; // @[:@24584.4]
  assign RetimeWrapper_180_reset = reset; // @[:@24585.4]
  assign RetimeWrapper_180_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24587.4]
  assign RetimeWrapper_180_io_in = _T_1317 & io_rPort_15_en_0; // @[package.scala 94:16:@24586.4]
  assign RetimeWrapper_181_clock = clock; // @[:@24592.4]
  assign RetimeWrapper_181_reset = reset; // @[:@24593.4]
  assign RetimeWrapper_181_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24595.4]
  assign RetimeWrapper_181_io_in = _T_1501 & io_rPort_15_en_0; // @[package.scala 94:16:@24594.4]
  assign RetimeWrapper_182_clock = clock; // @[:@24600.4]
  assign RetimeWrapper_182_reset = reset; // @[:@24601.4]
  assign RetimeWrapper_182_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24603.4]
  assign RetimeWrapper_182_io_in = _T_1685 & io_rPort_15_en_0; // @[package.scala 94:16:@24602.4]
  assign RetimeWrapper_183_clock = clock; // @[:@24608.4]
  assign RetimeWrapper_183_reset = reset; // @[:@24609.4]
  assign RetimeWrapper_183_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24611.4]
  assign RetimeWrapper_183_io_in = _T_1869 & io_rPort_15_en_0; // @[package.scala 94:16:@24610.4]
  assign RetimeWrapper_184_clock = clock; // @[:@24616.4]
  assign RetimeWrapper_184_reset = reset; // @[:@24617.4]
  assign RetimeWrapper_184_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24619.4]
  assign RetimeWrapper_184_io_in = _T_2053 & io_rPort_15_en_0; // @[package.scala 94:16:@24618.4]
  assign RetimeWrapper_185_clock = clock; // @[:@24624.4]
  assign RetimeWrapper_185_reset = reset; // @[:@24625.4]
  assign RetimeWrapper_185_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24627.4]
  assign RetimeWrapper_185_io_in = _T_2237 & io_rPort_15_en_0; // @[package.scala 94:16:@24626.4]
  assign RetimeWrapper_186_clock = clock; // @[:@24632.4]
  assign RetimeWrapper_186_reset = reset; // @[:@24633.4]
  assign RetimeWrapper_186_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24635.4]
  assign RetimeWrapper_186_io_in = _T_2421 & io_rPort_15_en_0; // @[package.scala 94:16:@24634.4]
  assign RetimeWrapper_187_clock = clock; // @[:@24640.4]
  assign RetimeWrapper_187_reset = reset; // @[:@24641.4]
  assign RetimeWrapper_187_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24643.4]
  assign RetimeWrapper_187_io_in = _T_2605 & io_rPort_15_en_0; // @[package.scala 94:16:@24642.4]
  assign RetimeWrapper_188_clock = clock; // @[:@24648.4]
  assign RetimeWrapper_188_reset = reset; // @[:@24649.4]
  assign RetimeWrapper_188_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24651.4]
  assign RetimeWrapper_188_io_in = _T_2789 & io_rPort_15_en_0; // @[package.scala 94:16:@24650.4]
  assign RetimeWrapper_189_clock = clock; // @[:@24656.4]
  assign RetimeWrapper_189_reset = reset; // @[:@24657.4]
  assign RetimeWrapper_189_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24659.4]
  assign RetimeWrapper_189_io_in = _T_2973 & io_rPort_15_en_0; // @[package.scala 94:16:@24658.4]
  assign RetimeWrapper_190_clock = clock; // @[:@24664.4]
  assign RetimeWrapper_190_reset = reset; // @[:@24665.4]
  assign RetimeWrapper_190_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24667.4]
  assign RetimeWrapper_190_io_in = _T_3157 & io_rPort_15_en_0; // @[package.scala 94:16:@24666.4]
  assign RetimeWrapper_191_clock = clock; // @[:@24672.4]
  assign RetimeWrapper_191_reset = reset; // @[:@24673.4]
  assign RetimeWrapper_191_io_flow = io_rPort_15_backpressure; // @[package.scala 95:18:@24675.4]
  assign RetimeWrapper_191_io_in = _T_3341 & io_rPort_15_en_0; // @[package.scala 94:16:@24674.4]
  assign RetimeWrapper_192_clock = clock; // @[:@24728.4]
  assign RetimeWrapper_192_reset = reset; // @[:@24729.4]
  assign RetimeWrapper_192_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24731.4]
  assign RetimeWrapper_192_io_in = _T_1231 & io_rPort_16_en_0; // @[package.scala 94:16:@24730.4]
  assign RetimeWrapper_193_clock = clock; // @[:@24736.4]
  assign RetimeWrapper_193_reset = reset; // @[:@24737.4]
  assign RetimeWrapper_193_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24739.4]
  assign RetimeWrapper_193_io_in = _T_1415 & io_rPort_16_en_0; // @[package.scala 94:16:@24738.4]
  assign RetimeWrapper_194_clock = clock; // @[:@24744.4]
  assign RetimeWrapper_194_reset = reset; // @[:@24745.4]
  assign RetimeWrapper_194_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24747.4]
  assign RetimeWrapper_194_io_in = _T_1599 & io_rPort_16_en_0; // @[package.scala 94:16:@24746.4]
  assign RetimeWrapper_195_clock = clock; // @[:@24752.4]
  assign RetimeWrapper_195_reset = reset; // @[:@24753.4]
  assign RetimeWrapper_195_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24755.4]
  assign RetimeWrapper_195_io_in = _T_1783 & io_rPort_16_en_0; // @[package.scala 94:16:@24754.4]
  assign RetimeWrapper_196_clock = clock; // @[:@24760.4]
  assign RetimeWrapper_196_reset = reset; // @[:@24761.4]
  assign RetimeWrapper_196_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24763.4]
  assign RetimeWrapper_196_io_in = _T_1967 & io_rPort_16_en_0; // @[package.scala 94:16:@24762.4]
  assign RetimeWrapper_197_clock = clock; // @[:@24768.4]
  assign RetimeWrapper_197_reset = reset; // @[:@24769.4]
  assign RetimeWrapper_197_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24771.4]
  assign RetimeWrapper_197_io_in = _T_2151 & io_rPort_16_en_0; // @[package.scala 94:16:@24770.4]
  assign RetimeWrapper_198_clock = clock; // @[:@24776.4]
  assign RetimeWrapper_198_reset = reset; // @[:@24777.4]
  assign RetimeWrapper_198_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24779.4]
  assign RetimeWrapper_198_io_in = _T_2335 & io_rPort_16_en_0; // @[package.scala 94:16:@24778.4]
  assign RetimeWrapper_199_clock = clock; // @[:@24784.4]
  assign RetimeWrapper_199_reset = reset; // @[:@24785.4]
  assign RetimeWrapper_199_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24787.4]
  assign RetimeWrapper_199_io_in = _T_2519 & io_rPort_16_en_0; // @[package.scala 94:16:@24786.4]
  assign RetimeWrapper_200_clock = clock; // @[:@24792.4]
  assign RetimeWrapper_200_reset = reset; // @[:@24793.4]
  assign RetimeWrapper_200_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24795.4]
  assign RetimeWrapper_200_io_in = _T_2703 & io_rPort_16_en_0; // @[package.scala 94:16:@24794.4]
  assign RetimeWrapper_201_clock = clock; // @[:@24800.4]
  assign RetimeWrapper_201_reset = reset; // @[:@24801.4]
  assign RetimeWrapper_201_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24803.4]
  assign RetimeWrapper_201_io_in = _T_2887 & io_rPort_16_en_0; // @[package.scala 94:16:@24802.4]
  assign RetimeWrapper_202_clock = clock; // @[:@24808.4]
  assign RetimeWrapper_202_reset = reset; // @[:@24809.4]
  assign RetimeWrapper_202_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24811.4]
  assign RetimeWrapper_202_io_in = _T_3071 & io_rPort_16_en_0; // @[package.scala 94:16:@24810.4]
  assign RetimeWrapper_203_clock = clock; // @[:@24816.4]
  assign RetimeWrapper_203_reset = reset; // @[:@24817.4]
  assign RetimeWrapper_203_io_flow = io_rPort_16_backpressure; // @[package.scala 95:18:@24819.4]
  assign RetimeWrapper_203_io_in = _T_3255 & io_rPort_16_en_0; // @[package.scala 94:16:@24818.4]
  assign RetimeWrapper_204_clock = clock; // @[:@24872.4]
  assign RetimeWrapper_204_reset = reset; // @[:@24873.4]
  assign RetimeWrapper_204_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24875.4]
  assign RetimeWrapper_204_io_in = _T_1323 & io_rPort_17_en_0; // @[package.scala 94:16:@24874.4]
  assign RetimeWrapper_205_clock = clock; // @[:@24880.4]
  assign RetimeWrapper_205_reset = reset; // @[:@24881.4]
  assign RetimeWrapper_205_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24883.4]
  assign RetimeWrapper_205_io_in = _T_1507 & io_rPort_17_en_0; // @[package.scala 94:16:@24882.4]
  assign RetimeWrapper_206_clock = clock; // @[:@24888.4]
  assign RetimeWrapper_206_reset = reset; // @[:@24889.4]
  assign RetimeWrapper_206_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24891.4]
  assign RetimeWrapper_206_io_in = _T_1691 & io_rPort_17_en_0; // @[package.scala 94:16:@24890.4]
  assign RetimeWrapper_207_clock = clock; // @[:@24896.4]
  assign RetimeWrapper_207_reset = reset; // @[:@24897.4]
  assign RetimeWrapper_207_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24899.4]
  assign RetimeWrapper_207_io_in = _T_1875 & io_rPort_17_en_0; // @[package.scala 94:16:@24898.4]
  assign RetimeWrapper_208_clock = clock; // @[:@24904.4]
  assign RetimeWrapper_208_reset = reset; // @[:@24905.4]
  assign RetimeWrapper_208_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24907.4]
  assign RetimeWrapper_208_io_in = _T_2059 & io_rPort_17_en_0; // @[package.scala 94:16:@24906.4]
  assign RetimeWrapper_209_clock = clock; // @[:@24912.4]
  assign RetimeWrapper_209_reset = reset; // @[:@24913.4]
  assign RetimeWrapper_209_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24915.4]
  assign RetimeWrapper_209_io_in = _T_2243 & io_rPort_17_en_0; // @[package.scala 94:16:@24914.4]
  assign RetimeWrapper_210_clock = clock; // @[:@24920.4]
  assign RetimeWrapper_210_reset = reset; // @[:@24921.4]
  assign RetimeWrapper_210_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24923.4]
  assign RetimeWrapper_210_io_in = _T_2427 & io_rPort_17_en_0; // @[package.scala 94:16:@24922.4]
  assign RetimeWrapper_211_clock = clock; // @[:@24928.4]
  assign RetimeWrapper_211_reset = reset; // @[:@24929.4]
  assign RetimeWrapper_211_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24931.4]
  assign RetimeWrapper_211_io_in = _T_2611 & io_rPort_17_en_0; // @[package.scala 94:16:@24930.4]
  assign RetimeWrapper_212_clock = clock; // @[:@24936.4]
  assign RetimeWrapper_212_reset = reset; // @[:@24937.4]
  assign RetimeWrapper_212_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24939.4]
  assign RetimeWrapper_212_io_in = _T_2795 & io_rPort_17_en_0; // @[package.scala 94:16:@24938.4]
  assign RetimeWrapper_213_clock = clock; // @[:@24944.4]
  assign RetimeWrapper_213_reset = reset; // @[:@24945.4]
  assign RetimeWrapper_213_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24947.4]
  assign RetimeWrapper_213_io_in = _T_2979 & io_rPort_17_en_0; // @[package.scala 94:16:@24946.4]
  assign RetimeWrapper_214_clock = clock; // @[:@24952.4]
  assign RetimeWrapper_214_reset = reset; // @[:@24953.4]
  assign RetimeWrapper_214_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24955.4]
  assign RetimeWrapper_214_io_in = _T_3163 & io_rPort_17_en_0; // @[package.scala 94:16:@24954.4]
  assign RetimeWrapper_215_clock = clock; // @[:@24960.4]
  assign RetimeWrapper_215_reset = reset; // @[:@24961.4]
  assign RetimeWrapper_215_io_flow = io_rPort_17_backpressure; // @[package.scala 95:18:@24963.4]
  assign RetimeWrapper_215_io_in = _T_3347 & io_rPort_17_en_0; // @[package.scala 94:16:@24962.4]
endmodule
module StickySelects_25( // @[:@27547.2]
  input   clock, // @[:@27548.4]
  input   reset, // @[:@27549.4]
  input   io_ins_0, // @[:@27550.4]
  input   io_ins_1, // @[:@27550.4]
  input   io_ins_2, // @[:@27550.4]
  input   io_ins_3, // @[:@27550.4]
  output  io_outs_0, // @[:@27550.4]
  output  io_outs_1, // @[:@27550.4]
  output  io_outs_2, // @[:@27550.4]
  output  io_outs_3 // @[:@27550.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@27552.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@27553.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@27554.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@27555.4]
  reg [31:0] _RAND_3;
  wire  _T_29; // @[StickySelects.scala 47:46:@27556.4]
  wire  _T_30; // @[StickySelects.scala 47:46:@27557.4]
  wire  _T_31; // @[StickySelects.scala 49:53:@27558.4]
  wire  _T_32; // @[StickySelects.scala 49:21:@27559.4]
  wire  _T_33; // @[StickySelects.scala 47:46:@27561.4]
  wire  _T_34; // @[StickySelects.scala 47:46:@27562.4]
  wire  _T_35; // @[StickySelects.scala 49:53:@27563.4]
  wire  _T_36; // @[StickySelects.scala 49:21:@27564.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@27566.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@27567.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@27568.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@27569.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@27572.4]
  wire  _T_43; // @[StickySelects.scala 49:53:@27573.4]
  wire  _T_44; // @[StickySelects.scala 49:21:@27574.4]
  assign _T_29 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@27556.4]
  assign _T_30 = _T_29 | io_ins_3; // @[StickySelects.scala 47:46:@27557.4]
  assign _T_31 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@27558.4]
  assign _T_32 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 49:21:@27559.4]
  assign _T_33 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@27561.4]
  assign _T_34 = _T_33 | io_ins_3; // @[StickySelects.scala 47:46:@27562.4]
  assign _T_35 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@27563.4]
  assign _T_36 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 49:21:@27564.4]
  assign _T_37 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@27566.4]
  assign _T_38 = _T_37 | io_ins_3; // @[StickySelects.scala 47:46:@27567.4]
  assign _T_39 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@27568.4]
  assign _T_40 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 49:21:@27569.4]
  assign _T_42 = _T_37 | io_ins_2; // @[StickySelects.scala 47:46:@27572.4]
  assign _T_43 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@27573.4]
  assign _T_44 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 49:21:@27574.4]
  assign io_outs_0 = _T_30 ? io_ins_0 : _T_31; // @[StickySelects.scala 53:57:@27576.4]
  assign io_outs_1 = _T_34 ? io_ins_1 : _T_35; // @[StickySelects.scala 53:57:@27577.4]
  assign io_outs_2 = _T_38 ? io_ins_2 : _T_39; // @[StickySelects.scala 53:57:@27578.4]
  assign io_outs_3 = _T_42 ? io_ins_3 : _T_43; // @[StickySelects.scala 53:57:@27579.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_30) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_31;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_34) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_35;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_39;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_42) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_43;
      end
    end
  end
endmodule
module StickySelects_26( // @[:@27581.2]
  input   clock, // @[:@27582.4]
  input   reset, // @[:@27583.4]
  input   io_ins_0, // @[:@27584.4]
  input   io_ins_1, // @[:@27584.4]
  input   io_ins_2, // @[:@27584.4]
  input   io_ins_3, // @[:@27584.4]
  input   io_ins_4, // @[:@27584.4]
  input   io_ins_5, // @[:@27584.4]
  output  io_outs_0, // @[:@27584.4]
  output  io_outs_1, // @[:@27584.4]
  output  io_outs_2, // @[:@27584.4]
  output  io_outs_3, // @[:@27584.4]
  output  io_outs_4, // @[:@27584.4]
  output  io_outs_5 // @[:@27584.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@27586.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@27587.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@27588.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@27589.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@27590.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@27591.4]
  reg [31:0] _RAND_5;
  wire  _T_35; // @[StickySelects.scala 47:46:@27592.4]
  wire  _T_36; // @[StickySelects.scala 47:46:@27593.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@27594.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@27595.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@27596.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@27597.4]
  wire  _T_41; // @[StickySelects.scala 47:46:@27599.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@27600.4]
  wire  _T_43; // @[StickySelects.scala 47:46:@27601.4]
  wire  _T_44; // @[StickySelects.scala 47:46:@27602.4]
  wire  _T_45; // @[StickySelects.scala 49:53:@27603.4]
  wire  _T_46; // @[StickySelects.scala 49:21:@27604.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@27606.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@27607.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@27608.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@27609.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@27610.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@27611.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@27614.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@27615.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@27616.4]
  wire  _T_57; // @[StickySelects.scala 49:53:@27617.4]
  wire  _T_58; // @[StickySelects.scala 49:21:@27618.4]
  wire  _T_61; // @[StickySelects.scala 47:46:@27622.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@27623.4]
  wire  _T_63; // @[StickySelects.scala 49:53:@27624.4]
  wire  _T_64; // @[StickySelects.scala 49:21:@27625.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@27630.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@27631.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@27632.4]
  assign _T_35 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@27592.4]
  assign _T_36 = _T_35 | io_ins_3; // @[StickySelects.scala 47:46:@27593.4]
  assign _T_37 = _T_36 | io_ins_4; // @[StickySelects.scala 47:46:@27594.4]
  assign _T_38 = _T_37 | io_ins_5; // @[StickySelects.scala 47:46:@27595.4]
  assign _T_39 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@27596.4]
  assign _T_40 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 49:21:@27597.4]
  assign _T_41 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@27599.4]
  assign _T_42 = _T_41 | io_ins_3; // @[StickySelects.scala 47:46:@27600.4]
  assign _T_43 = _T_42 | io_ins_4; // @[StickySelects.scala 47:46:@27601.4]
  assign _T_44 = _T_43 | io_ins_5; // @[StickySelects.scala 47:46:@27602.4]
  assign _T_45 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@27603.4]
  assign _T_46 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 49:21:@27604.4]
  assign _T_47 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@27606.4]
  assign _T_48 = _T_47 | io_ins_3; // @[StickySelects.scala 47:46:@27607.4]
  assign _T_49 = _T_48 | io_ins_4; // @[StickySelects.scala 47:46:@27608.4]
  assign _T_50 = _T_49 | io_ins_5; // @[StickySelects.scala 47:46:@27609.4]
  assign _T_51 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@27610.4]
  assign _T_52 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 49:21:@27611.4]
  assign _T_54 = _T_47 | io_ins_2; // @[StickySelects.scala 47:46:@27614.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@27615.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@27616.4]
  assign _T_57 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@27617.4]
  assign _T_58 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 49:21:@27618.4]
  assign _T_61 = _T_54 | io_ins_3; // @[StickySelects.scala 47:46:@27622.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 47:46:@27623.4]
  assign _T_63 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@27624.4]
  assign _T_64 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 49:21:@27625.4]
  assign _T_68 = _T_61 | io_ins_4; // @[StickySelects.scala 47:46:@27630.4]
  assign _T_69 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@27631.4]
  assign _T_70 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 49:21:@27632.4]
  assign io_outs_0 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 53:57:@27634.4]
  assign io_outs_1 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 53:57:@27635.4]
  assign io_outs_2 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 53:57:@27636.4]
  assign io_outs_3 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 53:57:@27637.4]
  assign io_outs_4 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 53:57:@27638.4]
  assign io_outs_5 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 53:57:@27639.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_39;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_45;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_51;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_56) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_57;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_62) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_63;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_69;
      end
    end
  end
endmodule
module x384_lb2_0( // @[:@32515.2]
  input         clock, // @[:@32516.4]
  input         reset, // @[:@32517.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@32518.4]
  input         io_rPort_9_en_0, // @[:@32518.4]
  input         io_rPort_9_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_9_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@32518.4]
  input         io_rPort_8_en_0, // @[:@32518.4]
  input         io_rPort_8_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_8_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@32518.4]
  input         io_rPort_7_en_0, // @[:@32518.4]
  input         io_rPort_7_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_7_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@32518.4]
  input         io_rPort_6_en_0, // @[:@32518.4]
  input         io_rPort_6_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_6_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@32518.4]
  input         io_rPort_5_en_0, // @[:@32518.4]
  input         io_rPort_5_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_5_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@32518.4]
  input         io_rPort_4_en_0, // @[:@32518.4]
  input         io_rPort_4_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_4_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@32518.4]
  input         io_rPort_3_en_0, // @[:@32518.4]
  input         io_rPort_3_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_3_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@32518.4]
  input         io_rPort_2_en_0, // @[:@32518.4]
  input         io_rPort_2_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_2_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@32518.4]
  input         io_rPort_1_en_0, // @[:@32518.4]
  input         io_rPort_1_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_1_output_0, // @[:@32518.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@32518.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@32518.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@32518.4]
  input         io_rPort_0_en_0, // @[:@32518.4]
  input         io_rPort_0_backpressure, // @[:@32518.4]
  output [31:0] io_rPort_0_output_0, // @[:@32518.4]
  input  [2:0]  io_wPort_3_banks_1, // @[:@32518.4]
  input  [2:0]  io_wPort_3_banks_0, // @[:@32518.4]
  input  [8:0]  io_wPort_3_ofs_0, // @[:@32518.4]
  input  [31:0] io_wPort_3_data_0, // @[:@32518.4]
  input         io_wPort_3_en_0, // @[:@32518.4]
  input  [2:0]  io_wPort_2_banks_1, // @[:@32518.4]
  input  [2:0]  io_wPort_2_banks_0, // @[:@32518.4]
  input  [8:0]  io_wPort_2_ofs_0, // @[:@32518.4]
  input  [31:0] io_wPort_2_data_0, // @[:@32518.4]
  input         io_wPort_2_en_0, // @[:@32518.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@32518.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@32518.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@32518.4]
  input  [31:0] io_wPort_1_data_0, // @[:@32518.4]
  input         io_wPort_1_en_0, // @[:@32518.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@32518.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@32518.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@32518.4]
  input  [31:0] io_wPort_0_data_0, // @[:@32518.4]
  input         io_wPort_0_en_0 // @[:@32518.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@32613.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@32613.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32613.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32613.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32613.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@32613.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@32613.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@32613.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@32629.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@32629.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32629.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32629.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32629.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@32629.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@32629.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@32629.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@32645.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@32645.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32645.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32645.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32645.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@32645.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@32645.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@32645.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@32661.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@32661.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32661.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32661.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32661.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@32661.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@32661.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@32661.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@32677.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@32677.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32677.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32677.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32677.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@32677.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@32677.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@32677.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@32693.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@32693.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32693.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32693.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32693.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@32693.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@32693.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@32693.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@32709.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@32709.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32709.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32709.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32709.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@32709.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@32709.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@32709.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@32725.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@32725.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32725.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32725.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32725.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@32725.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@32725.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@32725.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@32741.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@32741.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32741.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32741.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32741.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@32741.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@32741.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@32741.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@32757.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@32757.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32757.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32757.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32757.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@32757.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@32757.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@32757.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@32773.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@32773.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32773.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32773.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32773.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@32773.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@32773.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@32773.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@32789.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@32789.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32789.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32789.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32789.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@32789.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@32789.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@32789.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@32805.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@32805.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32805.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32805.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32805.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@32805.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@32805.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@32805.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@32821.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@32821.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32821.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32821.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32821.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@32821.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@32821.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@32821.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@32837.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@32837.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32837.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32837.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32837.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@32837.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@32837.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@32837.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@32853.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@32853.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32853.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32853.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32853.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@32853.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@32853.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@32853.4]
  wire  Mem1D_16_clock; // @[MemPrimitives.scala 64:21:@32869.4]
  wire  Mem1D_16_reset; // @[MemPrimitives.scala 64:21:@32869.4]
  wire [8:0] Mem1D_16_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32869.4]
  wire  Mem1D_16_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32869.4]
  wire [8:0] Mem1D_16_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32869.4]
  wire [31:0] Mem1D_16_io_w_data_0; // @[MemPrimitives.scala 64:21:@32869.4]
  wire  Mem1D_16_io_w_en_0; // @[MemPrimitives.scala 64:21:@32869.4]
  wire [31:0] Mem1D_16_io_output; // @[MemPrimitives.scala 64:21:@32869.4]
  wire  Mem1D_17_clock; // @[MemPrimitives.scala 64:21:@32885.4]
  wire  Mem1D_17_reset; // @[MemPrimitives.scala 64:21:@32885.4]
  wire [8:0] Mem1D_17_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32885.4]
  wire  Mem1D_17_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32885.4]
  wire [8:0] Mem1D_17_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32885.4]
  wire [31:0] Mem1D_17_io_w_data_0; // @[MemPrimitives.scala 64:21:@32885.4]
  wire  Mem1D_17_io_w_en_0; // @[MemPrimitives.scala 64:21:@32885.4]
  wire [31:0] Mem1D_17_io_output; // @[MemPrimitives.scala 64:21:@32885.4]
  wire  Mem1D_18_clock; // @[MemPrimitives.scala 64:21:@32901.4]
  wire  Mem1D_18_reset; // @[MemPrimitives.scala 64:21:@32901.4]
  wire [8:0] Mem1D_18_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32901.4]
  wire  Mem1D_18_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32901.4]
  wire [8:0] Mem1D_18_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32901.4]
  wire [31:0] Mem1D_18_io_w_data_0; // @[MemPrimitives.scala 64:21:@32901.4]
  wire  Mem1D_18_io_w_en_0; // @[MemPrimitives.scala 64:21:@32901.4]
  wire [31:0] Mem1D_18_io_output; // @[MemPrimitives.scala 64:21:@32901.4]
  wire  Mem1D_19_clock; // @[MemPrimitives.scala 64:21:@32917.4]
  wire  Mem1D_19_reset; // @[MemPrimitives.scala 64:21:@32917.4]
  wire [8:0] Mem1D_19_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32917.4]
  wire  Mem1D_19_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32917.4]
  wire [8:0] Mem1D_19_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32917.4]
  wire [31:0] Mem1D_19_io_w_data_0; // @[MemPrimitives.scala 64:21:@32917.4]
  wire  Mem1D_19_io_w_en_0; // @[MemPrimitives.scala 64:21:@32917.4]
  wire [31:0] Mem1D_19_io_output; // @[MemPrimitives.scala 64:21:@32917.4]
  wire  Mem1D_20_clock; // @[MemPrimitives.scala 64:21:@32933.4]
  wire  Mem1D_20_reset; // @[MemPrimitives.scala 64:21:@32933.4]
  wire [8:0] Mem1D_20_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32933.4]
  wire  Mem1D_20_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32933.4]
  wire [8:0] Mem1D_20_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32933.4]
  wire [31:0] Mem1D_20_io_w_data_0; // @[MemPrimitives.scala 64:21:@32933.4]
  wire  Mem1D_20_io_w_en_0; // @[MemPrimitives.scala 64:21:@32933.4]
  wire [31:0] Mem1D_20_io_output; // @[MemPrimitives.scala 64:21:@32933.4]
  wire  Mem1D_21_clock; // @[MemPrimitives.scala 64:21:@32949.4]
  wire  Mem1D_21_reset; // @[MemPrimitives.scala 64:21:@32949.4]
  wire [8:0] Mem1D_21_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32949.4]
  wire  Mem1D_21_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32949.4]
  wire [8:0] Mem1D_21_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32949.4]
  wire [31:0] Mem1D_21_io_w_data_0; // @[MemPrimitives.scala 64:21:@32949.4]
  wire  Mem1D_21_io_w_en_0; // @[MemPrimitives.scala 64:21:@32949.4]
  wire [31:0] Mem1D_21_io_output; // @[MemPrimitives.scala 64:21:@32949.4]
  wire  Mem1D_22_clock; // @[MemPrimitives.scala 64:21:@32965.4]
  wire  Mem1D_22_reset; // @[MemPrimitives.scala 64:21:@32965.4]
  wire [8:0] Mem1D_22_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32965.4]
  wire  Mem1D_22_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32965.4]
  wire [8:0] Mem1D_22_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32965.4]
  wire [31:0] Mem1D_22_io_w_data_0; // @[MemPrimitives.scala 64:21:@32965.4]
  wire  Mem1D_22_io_w_en_0; // @[MemPrimitives.scala 64:21:@32965.4]
  wire [31:0] Mem1D_22_io_output; // @[MemPrimitives.scala 64:21:@32965.4]
  wire  Mem1D_23_clock; // @[MemPrimitives.scala 64:21:@32981.4]
  wire  Mem1D_23_reset; // @[MemPrimitives.scala 64:21:@32981.4]
  wire [8:0] Mem1D_23_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@32981.4]
  wire  Mem1D_23_io_r_backpressure; // @[MemPrimitives.scala 64:21:@32981.4]
  wire [8:0] Mem1D_23_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@32981.4]
  wire [31:0] Mem1D_23_io_w_data_0; // @[MemPrimitives.scala 64:21:@32981.4]
  wire  Mem1D_23_io_w_en_0; // @[MemPrimitives.scala 64:21:@32981.4]
  wire [31:0] Mem1D_23_io_output; // @[MemPrimitives.scala 64:21:@32981.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@33469.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@33521.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@33575.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@33627.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@33681.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@33733.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@33787.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@33839.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@33893.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@33945.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@33999.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@34051.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@34105.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@34157.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@34211.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@34263.4]
  wire  StickySelects_16_clock; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_reset; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_io_ins_0; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_io_ins_1; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_io_ins_2; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_io_ins_3; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_io_outs_0; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_io_outs_1; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_io_outs_2; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_16_io_outs_3; // @[MemPrimitives.scala 124:33:@34317.4]
  wire  StickySelects_17_clock; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_reset; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_ins_0; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_ins_1; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_ins_2; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_ins_3; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_ins_4; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_ins_5; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_outs_0; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_outs_1; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_outs_2; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_outs_3; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_outs_4; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_17_io_outs_5; // @[MemPrimitives.scala 124:33:@34369.4]
  wire  StickySelects_18_clock; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_reset; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_io_ins_0; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_io_ins_1; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_io_ins_2; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_io_ins_3; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_io_outs_0; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_io_outs_1; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_io_outs_2; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_18_io_outs_3; // @[MemPrimitives.scala 124:33:@34423.4]
  wire  StickySelects_19_clock; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_reset; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_ins_0; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_ins_1; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_ins_2; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_ins_3; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_ins_4; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_ins_5; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_outs_0; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_outs_1; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_outs_2; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_outs_3; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_outs_4; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_19_io_outs_5; // @[MemPrimitives.scala 124:33:@34475.4]
  wire  StickySelects_20_clock; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_reset; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_io_ins_0; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_io_ins_1; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_io_ins_2; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_io_ins_3; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_io_outs_0; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_io_outs_1; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_io_outs_2; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_20_io_outs_3; // @[MemPrimitives.scala 124:33:@34529.4]
  wire  StickySelects_21_clock; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_reset; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_ins_0; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_ins_1; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_ins_2; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_ins_3; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_ins_4; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_ins_5; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_outs_0; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_outs_1; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_outs_2; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_outs_3; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_outs_4; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_21_io_outs_5; // @[MemPrimitives.scala 124:33:@34581.4]
  wire  StickySelects_22_clock; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_reset; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_io_ins_0; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_io_ins_1; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_io_ins_2; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_io_ins_3; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_io_outs_0; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_io_outs_1; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_io_outs_2; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_22_io_outs_3; // @[MemPrimitives.scala 124:33:@34635.4]
  wire  StickySelects_23_clock; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_reset; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_ins_0; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_ins_1; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_ins_2; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_ins_3; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_ins_4; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_ins_5; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_outs_0; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_outs_1; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_outs_2; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_outs_3; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_outs_4; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  StickySelects_23_io_outs_5; // @[MemPrimitives.scala 124:33:@34687.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@34762.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@34762.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@34762.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@34762.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@34762.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@34770.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@34770.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@34770.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@34770.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@34770.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@34778.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@34778.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@34778.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@34778.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@34778.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@34786.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@34786.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@34786.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@34786.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@34786.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@34794.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@34794.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@34794.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@34794.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@34794.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@34802.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@34802.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@34802.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@34802.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@34802.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@34810.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@34810.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@34810.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@34810.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@34810.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@34818.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@34818.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@34818.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@34818.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@34818.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@34826.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@34826.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@34826.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@34826.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@34826.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@34834.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@34834.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@34834.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@34834.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@34834.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@34842.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@34850.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@34850.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@34850.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@34850.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@34850.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@34906.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@34914.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@34922.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@34922.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@34922.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@34922.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@34922.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@34930.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@34930.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@34930.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@34930.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@34930.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@34938.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@34938.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@34938.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@34938.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@34938.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@34946.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@34946.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@34946.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@34946.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@34946.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@34954.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@34954.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@34954.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@34954.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@34954.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@34962.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@34962.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@34962.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@34962.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@34962.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@34970.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@34978.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@34978.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@34978.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@34978.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@34978.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@34986.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@34986.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@34986.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@34986.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@34986.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@34994.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@34994.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@34994.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@34994.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@34994.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@35050.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@35050.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@35050.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@35050.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@35050.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@35058.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@35058.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@35058.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@35058.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@35058.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@35066.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@35066.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@35066.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@35066.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@35066.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@35074.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@35074.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@35074.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@35074.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@35074.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@35082.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@35082.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@35082.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@35082.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@35082.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@35090.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@35090.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@35090.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@35090.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@35090.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@35098.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@35098.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@35098.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@35098.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@35098.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@35106.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@35106.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@35106.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@35106.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@35106.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@35114.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@35114.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@35114.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@35114.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@35114.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@35122.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@35122.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@35122.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@35122.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@35122.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@35130.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@35130.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@35130.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@35130.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@35130.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@35138.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@35138.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@35138.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@35138.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@35138.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@35194.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@35194.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@35194.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@35194.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@35194.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@35202.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@35202.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@35202.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@35202.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@35202.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@35210.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@35210.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@35210.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@35210.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@35210.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@35218.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@35218.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@35218.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@35218.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@35218.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@35226.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@35226.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@35226.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@35226.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@35226.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@35234.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@35234.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@35234.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@35234.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@35234.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@35242.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@35242.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@35242.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@35242.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@35242.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@35250.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@35258.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@35258.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@35258.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@35258.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@35258.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@35266.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@35266.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@35266.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@35266.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@35266.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@35274.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@35274.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@35274.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@35274.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@35274.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@35282.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@35282.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@35282.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@35282.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@35282.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@35338.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@35338.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@35338.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@35338.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@35338.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@35346.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@35346.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@35346.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@35346.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@35346.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@35354.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@35354.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@35354.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@35354.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@35354.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@35362.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@35362.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@35362.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@35362.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@35362.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@35370.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@35370.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@35370.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@35370.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@35370.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@35378.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@35378.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@35378.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@35378.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@35378.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@35386.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@35386.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@35386.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@35386.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@35386.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@35394.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@35394.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@35394.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@35394.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@35394.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@35402.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@35402.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@35402.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@35402.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@35402.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@35410.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@35410.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@35410.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@35410.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@35410.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@35418.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@35418.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@35418.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@35418.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@35418.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@35426.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@35426.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@35426.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@35426.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@35426.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@35482.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@35482.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@35482.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@35482.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@35482.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@35490.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@35490.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@35490.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@35490.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@35490.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@35498.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@35498.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@35498.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@35498.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@35498.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@35506.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@35506.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@35506.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@35506.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@35506.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@35514.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@35514.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@35514.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@35514.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@35514.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@35522.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@35522.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@35522.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@35522.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@35522.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@35530.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@35530.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@35530.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@35530.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@35530.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@35538.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@35538.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@35538.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@35538.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@35538.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@35546.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@35546.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@35546.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@35546.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@35546.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@35554.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@35554.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@35554.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@35554.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@35554.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@35562.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@35562.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@35562.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@35562.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@35562.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@35570.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@35570.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@35570.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@35570.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@35570.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@35626.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@35626.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@35626.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@35626.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@35626.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@35634.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@35634.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@35634.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@35634.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@35634.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@35642.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@35650.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@35650.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@35650.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@35650.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@35650.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@35658.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@35658.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@35658.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@35658.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@35658.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@35666.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@35666.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@35666.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@35666.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@35666.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@35674.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@35674.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@35674.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@35674.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@35674.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@35682.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@35682.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@35682.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@35682.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@35682.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@35690.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@35698.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@35698.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@35698.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@35698.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@35698.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@35706.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@35706.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@35706.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@35706.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@35706.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@35714.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@35714.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@35714.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@35714.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@35714.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@35770.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@35770.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@35770.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@35770.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@35770.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@35778.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@35778.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@35778.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@35778.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@35778.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@35786.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@35786.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@35786.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@35786.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@35786.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@35794.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@35794.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@35794.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@35794.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@35794.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@35802.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@35802.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@35802.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@35802.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@35802.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@35810.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@35810.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@35810.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@35810.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@35810.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@35818.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@35818.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@35818.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@35818.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@35818.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@35826.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@35826.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@35826.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@35826.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@35826.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@35834.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@35834.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@35834.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@35834.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@35834.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@35842.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@35842.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@35842.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@35842.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@35842.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@35850.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@35850.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@35850.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@35850.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@35850.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@35858.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@35858.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@35858.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@35858.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@35858.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@35914.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@35914.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@35914.4]
  wire  RetimeWrapper_96_io_in; // @[package.scala 93:22:@35914.4]
  wire  RetimeWrapper_96_io_out; // @[package.scala 93:22:@35914.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@35922.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@35922.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@35922.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@35922.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@35922.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@35930.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@35930.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@35930.4]
  wire  RetimeWrapper_98_io_in; // @[package.scala 93:22:@35930.4]
  wire  RetimeWrapper_98_io_out; // @[package.scala 93:22:@35930.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@35938.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@35938.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@35938.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@35938.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@35938.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@35946.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@35946.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@35946.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@35946.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@35946.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@35954.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@35954.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@35954.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@35954.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@35954.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@35962.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@35962.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@35962.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@35962.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@35962.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@35970.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@35970.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@35970.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@35970.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@35970.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@35978.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@35978.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@35978.4]
  wire  RetimeWrapper_104_io_in; // @[package.scala 93:22:@35978.4]
  wire  RetimeWrapper_104_io_out; // @[package.scala 93:22:@35978.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@35986.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@35986.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@35986.4]
  wire  RetimeWrapper_105_io_in; // @[package.scala 93:22:@35986.4]
  wire  RetimeWrapper_105_io_out; // @[package.scala 93:22:@35986.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@35994.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@35994.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@35994.4]
  wire  RetimeWrapper_106_io_in; // @[package.scala 93:22:@35994.4]
  wire  RetimeWrapper_106_io_out; // @[package.scala 93:22:@35994.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@36002.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@36002.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@36002.4]
  wire  RetimeWrapper_107_io_in; // @[package.scala 93:22:@36002.4]
  wire  RetimeWrapper_107_io_out; // @[package.scala 93:22:@36002.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@36058.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@36058.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@36058.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@36058.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@36058.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@36066.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@36066.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@36066.4]
  wire  RetimeWrapper_109_io_in; // @[package.scala 93:22:@36066.4]
  wire  RetimeWrapper_109_io_out; // @[package.scala 93:22:@36066.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@36074.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@36074.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@36074.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@36074.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@36074.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@36082.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@36082.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@36082.4]
  wire  RetimeWrapper_111_io_in; // @[package.scala 93:22:@36082.4]
  wire  RetimeWrapper_111_io_out; // @[package.scala 93:22:@36082.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@36090.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@36090.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@36090.4]
  wire  RetimeWrapper_112_io_in; // @[package.scala 93:22:@36090.4]
  wire  RetimeWrapper_112_io_out; // @[package.scala 93:22:@36090.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@36098.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@36098.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@36098.4]
  wire  RetimeWrapper_113_io_in; // @[package.scala 93:22:@36098.4]
  wire  RetimeWrapper_113_io_out; // @[package.scala 93:22:@36098.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@36106.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@36106.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@36106.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@36106.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@36106.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@36114.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@36114.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@36114.4]
  wire  RetimeWrapper_115_io_in; // @[package.scala 93:22:@36114.4]
  wire  RetimeWrapper_115_io_out; // @[package.scala 93:22:@36114.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_116_io_in; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_116_io_out; // @[package.scala 93:22:@36122.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@36130.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@36130.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@36130.4]
  wire  RetimeWrapper_117_io_in; // @[package.scala 93:22:@36130.4]
  wire  RetimeWrapper_117_io_out; // @[package.scala 93:22:@36130.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@36138.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@36138.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@36138.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@36138.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@36138.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@36146.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@36146.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@36146.4]
  wire  RetimeWrapper_119_io_in; // @[package.scala 93:22:@36146.4]
  wire  RetimeWrapper_119_io_out; // @[package.scala 93:22:@36146.4]
  wire  _T_460; // @[MemPrimitives.scala 82:210:@32997.4]
  wire  _T_462; // @[MemPrimitives.scala 82:210:@32998.4]
  wire  _T_463; // @[MemPrimitives.scala 82:228:@32999.4]
  wire  _T_464; // @[MemPrimitives.scala 83:102:@33000.4]
  wire  _T_466; // @[MemPrimitives.scala 82:210:@33001.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@33002.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@33003.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@33004.4]
  wire [41:0] _T_472; // @[Cat.scala 30:58:@33006.4]
  wire [41:0] _T_474; // @[Cat.scala 30:58:@33008.4]
  wire [41:0] _T_475; // @[Mux.scala 31:69:@33009.4]
  wire  _T_480; // @[MemPrimitives.scala 82:210:@33016.4]
  wire  _T_482; // @[MemPrimitives.scala 82:210:@33017.4]
  wire  _T_483; // @[MemPrimitives.scala 82:228:@33018.4]
  wire  _T_484; // @[MemPrimitives.scala 83:102:@33019.4]
  wire  _T_486; // @[MemPrimitives.scala 82:210:@33020.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@33021.4]
  wire  _T_489; // @[MemPrimitives.scala 82:228:@33022.4]
  wire  _T_490; // @[MemPrimitives.scala 83:102:@33023.4]
  wire [41:0] _T_492; // @[Cat.scala 30:58:@33025.4]
  wire [41:0] _T_494; // @[Cat.scala 30:58:@33027.4]
  wire [41:0] _T_495; // @[Mux.scala 31:69:@33028.4]
  wire  _T_502; // @[MemPrimitives.scala 82:210:@33036.4]
  wire  _T_503; // @[MemPrimitives.scala 82:228:@33037.4]
  wire  _T_504; // @[MemPrimitives.scala 83:102:@33038.4]
  wire  _T_508; // @[MemPrimitives.scala 82:210:@33040.4]
  wire  _T_509; // @[MemPrimitives.scala 82:228:@33041.4]
  wire  _T_510; // @[MemPrimitives.scala 83:102:@33042.4]
  wire [41:0] _T_512; // @[Cat.scala 30:58:@33044.4]
  wire [41:0] _T_514; // @[Cat.scala 30:58:@33046.4]
  wire [41:0] _T_515; // @[Mux.scala 31:69:@33047.4]
  wire  _T_522; // @[MemPrimitives.scala 82:210:@33055.4]
  wire  _T_523; // @[MemPrimitives.scala 82:228:@33056.4]
  wire  _T_524; // @[MemPrimitives.scala 83:102:@33057.4]
  wire  _T_528; // @[MemPrimitives.scala 82:210:@33059.4]
  wire  _T_529; // @[MemPrimitives.scala 82:228:@33060.4]
  wire  _T_530; // @[MemPrimitives.scala 83:102:@33061.4]
  wire [41:0] _T_532; // @[Cat.scala 30:58:@33063.4]
  wire [41:0] _T_534; // @[Cat.scala 30:58:@33065.4]
  wire [41:0] _T_535; // @[Mux.scala 31:69:@33066.4]
  wire  _T_542; // @[MemPrimitives.scala 82:210:@33074.4]
  wire  _T_543; // @[MemPrimitives.scala 82:228:@33075.4]
  wire  _T_544; // @[MemPrimitives.scala 83:102:@33076.4]
  wire  _T_548; // @[MemPrimitives.scala 82:210:@33078.4]
  wire  _T_549; // @[MemPrimitives.scala 82:228:@33079.4]
  wire  _T_550; // @[MemPrimitives.scala 83:102:@33080.4]
  wire [41:0] _T_552; // @[Cat.scala 30:58:@33082.4]
  wire [41:0] _T_554; // @[Cat.scala 30:58:@33084.4]
  wire [41:0] _T_555; // @[Mux.scala 31:69:@33085.4]
  wire  _T_562; // @[MemPrimitives.scala 82:210:@33093.4]
  wire  _T_563; // @[MemPrimitives.scala 82:228:@33094.4]
  wire  _T_564; // @[MemPrimitives.scala 83:102:@33095.4]
  wire  _T_568; // @[MemPrimitives.scala 82:210:@33097.4]
  wire  _T_569; // @[MemPrimitives.scala 82:228:@33098.4]
  wire  _T_570; // @[MemPrimitives.scala 83:102:@33099.4]
  wire [41:0] _T_572; // @[Cat.scala 30:58:@33101.4]
  wire [41:0] _T_574; // @[Cat.scala 30:58:@33103.4]
  wire [41:0] _T_575; // @[Mux.scala 31:69:@33104.4]
  wire  _T_580; // @[MemPrimitives.scala 82:210:@33111.4]
  wire  _T_583; // @[MemPrimitives.scala 82:228:@33113.4]
  wire  _T_584; // @[MemPrimitives.scala 83:102:@33114.4]
  wire  _T_586; // @[MemPrimitives.scala 82:210:@33115.4]
  wire  _T_589; // @[MemPrimitives.scala 82:228:@33117.4]
  wire  _T_590; // @[MemPrimitives.scala 83:102:@33118.4]
  wire [41:0] _T_592; // @[Cat.scala 30:58:@33120.4]
  wire [41:0] _T_594; // @[Cat.scala 30:58:@33122.4]
  wire [41:0] _T_595; // @[Mux.scala 31:69:@33123.4]
  wire  _T_600; // @[MemPrimitives.scala 82:210:@33130.4]
  wire  _T_603; // @[MemPrimitives.scala 82:228:@33132.4]
  wire  _T_604; // @[MemPrimitives.scala 83:102:@33133.4]
  wire  _T_606; // @[MemPrimitives.scala 82:210:@33134.4]
  wire  _T_609; // @[MemPrimitives.scala 82:228:@33136.4]
  wire  _T_610; // @[MemPrimitives.scala 83:102:@33137.4]
  wire [41:0] _T_612; // @[Cat.scala 30:58:@33139.4]
  wire [41:0] _T_614; // @[Cat.scala 30:58:@33141.4]
  wire [41:0] _T_615; // @[Mux.scala 31:69:@33142.4]
  wire  _T_623; // @[MemPrimitives.scala 82:228:@33151.4]
  wire  _T_624; // @[MemPrimitives.scala 83:102:@33152.4]
  wire  _T_629; // @[MemPrimitives.scala 82:228:@33155.4]
  wire  _T_630; // @[MemPrimitives.scala 83:102:@33156.4]
  wire [41:0] _T_632; // @[Cat.scala 30:58:@33158.4]
  wire [41:0] _T_634; // @[Cat.scala 30:58:@33160.4]
  wire [41:0] _T_635; // @[Mux.scala 31:69:@33161.4]
  wire  _T_643; // @[MemPrimitives.scala 82:228:@33170.4]
  wire  _T_644; // @[MemPrimitives.scala 83:102:@33171.4]
  wire  _T_649; // @[MemPrimitives.scala 82:228:@33174.4]
  wire  _T_650; // @[MemPrimitives.scala 83:102:@33175.4]
  wire [41:0] _T_652; // @[Cat.scala 30:58:@33177.4]
  wire [41:0] _T_654; // @[Cat.scala 30:58:@33179.4]
  wire [41:0] _T_655; // @[Mux.scala 31:69:@33180.4]
  wire  _T_663; // @[MemPrimitives.scala 82:228:@33189.4]
  wire  _T_664; // @[MemPrimitives.scala 83:102:@33190.4]
  wire  _T_669; // @[MemPrimitives.scala 82:228:@33193.4]
  wire  _T_670; // @[MemPrimitives.scala 83:102:@33194.4]
  wire [41:0] _T_672; // @[Cat.scala 30:58:@33196.4]
  wire [41:0] _T_674; // @[Cat.scala 30:58:@33198.4]
  wire [41:0] _T_675; // @[Mux.scala 31:69:@33199.4]
  wire  _T_683; // @[MemPrimitives.scala 82:228:@33208.4]
  wire  _T_684; // @[MemPrimitives.scala 83:102:@33209.4]
  wire  _T_689; // @[MemPrimitives.scala 82:228:@33212.4]
  wire  _T_690; // @[MemPrimitives.scala 83:102:@33213.4]
  wire [41:0] _T_692; // @[Cat.scala 30:58:@33215.4]
  wire [41:0] _T_694; // @[Cat.scala 30:58:@33217.4]
  wire [41:0] _T_695; // @[Mux.scala 31:69:@33218.4]
  wire  _T_700; // @[MemPrimitives.scala 82:210:@33225.4]
  wire  _T_703; // @[MemPrimitives.scala 82:228:@33227.4]
  wire  _T_704; // @[MemPrimitives.scala 83:102:@33228.4]
  wire  _T_706; // @[MemPrimitives.scala 82:210:@33229.4]
  wire  _T_709; // @[MemPrimitives.scala 82:228:@33231.4]
  wire  _T_710; // @[MemPrimitives.scala 83:102:@33232.4]
  wire [41:0] _T_712; // @[Cat.scala 30:58:@33234.4]
  wire [41:0] _T_714; // @[Cat.scala 30:58:@33236.4]
  wire [41:0] _T_715; // @[Mux.scala 31:69:@33237.4]
  wire  _T_720; // @[MemPrimitives.scala 82:210:@33244.4]
  wire  _T_723; // @[MemPrimitives.scala 82:228:@33246.4]
  wire  _T_724; // @[MemPrimitives.scala 83:102:@33247.4]
  wire  _T_726; // @[MemPrimitives.scala 82:210:@33248.4]
  wire  _T_729; // @[MemPrimitives.scala 82:228:@33250.4]
  wire  _T_730; // @[MemPrimitives.scala 83:102:@33251.4]
  wire [41:0] _T_732; // @[Cat.scala 30:58:@33253.4]
  wire [41:0] _T_734; // @[Cat.scala 30:58:@33255.4]
  wire [41:0] _T_735; // @[Mux.scala 31:69:@33256.4]
  wire  _T_743; // @[MemPrimitives.scala 82:228:@33265.4]
  wire  _T_744; // @[MemPrimitives.scala 83:102:@33266.4]
  wire  _T_749; // @[MemPrimitives.scala 82:228:@33269.4]
  wire  _T_750; // @[MemPrimitives.scala 83:102:@33270.4]
  wire [41:0] _T_752; // @[Cat.scala 30:58:@33272.4]
  wire [41:0] _T_754; // @[Cat.scala 30:58:@33274.4]
  wire [41:0] _T_755; // @[Mux.scala 31:69:@33275.4]
  wire  _T_763; // @[MemPrimitives.scala 82:228:@33284.4]
  wire  _T_764; // @[MemPrimitives.scala 83:102:@33285.4]
  wire  _T_769; // @[MemPrimitives.scala 82:228:@33288.4]
  wire  _T_770; // @[MemPrimitives.scala 83:102:@33289.4]
  wire [41:0] _T_772; // @[Cat.scala 30:58:@33291.4]
  wire [41:0] _T_774; // @[Cat.scala 30:58:@33293.4]
  wire [41:0] _T_775; // @[Mux.scala 31:69:@33294.4]
  wire  _T_783; // @[MemPrimitives.scala 82:228:@33303.4]
  wire  _T_784; // @[MemPrimitives.scala 83:102:@33304.4]
  wire  _T_789; // @[MemPrimitives.scala 82:228:@33307.4]
  wire  _T_790; // @[MemPrimitives.scala 83:102:@33308.4]
  wire [41:0] _T_792; // @[Cat.scala 30:58:@33310.4]
  wire [41:0] _T_794; // @[Cat.scala 30:58:@33312.4]
  wire [41:0] _T_795; // @[Mux.scala 31:69:@33313.4]
  wire  _T_803; // @[MemPrimitives.scala 82:228:@33322.4]
  wire  _T_804; // @[MemPrimitives.scala 83:102:@33323.4]
  wire  _T_809; // @[MemPrimitives.scala 82:228:@33326.4]
  wire  _T_810; // @[MemPrimitives.scala 83:102:@33327.4]
  wire [41:0] _T_812; // @[Cat.scala 30:58:@33329.4]
  wire [41:0] _T_814; // @[Cat.scala 30:58:@33331.4]
  wire [41:0] _T_815; // @[Mux.scala 31:69:@33332.4]
  wire  _T_820; // @[MemPrimitives.scala 82:210:@33339.4]
  wire  _T_823; // @[MemPrimitives.scala 82:228:@33341.4]
  wire  _T_824; // @[MemPrimitives.scala 83:102:@33342.4]
  wire  _T_826; // @[MemPrimitives.scala 82:210:@33343.4]
  wire  _T_829; // @[MemPrimitives.scala 82:228:@33345.4]
  wire  _T_830; // @[MemPrimitives.scala 83:102:@33346.4]
  wire [41:0] _T_832; // @[Cat.scala 30:58:@33348.4]
  wire [41:0] _T_834; // @[Cat.scala 30:58:@33350.4]
  wire [41:0] _T_835; // @[Mux.scala 31:69:@33351.4]
  wire  _T_840; // @[MemPrimitives.scala 82:210:@33358.4]
  wire  _T_843; // @[MemPrimitives.scala 82:228:@33360.4]
  wire  _T_844; // @[MemPrimitives.scala 83:102:@33361.4]
  wire  _T_846; // @[MemPrimitives.scala 82:210:@33362.4]
  wire  _T_849; // @[MemPrimitives.scala 82:228:@33364.4]
  wire  _T_850; // @[MemPrimitives.scala 83:102:@33365.4]
  wire [41:0] _T_852; // @[Cat.scala 30:58:@33367.4]
  wire [41:0] _T_854; // @[Cat.scala 30:58:@33369.4]
  wire [41:0] _T_855; // @[Mux.scala 31:69:@33370.4]
  wire  _T_863; // @[MemPrimitives.scala 82:228:@33379.4]
  wire  _T_864; // @[MemPrimitives.scala 83:102:@33380.4]
  wire  _T_869; // @[MemPrimitives.scala 82:228:@33383.4]
  wire  _T_870; // @[MemPrimitives.scala 83:102:@33384.4]
  wire [41:0] _T_872; // @[Cat.scala 30:58:@33386.4]
  wire [41:0] _T_874; // @[Cat.scala 30:58:@33388.4]
  wire [41:0] _T_875; // @[Mux.scala 31:69:@33389.4]
  wire  _T_883; // @[MemPrimitives.scala 82:228:@33398.4]
  wire  _T_884; // @[MemPrimitives.scala 83:102:@33399.4]
  wire  _T_889; // @[MemPrimitives.scala 82:228:@33402.4]
  wire  _T_890; // @[MemPrimitives.scala 83:102:@33403.4]
  wire [41:0] _T_892; // @[Cat.scala 30:58:@33405.4]
  wire [41:0] _T_894; // @[Cat.scala 30:58:@33407.4]
  wire [41:0] _T_895; // @[Mux.scala 31:69:@33408.4]
  wire  _T_903; // @[MemPrimitives.scala 82:228:@33417.4]
  wire  _T_904; // @[MemPrimitives.scala 83:102:@33418.4]
  wire  _T_909; // @[MemPrimitives.scala 82:228:@33421.4]
  wire  _T_910; // @[MemPrimitives.scala 83:102:@33422.4]
  wire [41:0] _T_912; // @[Cat.scala 30:58:@33424.4]
  wire [41:0] _T_914; // @[Cat.scala 30:58:@33426.4]
  wire [41:0] _T_915; // @[Mux.scala 31:69:@33427.4]
  wire  _T_923; // @[MemPrimitives.scala 82:228:@33436.4]
  wire  _T_924; // @[MemPrimitives.scala 83:102:@33437.4]
  wire  _T_929; // @[MemPrimitives.scala 82:228:@33440.4]
  wire  _T_930; // @[MemPrimitives.scala 83:102:@33441.4]
  wire [41:0] _T_932; // @[Cat.scala 30:58:@33443.4]
  wire [41:0] _T_934; // @[Cat.scala 30:58:@33445.4]
  wire [41:0] _T_935; // @[Mux.scala 31:69:@33446.4]
  wire  _T_940; // @[MemPrimitives.scala 110:210:@33453.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@33454.4]
  wire  _T_943; // @[MemPrimitives.scala 110:228:@33455.4]
  wire  _T_946; // @[MemPrimitives.scala 110:210:@33457.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@33458.4]
  wire  _T_949; // @[MemPrimitives.scala 110:228:@33459.4]
  wire  _T_952; // @[MemPrimitives.scala 110:210:@33461.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@33462.4]
  wire  _T_955; // @[MemPrimitives.scala 110:228:@33463.4]
  wire  _T_958; // @[MemPrimitives.scala 110:210:@33465.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@33466.4]
  wire  _T_961; // @[MemPrimitives.scala 110:228:@33467.4]
  wire  _T_963; // @[MemPrimitives.scala 126:35:@33476.4]
  wire  _T_964; // @[MemPrimitives.scala 126:35:@33477.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@33478.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@33479.4]
  wire [10:0] _T_968; // @[Cat.scala 30:58:@33481.4]
  wire [10:0] _T_970; // @[Cat.scala 30:58:@33483.4]
  wire [10:0] _T_972; // @[Cat.scala 30:58:@33485.4]
  wire [10:0] _T_974; // @[Cat.scala 30:58:@33487.4]
  wire [10:0] _T_975; // @[Mux.scala 31:69:@33488.4]
  wire [10:0] _T_976; // @[Mux.scala 31:69:@33489.4]
  wire [10:0] _T_977; // @[Mux.scala 31:69:@33490.4]
  wire  _T_982; // @[MemPrimitives.scala 110:210:@33497.4]
  wire  _T_984; // @[MemPrimitives.scala 110:210:@33498.4]
  wire  _T_985; // @[MemPrimitives.scala 110:228:@33499.4]
  wire  _T_988; // @[MemPrimitives.scala 110:210:@33501.4]
  wire  _T_990; // @[MemPrimitives.scala 110:210:@33502.4]
  wire  _T_991; // @[MemPrimitives.scala 110:228:@33503.4]
  wire  _T_994; // @[MemPrimitives.scala 110:210:@33505.4]
  wire  _T_996; // @[MemPrimitives.scala 110:210:@33506.4]
  wire  _T_997; // @[MemPrimitives.scala 110:228:@33507.4]
  wire  _T_1000; // @[MemPrimitives.scala 110:210:@33509.4]
  wire  _T_1002; // @[MemPrimitives.scala 110:210:@33510.4]
  wire  _T_1003; // @[MemPrimitives.scala 110:228:@33511.4]
  wire  _T_1006; // @[MemPrimitives.scala 110:210:@33513.4]
  wire  _T_1008; // @[MemPrimitives.scala 110:210:@33514.4]
  wire  _T_1009; // @[MemPrimitives.scala 110:228:@33515.4]
  wire  _T_1012; // @[MemPrimitives.scala 110:210:@33517.4]
  wire  _T_1014; // @[MemPrimitives.scala 110:210:@33518.4]
  wire  _T_1015; // @[MemPrimitives.scala 110:228:@33519.4]
  wire  _T_1017; // @[MemPrimitives.scala 126:35:@33530.4]
  wire  _T_1018; // @[MemPrimitives.scala 126:35:@33531.4]
  wire  _T_1019; // @[MemPrimitives.scala 126:35:@33532.4]
  wire  _T_1020; // @[MemPrimitives.scala 126:35:@33533.4]
  wire  _T_1021; // @[MemPrimitives.scala 126:35:@33534.4]
  wire  _T_1022; // @[MemPrimitives.scala 126:35:@33535.4]
  wire [10:0] _T_1024; // @[Cat.scala 30:58:@33537.4]
  wire [10:0] _T_1026; // @[Cat.scala 30:58:@33539.4]
  wire [10:0] _T_1028; // @[Cat.scala 30:58:@33541.4]
  wire [10:0] _T_1030; // @[Cat.scala 30:58:@33543.4]
  wire [10:0] _T_1032; // @[Cat.scala 30:58:@33545.4]
  wire [10:0] _T_1034; // @[Cat.scala 30:58:@33547.4]
  wire [10:0] _T_1035; // @[Mux.scala 31:69:@33548.4]
  wire [10:0] _T_1036; // @[Mux.scala 31:69:@33549.4]
  wire [10:0] _T_1037; // @[Mux.scala 31:69:@33550.4]
  wire [10:0] _T_1038; // @[Mux.scala 31:69:@33551.4]
  wire [10:0] _T_1039; // @[Mux.scala 31:69:@33552.4]
  wire  _T_1046; // @[MemPrimitives.scala 110:210:@33560.4]
  wire  _T_1047; // @[MemPrimitives.scala 110:228:@33561.4]
  wire  _T_1052; // @[MemPrimitives.scala 110:210:@33564.4]
  wire  _T_1053; // @[MemPrimitives.scala 110:228:@33565.4]
  wire  _T_1058; // @[MemPrimitives.scala 110:210:@33568.4]
  wire  _T_1059; // @[MemPrimitives.scala 110:228:@33569.4]
  wire  _T_1064; // @[MemPrimitives.scala 110:210:@33572.4]
  wire  _T_1065; // @[MemPrimitives.scala 110:228:@33573.4]
  wire  _T_1067; // @[MemPrimitives.scala 126:35:@33582.4]
  wire  _T_1068; // @[MemPrimitives.scala 126:35:@33583.4]
  wire  _T_1069; // @[MemPrimitives.scala 126:35:@33584.4]
  wire  _T_1070; // @[MemPrimitives.scala 126:35:@33585.4]
  wire [10:0] _T_1072; // @[Cat.scala 30:58:@33587.4]
  wire [10:0] _T_1074; // @[Cat.scala 30:58:@33589.4]
  wire [10:0] _T_1076; // @[Cat.scala 30:58:@33591.4]
  wire [10:0] _T_1078; // @[Cat.scala 30:58:@33593.4]
  wire [10:0] _T_1079; // @[Mux.scala 31:69:@33594.4]
  wire [10:0] _T_1080; // @[Mux.scala 31:69:@33595.4]
  wire [10:0] _T_1081; // @[Mux.scala 31:69:@33596.4]
  wire  _T_1088; // @[MemPrimitives.scala 110:210:@33604.4]
  wire  _T_1089; // @[MemPrimitives.scala 110:228:@33605.4]
  wire  _T_1094; // @[MemPrimitives.scala 110:210:@33608.4]
  wire  _T_1095; // @[MemPrimitives.scala 110:228:@33609.4]
  wire  _T_1100; // @[MemPrimitives.scala 110:210:@33612.4]
  wire  _T_1101; // @[MemPrimitives.scala 110:228:@33613.4]
  wire  _T_1106; // @[MemPrimitives.scala 110:210:@33616.4]
  wire  _T_1107; // @[MemPrimitives.scala 110:228:@33617.4]
  wire  _T_1112; // @[MemPrimitives.scala 110:210:@33620.4]
  wire  _T_1113; // @[MemPrimitives.scala 110:228:@33621.4]
  wire  _T_1118; // @[MemPrimitives.scala 110:210:@33624.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@33625.4]
  wire  _T_1121; // @[MemPrimitives.scala 126:35:@33636.4]
  wire  _T_1122; // @[MemPrimitives.scala 126:35:@33637.4]
  wire  _T_1123; // @[MemPrimitives.scala 126:35:@33638.4]
  wire  _T_1124; // @[MemPrimitives.scala 126:35:@33639.4]
  wire  _T_1125; // @[MemPrimitives.scala 126:35:@33640.4]
  wire  _T_1126; // @[MemPrimitives.scala 126:35:@33641.4]
  wire [10:0] _T_1128; // @[Cat.scala 30:58:@33643.4]
  wire [10:0] _T_1130; // @[Cat.scala 30:58:@33645.4]
  wire [10:0] _T_1132; // @[Cat.scala 30:58:@33647.4]
  wire [10:0] _T_1134; // @[Cat.scala 30:58:@33649.4]
  wire [10:0] _T_1136; // @[Cat.scala 30:58:@33651.4]
  wire [10:0] _T_1138; // @[Cat.scala 30:58:@33653.4]
  wire [10:0] _T_1139; // @[Mux.scala 31:69:@33654.4]
  wire [10:0] _T_1140; // @[Mux.scala 31:69:@33655.4]
  wire [10:0] _T_1141; // @[Mux.scala 31:69:@33656.4]
  wire [10:0] _T_1142; // @[Mux.scala 31:69:@33657.4]
  wire [10:0] _T_1143; // @[Mux.scala 31:69:@33658.4]
  wire  _T_1150; // @[MemPrimitives.scala 110:210:@33666.4]
  wire  _T_1151; // @[MemPrimitives.scala 110:228:@33667.4]
  wire  _T_1156; // @[MemPrimitives.scala 110:210:@33670.4]
  wire  _T_1157; // @[MemPrimitives.scala 110:228:@33671.4]
  wire  _T_1162; // @[MemPrimitives.scala 110:210:@33674.4]
  wire  _T_1163; // @[MemPrimitives.scala 110:228:@33675.4]
  wire  _T_1168; // @[MemPrimitives.scala 110:210:@33678.4]
  wire  _T_1169; // @[MemPrimitives.scala 110:228:@33679.4]
  wire  _T_1171; // @[MemPrimitives.scala 126:35:@33688.4]
  wire  _T_1172; // @[MemPrimitives.scala 126:35:@33689.4]
  wire  _T_1173; // @[MemPrimitives.scala 126:35:@33690.4]
  wire  _T_1174; // @[MemPrimitives.scala 126:35:@33691.4]
  wire [10:0] _T_1176; // @[Cat.scala 30:58:@33693.4]
  wire [10:0] _T_1178; // @[Cat.scala 30:58:@33695.4]
  wire [10:0] _T_1180; // @[Cat.scala 30:58:@33697.4]
  wire [10:0] _T_1182; // @[Cat.scala 30:58:@33699.4]
  wire [10:0] _T_1183; // @[Mux.scala 31:69:@33700.4]
  wire [10:0] _T_1184; // @[Mux.scala 31:69:@33701.4]
  wire [10:0] _T_1185; // @[Mux.scala 31:69:@33702.4]
  wire  _T_1192; // @[MemPrimitives.scala 110:210:@33710.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@33711.4]
  wire  _T_1198; // @[MemPrimitives.scala 110:210:@33714.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@33715.4]
  wire  _T_1204; // @[MemPrimitives.scala 110:210:@33718.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@33719.4]
  wire  _T_1210; // @[MemPrimitives.scala 110:210:@33722.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@33723.4]
  wire  _T_1216; // @[MemPrimitives.scala 110:210:@33726.4]
  wire  _T_1217; // @[MemPrimitives.scala 110:228:@33727.4]
  wire  _T_1222; // @[MemPrimitives.scala 110:210:@33730.4]
  wire  _T_1223; // @[MemPrimitives.scala 110:228:@33731.4]
  wire  _T_1225; // @[MemPrimitives.scala 126:35:@33742.4]
  wire  _T_1226; // @[MemPrimitives.scala 126:35:@33743.4]
  wire  _T_1227; // @[MemPrimitives.scala 126:35:@33744.4]
  wire  _T_1228; // @[MemPrimitives.scala 126:35:@33745.4]
  wire  _T_1229; // @[MemPrimitives.scala 126:35:@33746.4]
  wire  _T_1230; // @[MemPrimitives.scala 126:35:@33747.4]
  wire [10:0] _T_1232; // @[Cat.scala 30:58:@33749.4]
  wire [10:0] _T_1234; // @[Cat.scala 30:58:@33751.4]
  wire [10:0] _T_1236; // @[Cat.scala 30:58:@33753.4]
  wire [10:0] _T_1238; // @[Cat.scala 30:58:@33755.4]
  wire [10:0] _T_1240; // @[Cat.scala 30:58:@33757.4]
  wire [10:0] _T_1242; // @[Cat.scala 30:58:@33759.4]
  wire [10:0] _T_1243; // @[Mux.scala 31:69:@33760.4]
  wire [10:0] _T_1244; // @[Mux.scala 31:69:@33761.4]
  wire [10:0] _T_1245; // @[Mux.scala 31:69:@33762.4]
  wire [10:0] _T_1246; // @[Mux.scala 31:69:@33763.4]
  wire [10:0] _T_1247; // @[Mux.scala 31:69:@33764.4]
  wire  _T_1252; // @[MemPrimitives.scala 110:210:@33771.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@33773.4]
  wire  _T_1258; // @[MemPrimitives.scala 110:210:@33775.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@33777.4]
  wire  _T_1264; // @[MemPrimitives.scala 110:210:@33779.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@33781.4]
  wire  _T_1270; // @[MemPrimitives.scala 110:210:@33783.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@33785.4]
  wire  _T_1275; // @[MemPrimitives.scala 126:35:@33794.4]
  wire  _T_1276; // @[MemPrimitives.scala 126:35:@33795.4]
  wire  _T_1277; // @[MemPrimitives.scala 126:35:@33796.4]
  wire  _T_1278; // @[MemPrimitives.scala 126:35:@33797.4]
  wire [10:0] _T_1280; // @[Cat.scala 30:58:@33799.4]
  wire [10:0] _T_1282; // @[Cat.scala 30:58:@33801.4]
  wire [10:0] _T_1284; // @[Cat.scala 30:58:@33803.4]
  wire [10:0] _T_1286; // @[Cat.scala 30:58:@33805.4]
  wire [10:0] _T_1287; // @[Mux.scala 31:69:@33806.4]
  wire [10:0] _T_1288; // @[Mux.scala 31:69:@33807.4]
  wire [10:0] _T_1289; // @[Mux.scala 31:69:@33808.4]
  wire  _T_1294; // @[MemPrimitives.scala 110:210:@33815.4]
  wire  _T_1297; // @[MemPrimitives.scala 110:228:@33817.4]
  wire  _T_1300; // @[MemPrimitives.scala 110:210:@33819.4]
  wire  _T_1303; // @[MemPrimitives.scala 110:228:@33821.4]
  wire  _T_1306; // @[MemPrimitives.scala 110:210:@33823.4]
  wire  _T_1309; // @[MemPrimitives.scala 110:228:@33825.4]
  wire  _T_1312; // @[MemPrimitives.scala 110:210:@33827.4]
  wire  _T_1315; // @[MemPrimitives.scala 110:228:@33829.4]
  wire  _T_1318; // @[MemPrimitives.scala 110:210:@33831.4]
  wire  _T_1321; // @[MemPrimitives.scala 110:228:@33833.4]
  wire  _T_1324; // @[MemPrimitives.scala 110:210:@33835.4]
  wire  _T_1327; // @[MemPrimitives.scala 110:228:@33837.4]
  wire  _T_1329; // @[MemPrimitives.scala 126:35:@33848.4]
  wire  _T_1330; // @[MemPrimitives.scala 126:35:@33849.4]
  wire  _T_1331; // @[MemPrimitives.scala 126:35:@33850.4]
  wire  _T_1332; // @[MemPrimitives.scala 126:35:@33851.4]
  wire  _T_1333; // @[MemPrimitives.scala 126:35:@33852.4]
  wire  _T_1334; // @[MemPrimitives.scala 126:35:@33853.4]
  wire [10:0] _T_1336; // @[Cat.scala 30:58:@33855.4]
  wire [10:0] _T_1338; // @[Cat.scala 30:58:@33857.4]
  wire [10:0] _T_1340; // @[Cat.scala 30:58:@33859.4]
  wire [10:0] _T_1342; // @[Cat.scala 30:58:@33861.4]
  wire [10:0] _T_1344; // @[Cat.scala 30:58:@33863.4]
  wire [10:0] _T_1346; // @[Cat.scala 30:58:@33865.4]
  wire [10:0] _T_1347; // @[Mux.scala 31:69:@33866.4]
  wire [10:0] _T_1348; // @[Mux.scala 31:69:@33867.4]
  wire [10:0] _T_1349; // @[Mux.scala 31:69:@33868.4]
  wire [10:0] _T_1350; // @[Mux.scala 31:69:@33869.4]
  wire [10:0] _T_1351; // @[Mux.scala 31:69:@33870.4]
  wire  _T_1359; // @[MemPrimitives.scala 110:228:@33879.4]
  wire  _T_1365; // @[MemPrimitives.scala 110:228:@33883.4]
  wire  _T_1371; // @[MemPrimitives.scala 110:228:@33887.4]
  wire  _T_1377; // @[MemPrimitives.scala 110:228:@33891.4]
  wire  _T_1379; // @[MemPrimitives.scala 126:35:@33900.4]
  wire  _T_1380; // @[MemPrimitives.scala 126:35:@33901.4]
  wire  _T_1381; // @[MemPrimitives.scala 126:35:@33902.4]
  wire  _T_1382; // @[MemPrimitives.scala 126:35:@33903.4]
  wire [10:0] _T_1384; // @[Cat.scala 30:58:@33905.4]
  wire [10:0] _T_1386; // @[Cat.scala 30:58:@33907.4]
  wire [10:0] _T_1388; // @[Cat.scala 30:58:@33909.4]
  wire [10:0] _T_1390; // @[Cat.scala 30:58:@33911.4]
  wire [10:0] _T_1391; // @[Mux.scala 31:69:@33912.4]
  wire [10:0] _T_1392; // @[Mux.scala 31:69:@33913.4]
  wire [10:0] _T_1393; // @[Mux.scala 31:69:@33914.4]
  wire  _T_1401; // @[MemPrimitives.scala 110:228:@33923.4]
  wire  _T_1407; // @[MemPrimitives.scala 110:228:@33927.4]
  wire  _T_1413; // @[MemPrimitives.scala 110:228:@33931.4]
  wire  _T_1419; // @[MemPrimitives.scala 110:228:@33935.4]
  wire  _T_1425; // @[MemPrimitives.scala 110:228:@33939.4]
  wire  _T_1431; // @[MemPrimitives.scala 110:228:@33943.4]
  wire  _T_1433; // @[MemPrimitives.scala 126:35:@33954.4]
  wire  _T_1434; // @[MemPrimitives.scala 126:35:@33955.4]
  wire  _T_1435; // @[MemPrimitives.scala 126:35:@33956.4]
  wire  _T_1436; // @[MemPrimitives.scala 126:35:@33957.4]
  wire  _T_1437; // @[MemPrimitives.scala 126:35:@33958.4]
  wire  _T_1438; // @[MemPrimitives.scala 126:35:@33959.4]
  wire [10:0] _T_1440; // @[Cat.scala 30:58:@33961.4]
  wire [10:0] _T_1442; // @[Cat.scala 30:58:@33963.4]
  wire [10:0] _T_1444; // @[Cat.scala 30:58:@33965.4]
  wire [10:0] _T_1446; // @[Cat.scala 30:58:@33967.4]
  wire [10:0] _T_1448; // @[Cat.scala 30:58:@33969.4]
  wire [10:0] _T_1450; // @[Cat.scala 30:58:@33971.4]
  wire [10:0] _T_1451; // @[Mux.scala 31:69:@33972.4]
  wire [10:0] _T_1452; // @[Mux.scala 31:69:@33973.4]
  wire [10:0] _T_1453; // @[Mux.scala 31:69:@33974.4]
  wire [10:0] _T_1454; // @[Mux.scala 31:69:@33975.4]
  wire [10:0] _T_1455; // @[Mux.scala 31:69:@33976.4]
  wire  _T_1463; // @[MemPrimitives.scala 110:228:@33985.4]
  wire  _T_1469; // @[MemPrimitives.scala 110:228:@33989.4]
  wire  _T_1475; // @[MemPrimitives.scala 110:228:@33993.4]
  wire  _T_1481; // @[MemPrimitives.scala 110:228:@33997.4]
  wire  _T_1483; // @[MemPrimitives.scala 126:35:@34006.4]
  wire  _T_1484; // @[MemPrimitives.scala 126:35:@34007.4]
  wire  _T_1485; // @[MemPrimitives.scala 126:35:@34008.4]
  wire  _T_1486; // @[MemPrimitives.scala 126:35:@34009.4]
  wire [10:0] _T_1488; // @[Cat.scala 30:58:@34011.4]
  wire [10:0] _T_1490; // @[Cat.scala 30:58:@34013.4]
  wire [10:0] _T_1492; // @[Cat.scala 30:58:@34015.4]
  wire [10:0] _T_1494; // @[Cat.scala 30:58:@34017.4]
  wire [10:0] _T_1495; // @[Mux.scala 31:69:@34018.4]
  wire [10:0] _T_1496; // @[Mux.scala 31:69:@34019.4]
  wire [10:0] _T_1497; // @[Mux.scala 31:69:@34020.4]
  wire  _T_1505; // @[MemPrimitives.scala 110:228:@34029.4]
  wire  _T_1511; // @[MemPrimitives.scala 110:228:@34033.4]
  wire  _T_1517; // @[MemPrimitives.scala 110:228:@34037.4]
  wire  _T_1523; // @[MemPrimitives.scala 110:228:@34041.4]
  wire  _T_1529; // @[MemPrimitives.scala 110:228:@34045.4]
  wire  _T_1535; // @[MemPrimitives.scala 110:228:@34049.4]
  wire  _T_1537; // @[MemPrimitives.scala 126:35:@34060.4]
  wire  _T_1538; // @[MemPrimitives.scala 126:35:@34061.4]
  wire  _T_1539; // @[MemPrimitives.scala 126:35:@34062.4]
  wire  _T_1540; // @[MemPrimitives.scala 126:35:@34063.4]
  wire  _T_1541; // @[MemPrimitives.scala 126:35:@34064.4]
  wire  _T_1542; // @[MemPrimitives.scala 126:35:@34065.4]
  wire [10:0] _T_1544; // @[Cat.scala 30:58:@34067.4]
  wire [10:0] _T_1546; // @[Cat.scala 30:58:@34069.4]
  wire [10:0] _T_1548; // @[Cat.scala 30:58:@34071.4]
  wire [10:0] _T_1550; // @[Cat.scala 30:58:@34073.4]
  wire [10:0] _T_1552; // @[Cat.scala 30:58:@34075.4]
  wire [10:0] _T_1554; // @[Cat.scala 30:58:@34077.4]
  wire [10:0] _T_1555; // @[Mux.scala 31:69:@34078.4]
  wire [10:0] _T_1556; // @[Mux.scala 31:69:@34079.4]
  wire [10:0] _T_1557; // @[Mux.scala 31:69:@34080.4]
  wire [10:0] _T_1558; // @[Mux.scala 31:69:@34081.4]
  wire [10:0] _T_1559; // @[Mux.scala 31:69:@34082.4]
  wire  _T_1564; // @[MemPrimitives.scala 110:210:@34089.4]
  wire  _T_1567; // @[MemPrimitives.scala 110:228:@34091.4]
  wire  _T_1570; // @[MemPrimitives.scala 110:210:@34093.4]
  wire  _T_1573; // @[MemPrimitives.scala 110:228:@34095.4]
  wire  _T_1576; // @[MemPrimitives.scala 110:210:@34097.4]
  wire  _T_1579; // @[MemPrimitives.scala 110:228:@34099.4]
  wire  _T_1582; // @[MemPrimitives.scala 110:210:@34101.4]
  wire  _T_1585; // @[MemPrimitives.scala 110:228:@34103.4]
  wire  _T_1587; // @[MemPrimitives.scala 126:35:@34112.4]
  wire  _T_1588; // @[MemPrimitives.scala 126:35:@34113.4]
  wire  _T_1589; // @[MemPrimitives.scala 126:35:@34114.4]
  wire  _T_1590; // @[MemPrimitives.scala 126:35:@34115.4]
  wire [10:0] _T_1592; // @[Cat.scala 30:58:@34117.4]
  wire [10:0] _T_1594; // @[Cat.scala 30:58:@34119.4]
  wire [10:0] _T_1596; // @[Cat.scala 30:58:@34121.4]
  wire [10:0] _T_1598; // @[Cat.scala 30:58:@34123.4]
  wire [10:0] _T_1599; // @[Mux.scala 31:69:@34124.4]
  wire [10:0] _T_1600; // @[Mux.scala 31:69:@34125.4]
  wire [10:0] _T_1601; // @[Mux.scala 31:69:@34126.4]
  wire  _T_1606; // @[MemPrimitives.scala 110:210:@34133.4]
  wire  _T_1609; // @[MemPrimitives.scala 110:228:@34135.4]
  wire  _T_1612; // @[MemPrimitives.scala 110:210:@34137.4]
  wire  _T_1615; // @[MemPrimitives.scala 110:228:@34139.4]
  wire  _T_1618; // @[MemPrimitives.scala 110:210:@34141.4]
  wire  _T_1621; // @[MemPrimitives.scala 110:228:@34143.4]
  wire  _T_1624; // @[MemPrimitives.scala 110:210:@34145.4]
  wire  _T_1627; // @[MemPrimitives.scala 110:228:@34147.4]
  wire  _T_1630; // @[MemPrimitives.scala 110:210:@34149.4]
  wire  _T_1633; // @[MemPrimitives.scala 110:228:@34151.4]
  wire  _T_1636; // @[MemPrimitives.scala 110:210:@34153.4]
  wire  _T_1639; // @[MemPrimitives.scala 110:228:@34155.4]
  wire  _T_1641; // @[MemPrimitives.scala 126:35:@34166.4]
  wire  _T_1642; // @[MemPrimitives.scala 126:35:@34167.4]
  wire  _T_1643; // @[MemPrimitives.scala 126:35:@34168.4]
  wire  _T_1644; // @[MemPrimitives.scala 126:35:@34169.4]
  wire  _T_1645; // @[MemPrimitives.scala 126:35:@34170.4]
  wire  _T_1646; // @[MemPrimitives.scala 126:35:@34171.4]
  wire [10:0] _T_1648; // @[Cat.scala 30:58:@34173.4]
  wire [10:0] _T_1650; // @[Cat.scala 30:58:@34175.4]
  wire [10:0] _T_1652; // @[Cat.scala 30:58:@34177.4]
  wire [10:0] _T_1654; // @[Cat.scala 30:58:@34179.4]
  wire [10:0] _T_1656; // @[Cat.scala 30:58:@34181.4]
  wire [10:0] _T_1658; // @[Cat.scala 30:58:@34183.4]
  wire [10:0] _T_1659; // @[Mux.scala 31:69:@34184.4]
  wire [10:0] _T_1660; // @[Mux.scala 31:69:@34185.4]
  wire [10:0] _T_1661; // @[Mux.scala 31:69:@34186.4]
  wire [10:0] _T_1662; // @[Mux.scala 31:69:@34187.4]
  wire [10:0] _T_1663; // @[Mux.scala 31:69:@34188.4]
  wire  _T_1671; // @[MemPrimitives.scala 110:228:@34197.4]
  wire  _T_1677; // @[MemPrimitives.scala 110:228:@34201.4]
  wire  _T_1683; // @[MemPrimitives.scala 110:228:@34205.4]
  wire  _T_1689; // @[MemPrimitives.scala 110:228:@34209.4]
  wire  _T_1691; // @[MemPrimitives.scala 126:35:@34218.4]
  wire  _T_1692; // @[MemPrimitives.scala 126:35:@34219.4]
  wire  _T_1693; // @[MemPrimitives.scala 126:35:@34220.4]
  wire  _T_1694; // @[MemPrimitives.scala 126:35:@34221.4]
  wire [10:0] _T_1696; // @[Cat.scala 30:58:@34223.4]
  wire [10:0] _T_1698; // @[Cat.scala 30:58:@34225.4]
  wire [10:0] _T_1700; // @[Cat.scala 30:58:@34227.4]
  wire [10:0] _T_1702; // @[Cat.scala 30:58:@34229.4]
  wire [10:0] _T_1703; // @[Mux.scala 31:69:@34230.4]
  wire [10:0] _T_1704; // @[Mux.scala 31:69:@34231.4]
  wire [10:0] _T_1705; // @[Mux.scala 31:69:@34232.4]
  wire  _T_1713; // @[MemPrimitives.scala 110:228:@34241.4]
  wire  _T_1719; // @[MemPrimitives.scala 110:228:@34245.4]
  wire  _T_1725; // @[MemPrimitives.scala 110:228:@34249.4]
  wire  _T_1731; // @[MemPrimitives.scala 110:228:@34253.4]
  wire  _T_1737; // @[MemPrimitives.scala 110:228:@34257.4]
  wire  _T_1743; // @[MemPrimitives.scala 110:228:@34261.4]
  wire  _T_1745; // @[MemPrimitives.scala 126:35:@34272.4]
  wire  _T_1746; // @[MemPrimitives.scala 126:35:@34273.4]
  wire  _T_1747; // @[MemPrimitives.scala 126:35:@34274.4]
  wire  _T_1748; // @[MemPrimitives.scala 126:35:@34275.4]
  wire  _T_1749; // @[MemPrimitives.scala 126:35:@34276.4]
  wire  _T_1750; // @[MemPrimitives.scala 126:35:@34277.4]
  wire [10:0] _T_1752; // @[Cat.scala 30:58:@34279.4]
  wire [10:0] _T_1754; // @[Cat.scala 30:58:@34281.4]
  wire [10:0] _T_1756; // @[Cat.scala 30:58:@34283.4]
  wire [10:0] _T_1758; // @[Cat.scala 30:58:@34285.4]
  wire [10:0] _T_1760; // @[Cat.scala 30:58:@34287.4]
  wire [10:0] _T_1762; // @[Cat.scala 30:58:@34289.4]
  wire [10:0] _T_1763; // @[Mux.scala 31:69:@34290.4]
  wire [10:0] _T_1764; // @[Mux.scala 31:69:@34291.4]
  wire [10:0] _T_1765; // @[Mux.scala 31:69:@34292.4]
  wire [10:0] _T_1766; // @[Mux.scala 31:69:@34293.4]
  wire [10:0] _T_1767; // @[Mux.scala 31:69:@34294.4]
  wire  _T_1775; // @[MemPrimitives.scala 110:228:@34303.4]
  wire  _T_1781; // @[MemPrimitives.scala 110:228:@34307.4]
  wire  _T_1787; // @[MemPrimitives.scala 110:228:@34311.4]
  wire  _T_1793; // @[MemPrimitives.scala 110:228:@34315.4]
  wire  _T_1795; // @[MemPrimitives.scala 126:35:@34324.4]
  wire  _T_1796; // @[MemPrimitives.scala 126:35:@34325.4]
  wire  _T_1797; // @[MemPrimitives.scala 126:35:@34326.4]
  wire  _T_1798; // @[MemPrimitives.scala 126:35:@34327.4]
  wire [10:0] _T_1800; // @[Cat.scala 30:58:@34329.4]
  wire [10:0] _T_1802; // @[Cat.scala 30:58:@34331.4]
  wire [10:0] _T_1804; // @[Cat.scala 30:58:@34333.4]
  wire [10:0] _T_1806; // @[Cat.scala 30:58:@34335.4]
  wire [10:0] _T_1807; // @[Mux.scala 31:69:@34336.4]
  wire [10:0] _T_1808; // @[Mux.scala 31:69:@34337.4]
  wire [10:0] _T_1809; // @[Mux.scala 31:69:@34338.4]
  wire  _T_1817; // @[MemPrimitives.scala 110:228:@34347.4]
  wire  _T_1823; // @[MemPrimitives.scala 110:228:@34351.4]
  wire  _T_1829; // @[MemPrimitives.scala 110:228:@34355.4]
  wire  _T_1835; // @[MemPrimitives.scala 110:228:@34359.4]
  wire  _T_1841; // @[MemPrimitives.scala 110:228:@34363.4]
  wire  _T_1847; // @[MemPrimitives.scala 110:228:@34367.4]
  wire  _T_1849; // @[MemPrimitives.scala 126:35:@34378.4]
  wire  _T_1850; // @[MemPrimitives.scala 126:35:@34379.4]
  wire  _T_1851; // @[MemPrimitives.scala 126:35:@34380.4]
  wire  _T_1852; // @[MemPrimitives.scala 126:35:@34381.4]
  wire  _T_1853; // @[MemPrimitives.scala 126:35:@34382.4]
  wire  _T_1854; // @[MemPrimitives.scala 126:35:@34383.4]
  wire [10:0] _T_1856; // @[Cat.scala 30:58:@34385.4]
  wire [10:0] _T_1858; // @[Cat.scala 30:58:@34387.4]
  wire [10:0] _T_1860; // @[Cat.scala 30:58:@34389.4]
  wire [10:0] _T_1862; // @[Cat.scala 30:58:@34391.4]
  wire [10:0] _T_1864; // @[Cat.scala 30:58:@34393.4]
  wire [10:0] _T_1866; // @[Cat.scala 30:58:@34395.4]
  wire [10:0] _T_1867; // @[Mux.scala 31:69:@34396.4]
  wire [10:0] _T_1868; // @[Mux.scala 31:69:@34397.4]
  wire [10:0] _T_1869; // @[Mux.scala 31:69:@34398.4]
  wire [10:0] _T_1870; // @[Mux.scala 31:69:@34399.4]
  wire [10:0] _T_1871; // @[Mux.scala 31:69:@34400.4]
  wire  _T_1876; // @[MemPrimitives.scala 110:210:@34407.4]
  wire  _T_1879; // @[MemPrimitives.scala 110:228:@34409.4]
  wire  _T_1882; // @[MemPrimitives.scala 110:210:@34411.4]
  wire  _T_1885; // @[MemPrimitives.scala 110:228:@34413.4]
  wire  _T_1888; // @[MemPrimitives.scala 110:210:@34415.4]
  wire  _T_1891; // @[MemPrimitives.scala 110:228:@34417.4]
  wire  _T_1894; // @[MemPrimitives.scala 110:210:@34419.4]
  wire  _T_1897; // @[MemPrimitives.scala 110:228:@34421.4]
  wire  _T_1899; // @[MemPrimitives.scala 126:35:@34430.4]
  wire  _T_1900; // @[MemPrimitives.scala 126:35:@34431.4]
  wire  _T_1901; // @[MemPrimitives.scala 126:35:@34432.4]
  wire  _T_1902; // @[MemPrimitives.scala 126:35:@34433.4]
  wire [10:0] _T_1904; // @[Cat.scala 30:58:@34435.4]
  wire [10:0] _T_1906; // @[Cat.scala 30:58:@34437.4]
  wire [10:0] _T_1908; // @[Cat.scala 30:58:@34439.4]
  wire [10:0] _T_1910; // @[Cat.scala 30:58:@34441.4]
  wire [10:0] _T_1911; // @[Mux.scala 31:69:@34442.4]
  wire [10:0] _T_1912; // @[Mux.scala 31:69:@34443.4]
  wire [10:0] _T_1913; // @[Mux.scala 31:69:@34444.4]
  wire  _T_1918; // @[MemPrimitives.scala 110:210:@34451.4]
  wire  _T_1921; // @[MemPrimitives.scala 110:228:@34453.4]
  wire  _T_1924; // @[MemPrimitives.scala 110:210:@34455.4]
  wire  _T_1927; // @[MemPrimitives.scala 110:228:@34457.4]
  wire  _T_1930; // @[MemPrimitives.scala 110:210:@34459.4]
  wire  _T_1933; // @[MemPrimitives.scala 110:228:@34461.4]
  wire  _T_1936; // @[MemPrimitives.scala 110:210:@34463.4]
  wire  _T_1939; // @[MemPrimitives.scala 110:228:@34465.4]
  wire  _T_1942; // @[MemPrimitives.scala 110:210:@34467.4]
  wire  _T_1945; // @[MemPrimitives.scala 110:228:@34469.4]
  wire  _T_1948; // @[MemPrimitives.scala 110:210:@34471.4]
  wire  _T_1951; // @[MemPrimitives.scala 110:228:@34473.4]
  wire  _T_1953; // @[MemPrimitives.scala 126:35:@34484.4]
  wire  _T_1954; // @[MemPrimitives.scala 126:35:@34485.4]
  wire  _T_1955; // @[MemPrimitives.scala 126:35:@34486.4]
  wire  _T_1956; // @[MemPrimitives.scala 126:35:@34487.4]
  wire  _T_1957; // @[MemPrimitives.scala 126:35:@34488.4]
  wire  _T_1958; // @[MemPrimitives.scala 126:35:@34489.4]
  wire [10:0] _T_1960; // @[Cat.scala 30:58:@34491.4]
  wire [10:0] _T_1962; // @[Cat.scala 30:58:@34493.4]
  wire [10:0] _T_1964; // @[Cat.scala 30:58:@34495.4]
  wire [10:0] _T_1966; // @[Cat.scala 30:58:@34497.4]
  wire [10:0] _T_1968; // @[Cat.scala 30:58:@34499.4]
  wire [10:0] _T_1970; // @[Cat.scala 30:58:@34501.4]
  wire [10:0] _T_1971; // @[Mux.scala 31:69:@34502.4]
  wire [10:0] _T_1972; // @[Mux.scala 31:69:@34503.4]
  wire [10:0] _T_1973; // @[Mux.scala 31:69:@34504.4]
  wire [10:0] _T_1974; // @[Mux.scala 31:69:@34505.4]
  wire [10:0] _T_1975; // @[Mux.scala 31:69:@34506.4]
  wire  _T_1983; // @[MemPrimitives.scala 110:228:@34515.4]
  wire  _T_1989; // @[MemPrimitives.scala 110:228:@34519.4]
  wire  _T_1995; // @[MemPrimitives.scala 110:228:@34523.4]
  wire  _T_2001; // @[MemPrimitives.scala 110:228:@34527.4]
  wire  _T_2003; // @[MemPrimitives.scala 126:35:@34536.4]
  wire  _T_2004; // @[MemPrimitives.scala 126:35:@34537.4]
  wire  _T_2005; // @[MemPrimitives.scala 126:35:@34538.4]
  wire  _T_2006; // @[MemPrimitives.scala 126:35:@34539.4]
  wire [10:0] _T_2008; // @[Cat.scala 30:58:@34541.4]
  wire [10:0] _T_2010; // @[Cat.scala 30:58:@34543.4]
  wire [10:0] _T_2012; // @[Cat.scala 30:58:@34545.4]
  wire [10:0] _T_2014; // @[Cat.scala 30:58:@34547.4]
  wire [10:0] _T_2015; // @[Mux.scala 31:69:@34548.4]
  wire [10:0] _T_2016; // @[Mux.scala 31:69:@34549.4]
  wire [10:0] _T_2017; // @[Mux.scala 31:69:@34550.4]
  wire  _T_2025; // @[MemPrimitives.scala 110:228:@34559.4]
  wire  _T_2031; // @[MemPrimitives.scala 110:228:@34563.4]
  wire  _T_2037; // @[MemPrimitives.scala 110:228:@34567.4]
  wire  _T_2043; // @[MemPrimitives.scala 110:228:@34571.4]
  wire  _T_2049; // @[MemPrimitives.scala 110:228:@34575.4]
  wire  _T_2055; // @[MemPrimitives.scala 110:228:@34579.4]
  wire  _T_2057; // @[MemPrimitives.scala 126:35:@34590.4]
  wire  _T_2058; // @[MemPrimitives.scala 126:35:@34591.4]
  wire  _T_2059; // @[MemPrimitives.scala 126:35:@34592.4]
  wire  _T_2060; // @[MemPrimitives.scala 126:35:@34593.4]
  wire  _T_2061; // @[MemPrimitives.scala 126:35:@34594.4]
  wire  _T_2062; // @[MemPrimitives.scala 126:35:@34595.4]
  wire [10:0] _T_2064; // @[Cat.scala 30:58:@34597.4]
  wire [10:0] _T_2066; // @[Cat.scala 30:58:@34599.4]
  wire [10:0] _T_2068; // @[Cat.scala 30:58:@34601.4]
  wire [10:0] _T_2070; // @[Cat.scala 30:58:@34603.4]
  wire [10:0] _T_2072; // @[Cat.scala 30:58:@34605.4]
  wire [10:0] _T_2074; // @[Cat.scala 30:58:@34607.4]
  wire [10:0] _T_2075; // @[Mux.scala 31:69:@34608.4]
  wire [10:0] _T_2076; // @[Mux.scala 31:69:@34609.4]
  wire [10:0] _T_2077; // @[Mux.scala 31:69:@34610.4]
  wire [10:0] _T_2078; // @[Mux.scala 31:69:@34611.4]
  wire [10:0] _T_2079; // @[Mux.scala 31:69:@34612.4]
  wire  _T_2087; // @[MemPrimitives.scala 110:228:@34621.4]
  wire  _T_2093; // @[MemPrimitives.scala 110:228:@34625.4]
  wire  _T_2099; // @[MemPrimitives.scala 110:228:@34629.4]
  wire  _T_2105; // @[MemPrimitives.scala 110:228:@34633.4]
  wire  _T_2107; // @[MemPrimitives.scala 126:35:@34642.4]
  wire  _T_2108; // @[MemPrimitives.scala 126:35:@34643.4]
  wire  _T_2109; // @[MemPrimitives.scala 126:35:@34644.4]
  wire  _T_2110; // @[MemPrimitives.scala 126:35:@34645.4]
  wire [10:0] _T_2112; // @[Cat.scala 30:58:@34647.4]
  wire [10:0] _T_2114; // @[Cat.scala 30:58:@34649.4]
  wire [10:0] _T_2116; // @[Cat.scala 30:58:@34651.4]
  wire [10:0] _T_2118; // @[Cat.scala 30:58:@34653.4]
  wire [10:0] _T_2119; // @[Mux.scala 31:69:@34654.4]
  wire [10:0] _T_2120; // @[Mux.scala 31:69:@34655.4]
  wire [10:0] _T_2121; // @[Mux.scala 31:69:@34656.4]
  wire  _T_2129; // @[MemPrimitives.scala 110:228:@34665.4]
  wire  _T_2135; // @[MemPrimitives.scala 110:228:@34669.4]
  wire  _T_2141; // @[MemPrimitives.scala 110:228:@34673.4]
  wire  _T_2147; // @[MemPrimitives.scala 110:228:@34677.4]
  wire  _T_2153; // @[MemPrimitives.scala 110:228:@34681.4]
  wire  _T_2159; // @[MemPrimitives.scala 110:228:@34685.4]
  wire  _T_2161; // @[MemPrimitives.scala 126:35:@34696.4]
  wire  _T_2162; // @[MemPrimitives.scala 126:35:@34697.4]
  wire  _T_2163; // @[MemPrimitives.scala 126:35:@34698.4]
  wire  _T_2164; // @[MemPrimitives.scala 126:35:@34699.4]
  wire  _T_2165; // @[MemPrimitives.scala 126:35:@34700.4]
  wire  _T_2166; // @[MemPrimitives.scala 126:35:@34701.4]
  wire [10:0] _T_2168; // @[Cat.scala 30:58:@34703.4]
  wire [10:0] _T_2170; // @[Cat.scala 30:58:@34705.4]
  wire [10:0] _T_2172; // @[Cat.scala 30:58:@34707.4]
  wire [10:0] _T_2174; // @[Cat.scala 30:58:@34709.4]
  wire [10:0] _T_2176; // @[Cat.scala 30:58:@34711.4]
  wire [10:0] _T_2178; // @[Cat.scala 30:58:@34713.4]
  wire [10:0] _T_2179; // @[Mux.scala 31:69:@34714.4]
  wire [10:0] _T_2180; // @[Mux.scala 31:69:@34715.4]
  wire [10:0] _T_2181; // @[Mux.scala 31:69:@34716.4]
  wire [10:0] _T_2182; // @[Mux.scala 31:69:@34717.4]
  wire [10:0] _T_2183; // @[Mux.scala 31:69:@34718.4]
  wire  _T_2279; // @[package.scala 96:25:@34847.4 package.scala 96:25:@34848.4]
  wire [31:0] _T_2283; // @[Mux.scala 31:69:@34857.4]
  wire  _T_2276; // @[package.scala 96:25:@34839.4 package.scala 96:25:@34840.4]
  wire [31:0] _T_2284; // @[Mux.scala 31:69:@34858.4]
  wire  _T_2273; // @[package.scala 96:25:@34831.4 package.scala 96:25:@34832.4]
  wire [31:0] _T_2285; // @[Mux.scala 31:69:@34859.4]
  wire  _T_2270; // @[package.scala 96:25:@34823.4 package.scala 96:25:@34824.4]
  wire [31:0] _T_2286; // @[Mux.scala 31:69:@34860.4]
  wire  _T_2267; // @[package.scala 96:25:@34815.4 package.scala 96:25:@34816.4]
  wire [31:0] _T_2287; // @[Mux.scala 31:69:@34861.4]
  wire  _T_2264; // @[package.scala 96:25:@34807.4 package.scala 96:25:@34808.4]
  wire [31:0] _T_2288; // @[Mux.scala 31:69:@34862.4]
  wire  _T_2261; // @[package.scala 96:25:@34799.4 package.scala 96:25:@34800.4]
  wire [31:0] _T_2289; // @[Mux.scala 31:69:@34863.4]
  wire  _T_2258; // @[package.scala 96:25:@34791.4 package.scala 96:25:@34792.4]
  wire [31:0] _T_2290; // @[Mux.scala 31:69:@34864.4]
  wire  _T_2255; // @[package.scala 96:25:@34783.4 package.scala 96:25:@34784.4]
  wire [31:0] _T_2291; // @[Mux.scala 31:69:@34865.4]
  wire  _T_2252; // @[package.scala 96:25:@34775.4 package.scala 96:25:@34776.4]
  wire [31:0] _T_2292; // @[Mux.scala 31:69:@34866.4]
  wire  _T_2249; // @[package.scala 96:25:@34767.4 package.scala 96:25:@34768.4]
  wire  _T_2386; // @[package.scala 96:25:@34991.4 package.scala 96:25:@34992.4]
  wire [31:0] _T_2390; // @[Mux.scala 31:69:@35001.4]
  wire  _T_2383; // @[package.scala 96:25:@34983.4 package.scala 96:25:@34984.4]
  wire [31:0] _T_2391; // @[Mux.scala 31:69:@35002.4]
  wire  _T_2380; // @[package.scala 96:25:@34975.4 package.scala 96:25:@34976.4]
  wire [31:0] _T_2392; // @[Mux.scala 31:69:@35003.4]
  wire  _T_2377; // @[package.scala 96:25:@34967.4 package.scala 96:25:@34968.4]
  wire [31:0] _T_2393; // @[Mux.scala 31:69:@35004.4]
  wire  _T_2374; // @[package.scala 96:25:@34959.4 package.scala 96:25:@34960.4]
  wire [31:0] _T_2394; // @[Mux.scala 31:69:@35005.4]
  wire  _T_2371; // @[package.scala 96:25:@34951.4 package.scala 96:25:@34952.4]
  wire [31:0] _T_2395; // @[Mux.scala 31:69:@35006.4]
  wire  _T_2368; // @[package.scala 96:25:@34943.4 package.scala 96:25:@34944.4]
  wire [31:0] _T_2396; // @[Mux.scala 31:69:@35007.4]
  wire  _T_2365; // @[package.scala 96:25:@34935.4 package.scala 96:25:@34936.4]
  wire [31:0] _T_2397; // @[Mux.scala 31:69:@35008.4]
  wire  _T_2362; // @[package.scala 96:25:@34927.4 package.scala 96:25:@34928.4]
  wire [31:0] _T_2398; // @[Mux.scala 31:69:@35009.4]
  wire  _T_2359; // @[package.scala 96:25:@34919.4 package.scala 96:25:@34920.4]
  wire [31:0] _T_2399; // @[Mux.scala 31:69:@35010.4]
  wire  _T_2356; // @[package.scala 96:25:@34911.4 package.scala 96:25:@34912.4]
  wire  _T_2493; // @[package.scala 96:25:@35135.4 package.scala 96:25:@35136.4]
  wire [31:0] _T_2497; // @[Mux.scala 31:69:@35145.4]
  wire  _T_2490; // @[package.scala 96:25:@35127.4 package.scala 96:25:@35128.4]
  wire [31:0] _T_2498; // @[Mux.scala 31:69:@35146.4]
  wire  _T_2487; // @[package.scala 96:25:@35119.4 package.scala 96:25:@35120.4]
  wire [31:0] _T_2499; // @[Mux.scala 31:69:@35147.4]
  wire  _T_2484; // @[package.scala 96:25:@35111.4 package.scala 96:25:@35112.4]
  wire [31:0] _T_2500; // @[Mux.scala 31:69:@35148.4]
  wire  _T_2481; // @[package.scala 96:25:@35103.4 package.scala 96:25:@35104.4]
  wire [31:0] _T_2501; // @[Mux.scala 31:69:@35149.4]
  wire  _T_2478; // @[package.scala 96:25:@35095.4 package.scala 96:25:@35096.4]
  wire [31:0] _T_2502; // @[Mux.scala 31:69:@35150.4]
  wire  _T_2475; // @[package.scala 96:25:@35087.4 package.scala 96:25:@35088.4]
  wire [31:0] _T_2503; // @[Mux.scala 31:69:@35151.4]
  wire  _T_2472; // @[package.scala 96:25:@35079.4 package.scala 96:25:@35080.4]
  wire [31:0] _T_2504; // @[Mux.scala 31:69:@35152.4]
  wire  _T_2469; // @[package.scala 96:25:@35071.4 package.scala 96:25:@35072.4]
  wire [31:0] _T_2505; // @[Mux.scala 31:69:@35153.4]
  wire  _T_2466; // @[package.scala 96:25:@35063.4 package.scala 96:25:@35064.4]
  wire [31:0] _T_2506; // @[Mux.scala 31:69:@35154.4]
  wire  _T_2463; // @[package.scala 96:25:@35055.4 package.scala 96:25:@35056.4]
  wire  _T_2600; // @[package.scala 96:25:@35279.4 package.scala 96:25:@35280.4]
  wire [31:0] _T_2604; // @[Mux.scala 31:69:@35289.4]
  wire  _T_2597; // @[package.scala 96:25:@35271.4 package.scala 96:25:@35272.4]
  wire [31:0] _T_2605; // @[Mux.scala 31:69:@35290.4]
  wire  _T_2594; // @[package.scala 96:25:@35263.4 package.scala 96:25:@35264.4]
  wire [31:0] _T_2606; // @[Mux.scala 31:69:@35291.4]
  wire  _T_2591; // @[package.scala 96:25:@35255.4 package.scala 96:25:@35256.4]
  wire [31:0] _T_2607; // @[Mux.scala 31:69:@35292.4]
  wire  _T_2588; // @[package.scala 96:25:@35247.4 package.scala 96:25:@35248.4]
  wire [31:0] _T_2608; // @[Mux.scala 31:69:@35293.4]
  wire  _T_2585; // @[package.scala 96:25:@35239.4 package.scala 96:25:@35240.4]
  wire [31:0] _T_2609; // @[Mux.scala 31:69:@35294.4]
  wire  _T_2582; // @[package.scala 96:25:@35231.4 package.scala 96:25:@35232.4]
  wire [31:0] _T_2610; // @[Mux.scala 31:69:@35295.4]
  wire  _T_2579; // @[package.scala 96:25:@35223.4 package.scala 96:25:@35224.4]
  wire [31:0] _T_2611; // @[Mux.scala 31:69:@35296.4]
  wire  _T_2576; // @[package.scala 96:25:@35215.4 package.scala 96:25:@35216.4]
  wire [31:0] _T_2612; // @[Mux.scala 31:69:@35297.4]
  wire  _T_2573; // @[package.scala 96:25:@35207.4 package.scala 96:25:@35208.4]
  wire [31:0] _T_2613; // @[Mux.scala 31:69:@35298.4]
  wire  _T_2570; // @[package.scala 96:25:@35199.4 package.scala 96:25:@35200.4]
  wire  _T_2707; // @[package.scala 96:25:@35423.4 package.scala 96:25:@35424.4]
  wire [31:0] _T_2711; // @[Mux.scala 31:69:@35433.4]
  wire  _T_2704; // @[package.scala 96:25:@35415.4 package.scala 96:25:@35416.4]
  wire [31:0] _T_2712; // @[Mux.scala 31:69:@35434.4]
  wire  _T_2701; // @[package.scala 96:25:@35407.4 package.scala 96:25:@35408.4]
  wire [31:0] _T_2713; // @[Mux.scala 31:69:@35435.4]
  wire  _T_2698; // @[package.scala 96:25:@35399.4 package.scala 96:25:@35400.4]
  wire [31:0] _T_2714; // @[Mux.scala 31:69:@35436.4]
  wire  _T_2695; // @[package.scala 96:25:@35391.4 package.scala 96:25:@35392.4]
  wire [31:0] _T_2715; // @[Mux.scala 31:69:@35437.4]
  wire  _T_2692; // @[package.scala 96:25:@35383.4 package.scala 96:25:@35384.4]
  wire [31:0] _T_2716; // @[Mux.scala 31:69:@35438.4]
  wire  _T_2689; // @[package.scala 96:25:@35375.4 package.scala 96:25:@35376.4]
  wire [31:0] _T_2717; // @[Mux.scala 31:69:@35439.4]
  wire  _T_2686; // @[package.scala 96:25:@35367.4 package.scala 96:25:@35368.4]
  wire [31:0] _T_2718; // @[Mux.scala 31:69:@35440.4]
  wire  _T_2683; // @[package.scala 96:25:@35359.4 package.scala 96:25:@35360.4]
  wire [31:0] _T_2719; // @[Mux.scala 31:69:@35441.4]
  wire  _T_2680; // @[package.scala 96:25:@35351.4 package.scala 96:25:@35352.4]
  wire [31:0] _T_2720; // @[Mux.scala 31:69:@35442.4]
  wire  _T_2677; // @[package.scala 96:25:@35343.4 package.scala 96:25:@35344.4]
  wire  _T_2814; // @[package.scala 96:25:@35567.4 package.scala 96:25:@35568.4]
  wire [31:0] _T_2818; // @[Mux.scala 31:69:@35577.4]
  wire  _T_2811; // @[package.scala 96:25:@35559.4 package.scala 96:25:@35560.4]
  wire [31:0] _T_2819; // @[Mux.scala 31:69:@35578.4]
  wire  _T_2808; // @[package.scala 96:25:@35551.4 package.scala 96:25:@35552.4]
  wire [31:0] _T_2820; // @[Mux.scala 31:69:@35579.4]
  wire  _T_2805; // @[package.scala 96:25:@35543.4 package.scala 96:25:@35544.4]
  wire [31:0] _T_2821; // @[Mux.scala 31:69:@35580.4]
  wire  _T_2802; // @[package.scala 96:25:@35535.4 package.scala 96:25:@35536.4]
  wire [31:0] _T_2822; // @[Mux.scala 31:69:@35581.4]
  wire  _T_2799; // @[package.scala 96:25:@35527.4 package.scala 96:25:@35528.4]
  wire [31:0] _T_2823; // @[Mux.scala 31:69:@35582.4]
  wire  _T_2796; // @[package.scala 96:25:@35519.4 package.scala 96:25:@35520.4]
  wire [31:0] _T_2824; // @[Mux.scala 31:69:@35583.4]
  wire  _T_2793; // @[package.scala 96:25:@35511.4 package.scala 96:25:@35512.4]
  wire [31:0] _T_2825; // @[Mux.scala 31:69:@35584.4]
  wire  _T_2790; // @[package.scala 96:25:@35503.4 package.scala 96:25:@35504.4]
  wire [31:0] _T_2826; // @[Mux.scala 31:69:@35585.4]
  wire  _T_2787; // @[package.scala 96:25:@35495.4 package.scala 96:25:@35496.4]
  wire [31:0] _T_2827; // @[Mux.scala 31:69:@35586.4]
  wire  _T_2784; // @[package.scala 96:25:@35487.4 package.scala 96:25:@35488.4]
  wire  _T_2921; // @[package.scala 96:25:@35711.4 package.scala 96:25:@35712.4]
  wire [31:0] _T_2925; // @[Mux.scala 31:69:@35721.4]
  wire  _T_2918; // @[package.scala 96:25:@35703.4 package.scala 96:25:@35704.4]
  wire [31:0] _T_2926; // @[Mux.scala 31:69:@35722.4]
  wire  _T_2915; // @[package.scala 96:25:@35695.4 package.scala 96:25:@35696.4]
  wire [31:0] _T_2927; // @[Mux.scala 31:69:@35723.4]
  wire  _T_2912; // @[package.scala 96:25:@35687.4 package.scala 96:25:@35688.4]
  wire [31:0] _T_2928; // @[Mux.scala 31:69:@35724.4]
  wire  _T_2909; // @[package.scala 96:25:@35679.4 package.scala 96:25:@35680.4]
  wire [31:0] _T_2929; // @[Mux.scala 31:69:@35725.4]
  wire  _T_2906; // @[package.scala 96:25:@35671.4 package.scala 96:25:@35672.4]
  wire [31:0] _T_2930; // @[Mux.scala 31:69:@35726.4]
  wire  _T_2903; // @[package.scala 96:25:@35663.4 package.scala 96:25:@35664.4]
  wire [31:0] _T_2931; // @[Mux.scala 31:69:@35727.4]
  wire  _T_2900; // @[package.scala 96:25:@35655.4 package.scala 96:25:@35656.4]
  wire [31:0] _T_2932; // @[Mux.scala 31:69:@35728.4]
  wire  _T_2897; // @[package.scala 96:25:@35647.4 package.scala 96:25:@35648.4]
  wire [31:0] _T_2933; // @[Mux.scala 31:69:@35729.4]
  wire  _T_2894; // @[package.scala 96:25:@35639.4 package.scala 96:25:@35640.4]
  wire [31:0] _T_2934; // @[Mux.scala 31:69:@35730.4]
  wire  _T_2891; // @[package.scala 96:25:@35631.4 package.scala 96:25:@35632.4]
  wire  _T_3028; // @[package.scala 96:25:@35855.4 package.scala 96:25:@35856.4]
  wire [31:0] _T_3032; // @[Mux.scala 31:69:@35865.4]
  wire  _T_3025; // @[package.scala 96:25:@35847.4 package.scala 96:25:@35848.4]
  wire [31:0] _T_3033; // @[Mux.scala 31:69:@35866.4]
  wire  _T_3022; // @[package.scala 96:25:@35839.4 package.scala 96:25:@35840.4]
  wire [31:0] _T_3034; // @[Mux.scala 31:69:@35867.4]
  wire  _T_3019; // @[package.scala 96:25:@35831.4 package.scala 96:25:@35832.4]
  wire [31:0] _T_3035; // @[Mux.scala 31:69:@35868.4]
  wire  _T_3016; // @[package.scala 96:25:@35823.4 package.scala 96:25:@35824.4]
  wire [31:0] _T_3036; // @[Mux.scala 31:69:@35869.4]
  wire  _T_3013; // @[package.scala 96:25:@35815.4 package.scala 96:25:@35816.4]
  wire [31:0] _T_3037; // @[Mux.scala 31:69:@35870.4]
  wire  _T_3010; // @[package.scala 96:25:@35807.4 package.scala 96:25:@35808.4]
  wire [31:0] _T_3038; // @[Mux.scala 31:69:@35871.4]
  wire  _T_3007; // @[package.scala 96:25:@35799.4 package.scala 96:25:@35800.4]
  wire [31:0] _T_3039; // @[Mux.scala 31:69:@35872.4]
  wire  _T_3004; // @[package.scala 96:25:@35791.4 package.scala 96:25:@35792.4]
  wire [31:0] _T_3040; // @[Mux.scala 31:69:@35873.4]
  wire  _T_3001; // @[package.scala 96:25:@35783.4 package.scala 96:25:@35784.4]
  wire [31:0] _T_3041; // @[Mux.scala 31:69:@35874.4]
  wire  _T_2998; // @[package.scala 96:25:@35775.4 package.scala 96:25:@35776.4]
  wire  _T_3135; // @[package.scala 96:25:@35999.4 package.scala 96:25:@36000.4]
  wire [31:0] _T_3139; // @[Mux.scala 31:69:@36009.4]
  wire  _T_3132; // @[package.scala 96:25:@35991.4 package.scala 96:25:@35992.4]
  wire [31:0] _T_3140; // @[Mux.scala 31:69:@36010.4]
  wire  _T_3129; // @[package.scala 96:25:@35983.4 package.scala 96:25:@35984.4]
  wire [31:0] _T_3141; // @[Mux.scala 31:69:@36011.4]
  wire  _T_3126; // @[package.scala 96:25:@35975.4 package.scala 96:25:@35976.4]
  wire [31:0] _T_3142; // @[Mux.scala 31:69:@36012.4]
  wire  _T_3123; // @[package.scala 96:25:@35967.4 package.scala 96:25:@35968.4]
  wire [31:0] _T_3143; // @[Mux.scala 31:69:@36013.4]
  wire  _T_3120; // @[package.scala 96:25:@35959.4 package.scala 96:25:@35960.4]
  wire [31:0] _T_3144; // @[Mux.scala 31:69:@36014.4]
  wire  _T_3117; // @[package.scala 96:25:@35951.4 package.scala 96:25:@35952.4]
  wire [31:0] _T_3145; // @[Mux.scala 31:69:@36015.4]
  wire  _T_3114; // @[package.scala 96:25:@35943.4 package.scala 96:25:@35944.4]
  wire [31:0] _T_3146; // @[Mux.scala 31:69:@36016.4]
  wire  _T_3111; // @[package.scala 96:25:@35935.4 package.scala 96:25:@35936.4]
  wire [31:0] _T_3147; // @[Mux.scala 31:69:@36017.4]
  wire  _T_3108; // @[package.scala 96:25:@35927.4 package.scala 96:25:@35928.4]
  wire [31:0] _T_3148; // @[Mux.scala 31:69:@36018.4]
  wire  _T_3105; // @[package.scala 96:25:@35919.4 package.scala 96:25:@35920.4]
  wire  _T_3242; // @[package.scala 96:25:@36143.4 package.scala 96:25:@36144.4]
  wire [31:0] _T_3246; // @[Mux.scala 31:69:@36153.4]
  wire  _T_3239; // @[package.scala 96:25:@36135.4 package.scala 96:25:@36136.4]
  wire [31:0] _T_3247; // @[Mux.scala 31:69:@36154.4]
  wire  _T_3236; // @[package.scala 96:25:@36127.4 package.scala 96:25:@36128.4]
  wire [31:0] _T_3248; // @[Mux.scala 31:69:@36155.4]
  wire  _T_3233; // @[package.scala 96:25:@36119.4 package.scala 96:25:@36120.4]
  wire [31:0] _T_3249; // @[Mux.scala 31:69:@36156.4]
  wire  _T_3230; // @[package.scala 96:25:@36111.4 package.scala 96:25:@36112.4]
  wire [31:0] _T_3250; // @[Mux.scala 31:69:@36157.4]
  wire  _T_3227; // @[package.scala 96:25:@36103.4 package.scala 96:25:@36104.4]
  wire [31:0] _T_3251; // @[Mux.scala 31:69:@36158.4]
  wire  _T_3224; // @[package.scala 96:25:@36095.4 package.scala 96:25:@36096.4]
  wire [31:0] _T_3252; // @[Mux.scala 31:69:@36159.4]
  wire  _T_3221; // @[package.scala 96:25:@36087.4 package.scala 96:25:@36088.4]
  wire [31:0] _T_3253; // @[Mux.scala 31:69:@36160.4]
  wire  _T_3218; // @[package.scala 96:25:@36079.4 package.scala 96:25:@36080.4]
  wire [31:0] _T_3254; // @[Mux.scala 31:69:@36161.4]
  wire  _T_3215; // @[package.scala 96:25:@36071.4 package.scala 96:25:@36072.4]
  wire [31:0] _T_3255; // @[Mux.scala 31:69:@36162.4]
  wire  _T_3212; // @[package.scala 96:25:@36063.4 package.scala 96:25:@36064.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@32613.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@32629.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@32645.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@32661.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@32677.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@32693.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@32709.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@32725.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@32741.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@32757.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@32773.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@32789.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@32805.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@32821.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@32837.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@32853.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  Mem1D_5 Mem1D_16 ( // @[MemPrimitives.scala 64:21:@32869.4]
    .clock(Mem1D_16_clock),
    .reset(Mem1D_16_reset),
    .io_r_ofs_0(Mem1D_16_io_r_ofs_0),
    .io_r_backpressure(Mem1D_16_io_r_backpressure),
    .io_w_ofs_0(Mem1D_16_io_w_ofs_0),
    .io_w_data_0(Mem1D_16_io_w_data_0),
    .io_w_en_0(Mem1D_16_io_w_en_0),
    .io_output(Mem1D_16_io_output)
  );
  Mem1D_5 Mem1D_17 ( // @[MemPrimitives.scala 64:21:@32885.4]
    .clock(Mem1D_17_clock),
    .reset(Mem1D_17_reset),
    .io_r_ofs_0(Mem1D_17_io_r_ofs_0),
    .io_r_backpressure(Mem1D_17_io_r_backpressure),
    .io_w_ofs_0(Mem1D_17_io_w_ofs_0),
    .io_w_data_0(Mem1D_17_io_w_data_0),
    .io_w_en_0(Mem1D_17_io_w_en_0),
    .io_output(Mem1D_17_io_output)
  );
  Mem1D_5 Mem1D_18 ( // @[MemPrimitives.scala 64:21:@32901.4]
    .clock(Mem1D_18_clock),
    .reset(Mem1D_18_reset),
    .io_r_ofs_0(Mem1D_18_io_r_ofs_0),
    .io_r_backpressure(Mem1D_18_io_r_backpressure),
    .io_w_ofs_0(Mem1D_18_io_w_ofs_0),
    .io_w_data_0(Mem1D_18_io_w_data_0),
    .io_w_en_0(Mem1D_18_io_w_en_0),
    .io_output(Mem1D_18_io_output)
  );
  Mem1D_5 Mem1D_19 ( // @[MemPrimitives.scala 64:21:@32917.4]
    .clock(Mem1D_19_clock),
    .reset(Mem1D_19_reset),
    .io_r_ofs_0(Mem1D_19_io_r_ofs_0),
    .io_r_backpressure(Mem1D_19_io_r_backpressure),
    .io_w_ofs_0(Mem1D_19_io_w_ofs_0),
    .io_w_data_0(Mem1D_19_io_w_data_0),
    .io_w_en_0(Mem1D_19_io_w_en_0),
    .io_output(Mem1D_19_io_output)
  );
  Mem1D_5 Mem1D_20 ( // @[MemPrimitives.scala 64:21:@32933.4]
    .clock(Mem1D_20_clock),
    .reset(Mem1D_20_reset),
    .io_r_ofs_0(Mem1D_20_io_r_ofs_0),
    .io_r_backpressure(Mem1D_20_io_r_backpressure),
    .io_w_ofs_0(Mem1D_20_io_w_ofs_0),
    .io_w_data_0(Mem1D_20_io_w_data_0),
    .io_w_en_0(Mem1D_20_io_w_en_0),
    .io_output(Mem1D_20_io_output)
  );
  Mem1D_5 Mem1D_21 ( // @[MemPrimitives.scala 64:21:@32949.4]
    .clock(Mem1D_21_clock),
    .reset(Mem1D_21_reset),
    .io_r_ofs_0(Mem1D_21_io_r_ofs_0),
    .io_r_backpressure(Mem1D_21_io_r_backpressure),
    .io_w_ofs_0(Mem1D_21_io_w_ofs_0),
    .io_w_data_0(Mem1D_21_io_w_data_0),
    .io_w_en_0(Mem1D_21_io_w_en_0),
    .io_output(Mem1D_21_io_output)
  );
  Mem1D_5 Mem1D_22 ( // @[MemPrimitives.scala 64:21:@32965.4]
    .clock(Mem1D_22_clock),
    .reset(Mem1D_22_reset),
    .io_r_ofs_0(Mem1D_22_io_r_ofs_0),
    .io_r_backpressure(Mem1D_22_io_r_backpressure),
    .io_w_ofs_0(Mem1D_22_io_w_ofs_0),
    .io_w_data_0(Mem1D_22_io_w_data_0),
    .io_w_en_0(Mem1D_22_io_w_en_0),
    .io_output(Mem1D_22_io_output)
  );
  Mem1D_5 Mem1D_23 ( // @[MemPrimitives.scala 64:21:@32981.4]
    .clock(Mem1D_23_clock),
    .reset(Mem1D_23_reset),
    .io_r_ofs_0(Mem1D_23_io_r_ofs_0),
    .io_r_backpressure(Mem1D_23_io_r_backpressure),
    .io_w_ofs_0(Mem1D_23_io_w_ofs_0),
    .io_w_data_0(Mem1D_23_io_w_data_0),
    .io_w_en_0(Mem1D_23_io_w_en_0),
    .io_output(Mem1D_23_io_output)
  );
  StickySelects_25 StickySelects ( // @[MemPrimitives.scala 124:33:@33469.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3)
  );
  StickySelects_26 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@33521.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects_25 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@33575.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3)
  );
  StickySelects_26 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@33627.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects_25 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@33681.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3)
  );
  StickySelects_26 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@33733.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects_25 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@33787.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3)
  );
  StickySelects_26 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@33839.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects_25 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@33893.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3)
  );
  StickySelects_26 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@33945.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects_25 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@33999.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3)
  );
  StickySelects_26 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@34051.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects_25 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@34105.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3)
  );
  StickySelects_26 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@34157.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects_25 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@34211.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3)
  );
  StickySelects_26 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@34263.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  StickySelects_25 StickySelects_16 ( // @[MemPrimitives.scala 124:33:@34317.4]
    .clock(StickySelects_16_clock),
    .reset(StickySelects_16_reset),
    .io_ins_0(StickySelects_16_io_ins_0),
    .io_ins_1(StickySelects_16_io_ins_1),
    .io_ins_2(StickySelects_16_io_ins_2),
    .io_ins_3(StickySelects_16_io_ins_3),
    .io_outs_0(StickySelects_16_io_outs_0),
    .io_outs_1(StickySelects_16_io_outs_1),
    .io_outs_2(StickySelects_16_io_outs_2),
    .io_outs_3(StickySelects_16_io_outs_3)
  );
  StickySelects_26 StickySelects_17 ( // @[MemPrimitives.scala 124:33:@34369.4]
    .clock(StickySelects_17_clock),
    .reset(StickySelects_17_reset),
    .io_ins_0(StickySelects_17_io_ins_0),
    .io_ins_1(StickySelects_17_io_ins_1),
    .io_ins_2(StickySelects_17_io_ins_2),
    .io_ins_3(StickySelects_17_io_ins_3),
    .io_ins_4(StickySelects_17_io_ins_4),
    .io_ins_5(StickySelects_17_io_ins_5),
    .io_outs_0(StickySelects_17_io_outs_0),
    .io_outs_1(StickySelects_17_io_outs_1),
    .io_outs_2(StickySelects_17_io_outs_2),
    .io_outs_3(StickySelects_17_io_outs_3),
    .io_outs_4(StickySelects_17_io_outs_4),
    .io_outs_5(StickySelects_17_io_outs_5)
  );
  StickySelects_25 StickySelects_18 ( // @[MemPrimitives.scala 124:33:@34423.4]
    .clock(StickySelects_18_clock),
    .reset(StickySelects_18_reset),
    .io_ins_0(StickySelects_18_io_ins_0),
    .io_ins_1(StickySelects_18_io_ins_1),
    .io_ins_2(StickySelects_18_io_ins_2),
    .io_ins_3(StickySelects_18_io_ins_3),
    .io_outs_0(StickySelects_18_io_outs_0),
    .io_outs_1(StickySelects_18_io_outs_1),
    .io_outs_2(StickySelects_18_io_outs_2),
    .io_outs_3(StickySelects_18_io_outs_3)
  );
  StickySelects_26 StickySelects_19 ( // @[MemPrimitives.scala 124:33:@34475.4]
    .clock(StickySelects_19_clock),
    .reset(StickySelects_19_reset),
    .io_ins_0(StickySelects_19_io_ins_0),
    .io_ins_1(StickySelects_19_io_ins_1),
    .io_ins_2(StickySelects_19_io_ins_2),
    .io_ins_3(StickySelects_19_io_ins_3),
    .io_ins_4(StickySelects_19_io_ins_4),
    .io_ins_5(StickySelects_19_io_ins_5),
    .io_outs_0(StickySelects_19_io_outs_0),
    .io_outs_1(StickySelects_19_io_outs_1),
    .io_outs_2(StickySelects_19_io_outs_2),
    .io_outs_3(StickySelects_19_io_outs_3),
    .io_outs_4(StickySelects_19_io_outs_4),
    .io_outs_5(StickySelects_19_io_outs_5)
  );
  StickySelects_25 StickySelects_20 ( // @[MemPrimitives.scala 124:33:@34529.4]
    .clock(StickySelects_20_clock),
    .reset(StickySelects_20_reset),
    .io_ins_0(StickySelects_20_io_ins_0),
    .io_ins_1(StickySelects_20_io_ins_1),
    .io_ins_2(StickySelects_20_io_ins_2),
    .io_ins_3(StickySelects_20_io_ins_3),
    .io_outs_0(StickySelects_20_io_outs_0),
    .io_outs_1(StickySelects_20_io_outs_1),
    .io_outs_2(StickySelects_20_io_outs_2),
    .io_outs_3(StickySelects_20_io_outs_3)
  );
  StickySelects_26 StickySelects_21 ( // @[MemPrimitives.scala 124:33:@34581.4]
    .clock(StickySelects_21_clock),
    .reset(StickySelects_21_reset),
    .io_ins_0(StickySelects_21_io_ins_0),
    .io_ins_1(StickySelects_21_io_ins_1),
    .io_ins_2(StickySelects_21_io_ins_2),
    .io_ins_3(StickySelects_21_io_ins_3),
    .io_ins_4(StickySelects_21_io_ins_4),
    .io_ins_5(StickySelects_21_io_ins_5),
    .io_outs_0(StickySelects_21_io_outs_0),
    .io_outs_1(StickySelects_21_io_outs_1),
    .io_outs_2(StickySelects_21_io_outs_2),
    .io_outs_3(StickySelects_21_io_outs_3),
    .io_outs_4(StickySelects_21_io_outs_4),
    .io_outs_5(StickySelects_21_io_outs_5)
  );
  StickySelects_25 StickySelects_22 ( // @[MemPrimitives.scala 124:33:@34635.4]
    .clock(StickySelects_22_clock),
    .reset(StickySelects_22_reset),
    .io_ins_0(StickySelects_22_io_ins_0),
    .io_ins_1(StickySelects_22_io_ins_1),
    .io_ins_2(StickySelects_22_io_ins_2),
    .io_ins_3(StickySelects_22_io_ins_3),
    .io_outs_0(StickySelects_22_io_outs_0),
    .io_outs_1(StickySelects_22_io_outs_1),
    .io_outs_2(StickySelects_22_io_outs_2),
    .io_outs_3(StickySelects_22_io_outs_3)
  );
  StickySelects_26 StickySelects_23 ( // @[MemPrimitives.scala 124:33:@34687.4]
    .clock(StickySelects_23_clock),
    .reset(StickySelects_23_reset),
    .io_ins_0(StickySelects_23_io_ins_0),
    .io_ins_1(StickySelects_23_io_ins_1),
    .io_ins_2(StickySelects_23_io_ins_2),
    .io_ins_3(StickySelects_23_io_ins_3),
    .io_ins_4(StickySelects_23_io_ins_4),
    .io_ins_5(StickySelects_23_io_ins_5),
    .io_outs_0(StickySelects_23_io_outs_0),
    .io_outs_1(StickySelects_23_io_outs_1),
    .io_outs_2(StickySelects_23_io_outs_2),
    .io_outs_3(StickySelects_23_io_outs_3),
    .io_outs_4(StickySelects_23_io_outs_4),
    .io_outs_5(StickySelects_23_io_outs_5)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@34762.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@34770.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@34778.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@34786.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@34794.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@34802.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@34810.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@34818.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@34826.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@34834.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@34842.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@34850.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@34906.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@34914.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@34922.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@34930.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@34938.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@34946.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@34954.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@34962.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@34970.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@34978.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@34986.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@34994.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@35050.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@35058.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@35066.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@35074.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@35082.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@35090.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@35098.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@35106.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@35114.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@35122.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@35130.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@35138.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@35194.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@35202.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@35210.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@35218.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@35226.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@35234.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@35242.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@35250.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@35258.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@35266.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@35274.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@35282.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@35338.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@35346.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@35354.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@35362.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@35370.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@35378.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@35386.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@35394.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@35402.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@35410.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@35418.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@35426.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@35482.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@35490.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@35498.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@35506.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@35514.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@35522.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@35530.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@35538.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@35546.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@35554.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@35562.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@35570.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@35626.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@35634.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@35642.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@35650.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@35658.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@35666.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@35674.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@35682.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@35690.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@35698.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@35706.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@35714.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@35770.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@35778.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@35786.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@35794.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@35802.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@35810.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@35818.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@35826.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@35834.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@35842.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@35850.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@35858.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_96 ( // @[package.scala 93:22:@35914.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_97 ( // @[package.scala 93:22:@35922.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_98 ( // @[package.scala 93:22:@35930.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_99 ( // @[package.scala 93:22:@35938.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_100 ( // @[package.scala 93:22:@35946.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_101 ( // @[package.scala 93:22:@35954.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_102 ( // @[package.scala 93:22:@35962.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_103 ( // @[package.scala 93:22:@35970.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_104 ( // @[package.scala 93:22:@35978.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_105 ( // @[package.scala 93:22:@35986.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_106 ( // @[package.scala 93:22:@35994.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_107 ( // @[package.scala 93:22:@36002.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_108 ( // @[package.scala 93:22:@36058.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_109 ( // @[package.scala 93:22:@36066.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_110 ( // @[package.scala 93:22:@36074.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_111 ( // @[package.scala 93:22:@36082.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_112 ( // @[package.scala 93:22:@36090.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_113 ( // @[package.scala 93:22:@36098.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_114 ( // @[package.scala 93:22:@36106.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_115 ( // @[package.scala 93:22:@36114.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_116 ( // @[package.scala 93:22:@36122.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_117 ( // @[package.scala 93:22:@36130.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_118 ( // @[package.scala 93:22:@36138.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_119 ( // @[package.scala 93:22:@36146.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  assign _T_460 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@32997.4]
  assign _T_462 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@32998.4]
  assign _T_463 = _T_460 & _T_462; // @[MemPrimitives.scala 82:228:@32999.4]
  assign _T_464 = io_wPort_0_en_0 & _T_463; // @[MemPrimitives.scala 83:102:@33000.4]
  assign _T_466 = io_wPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@33001.4]
  assign _T_468 = io_wPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@33002.4]
  assign _T_469 = _T_466 & _T_468; // @[MemPrimitives.scala 82:228:@33003.4]
  assign _T_470 = io_wPort_2_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@33004.4]
  assign _T_472 = {_T_464,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33006.4]
  assign _T_474 = {_T_470,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33008.4]
  assign _T_475 = _T_464 ? _T_472 : _T_474; // @[Mux.scala 31:69:@33009.4]
  assign _T_480 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@33016.4]
  assign _T_482 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@33017.4]
  assign _T_483 = _T_480 & _T_482; // @[MemPrimitives.scala 82:228:@33018.4]
  assign _T_484 = io_wPort_1_en_0 & _T_483; // @[MemPrimitives.scala 83:102:@33019.4]
  assign _T_486 = io_wPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@33020.4]
  assign _T_488 = io_wPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@33021.4]
  assign _T_489 = _T_486 & _T_488; // @[MemPrimitives.scala 82:228:@33022.4]
  assign _T_490 = io_wPort_3_en_0 & _T_489; // @[MemPrimitives.scala 83:102:@33023.4]
  assign _T_492 = {_T_484,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33025.4]
  assign _T_494 = {_T_490,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33027.4]
  assign _T_495 = _T_484 ? _T_492 : _T_494; // @[Mux.scala 31:69:@33028.4]
  assign _T_502 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@33036.4]
  assign _T_503 = _T_460 & _T_502; // @[MemPrimitives.scala 82:228:@33037.4]
  assign _T_504 = io_wPort_0_en_0 & _T_503; // @[MemPrimitives.scala 83:102:@33038.4]
  assign _T_508 = io_wPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@33040.4]
  assign _T_509 = _T_466 & _T_508; // @[MemPrimitives.scala 82:228:@33041.4]
  assign _T_510 = io_wPort_2_en_0 & _T_509; // @[MemPrimitives.scala 83:102:@33042.4]
  assign _T_512 = {_T_504,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33044.4]
  assign _T_514 = {_T_510,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33046.4]
  assign _T_515 = _T_504 ? _T_512 : _T_514; // @[Mux.scala 31:69:@33047.4]
  assign _T_522 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@33055.4]
  assign _T_523 = _T_480 & _T_522; // @[MemPrimitives.scala 82:228:@33056.4]
  assign _T_524 = io_wPort_1_en_0 & _T_523; // @[MemPrimitives.scala 83:102:@33057.4]
  assign _T_528 = io_wPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@33059.4]
  assign _T_529 = _T_486 & _T_528; // @[MemPrimitives.scala 82:228:@33060.4]
  assign _T_530 = io_wPort_3_en_0 & _T_529; // @[MemPrimitives.scala 83:102:@33061.4]
  assign _T_532 = {_T_524,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33063.4]
  assign _T_534 = {_T_530,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33065.4]
  assign _T_535 = _T_524 ? _T_532 : _T_534; // @[Mux.scala 31:69:@33066.4]
  assign _T_542 = io_wPort_0_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@33074.4]
  assign _T_543 = _T_460 & _T_542; // @[MemPrimitives.scala 82:228:@33075.4]
  assign _T_544 = io_wPort_0_en_0 & _T_543; // @[MemPrimitives.scala 83:102:@33076.4]
  assign _T_548 = io_wPort_2_banks_1 == 3'h4; // @[MemPrimitives.scala 82:210:@33078.4]
  assign _T_549 = _T_466 & _T_548; // @[MemPrimitives.scala 82:228:@33079.4]
  assign _T_550 = io_wPort_2_en_0 & _T_549; // @[MemPrimitives.scala 83:102:@33080.4]
  assign _T_552 = {_T_544,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33082.4]
  assign _T_554 = {_T_550,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33084.4]
  assign _T_555 = _T_544 ? _T_552 : _T_554; // @[Mux.scala 31:69:@33085.4]
  assign _T_562 = io_wPort_1_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@33093.4]
  assign _T_563 = _T_480 & _T_562; // @[MemPrimitives.scala 82:228:@33094.4]
  assign _T_564 = io_wPort_1_en_0 & _T_563; // @[MemPrimitives.scala 83:102:@33095.4]
  assign _T_568 = io_wPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 82:210:@33097.4]
  assign _T_569 = _T_486 & _T_568; // @[MemPrimitives.scala 82:228:@33098.4]
  assign _T_570 = io_wPort_3_en_0 & _T_569; // @[MemPrimitives.scala 83:102:@33099.4]
  assign _T_572 = {_T_564,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33101.4]
  assign _T_574 = {_T_570,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33103.4]
  assign _T_575 = _T_564 ? _T_572 : _T_574; // @[Mux.scala 31:69:@33104.4]
  assign _T_580 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@33111.4]
  assign _T_583 = _T_580 & _T_462; // @[MemPrimitives.scala 82:228:@33113.4]
  assign _T_584 = io_wPort_0_en_0 & _T_583; // @[MemPrimitives.scala 83:102:@33114.4]
  assign _T_586 = io_wPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@33115.4]
  assign _T_589 = _T_586 & _T_468; // @[MemPrimitives.scala 82:228:@33117.4]
  assign _T_590 = io_wPort_2_en_0 & _T_589; // @[MemPrimitives.scala 83:102:@33118.4]
  assign _T_592 = {_T_584,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33120.4]
  assign _T_594 = {_T_590,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33122.4]
  assign _T_595 = _T_584 ? _T_592 : _T_594; // @[Mux.scala 31:69:@33123.4]
  assign _T_600 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@33130.4]
  assign _T_603 = _T_600 & _T_482; // @[MemPrimitives.scala 82:228:@33132.4]
  assign _T_604 = io_wPort_1_en_0 & _T_603; // @[MemPrimitives.scala 83:102:@33133.4]
  assign _T_606 = io_wPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@33134.4]
  assign _T_609 = _T_606 & _T_488; // @[MemPrimitives.scala 82:228:@33136.4]
  assign _T_610 = io_wPort_3_en_0 & _T_609; // @[MemPrimitives.scala 83:102:@33137.4]
  assign _T_612 = {_T_604,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33139.4]
  assign _T_614 = {_T_610,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33141.4]
  assign _T_615 = _T_604 ? _T_612 : _T_614; // @[Mux.scala 31:69:@33142.4]
  assign _T_623 = _T_580 & _T_502; // @[MemPrimitives.scala 82:228:@33151.4]
  assign _T_624 = io_wPort_0_en_0 & _T_623; // @[MemPrimitives.scala 83:102:@33152.4]
  assign _T_629 = _T_586 & _T_508; // @[MemPrimitives.scala 82:228:@33155.4]
  assign _T_630 = io_wPort_2_en_0 & _T_629; // @[MemPrimitives.scala 83:102:@33156.4]
  assign _T_632 = {_T_624,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33158.4]
  assign _T_634 = {_T_630,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33160.4]
  assign _T_635 = _T_624 ? _T_632 : _T_634; // @[Mux.scala 31:69:@33161.4]
  assign _T_643 = _T_600 & _T_522; // @[MemPrimitives.scala 82:228:@33170.4]
  assign _T_644 = io_wPort_1_en_0 & _T_643; // @[MemPrimitives.scala 83:102:@33171.4]
  assign _T_649 = _T_606 & _T_528; // @[MemPrimitives.scala 82:228:@33174.4]
  assign _T_650 = io_wPort_3_en_0 & _T_649; // @[MemPrimitives.scala 83:102:@33175.4]
  assign _T_652 = {_T_644,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33177.4]
  assign _T_654 = {_T_650,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33179.4]
  assign _T_655 = _T_644 ? _T_652 : _T_654; // @[Mux.scala 31:69:@33180.4]
  assign _T_663 = _T_580 & _T_542; // @[MemPrimitives.scala 82:228:@33189.4]
  assign _T_664 = io_wPort_0_en_0 & _T_663; // @[MemPrimitives.scala 83:102:@33190.4]
  assign _T_669 = _T_586 & _T_548; // @[MemPrimitives.scala 82:228:@33193.4]
  assign _T_670 = io_wPort_2_en_0 & _T_669; // @[MemPrimitives.scala 83:102:@33194.4]
  assign _T_672 = {_T_664,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33196.4]
  assign _T_674 = {_T_670,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33198.4]
  assign _T_675 = _T_664 ? _T_672 : _T_674; // @[Mux.scala 31:69:@33199.4]
  assign _T_683 = _T_600 & _T_562; // @[MemPrimitives.scala 82:228:@33208.4]
  assign _T_684 = io_wPort_1_en_0 & _T_683; // @[MemPrimitives.scala 83:102:@33209.4]
  assign _T_689 = _T_606 & _T_568; // @[MemPrimitives.scala 82:228:@33212.4]
  assign _T_690 = io_wPort_3_en_0 & _T_689; // @[MemPrimitives.scala 83:102:@33213.4]
  assign _T_692 = {_T_684,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33215.4]
  assign _T_694 = {_T_690,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33217.4]
  assign _T_695 = _T_684 ? _T_692 : _T_694; // @[Mux.scala 31:69:@33218.4]
  assign _T_700 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@33225.4]
  assign _T_703 = _T_700 & _T_462; // @[MemPrimitives.scala 82:228:@33227.4]
  assign _T_704 = io_wPort_0_en_0 & _T_703; // @[MemPrimitives.scala 83:102:@33228.4]
  assign _T_706 = io_wPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@33229.4]
  assign _T_709 = _T_706 & _T_468; // @[MemPrimitives.scala 82:228:@33231.4]
  assign _T_710 = io_wPort_2_en_0 & _T_709; // @[MemPrimitives.scala 83:102:@33232.4]
  assign _T_712 = {_T_704,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33234.4]
  assign _T_714 = {_T_710,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33236.4]
  assign _T_715 = _T_704 ? _T_712 : _T_714; // @[Mux.scala 31:69:@33237.4]
  assign _T_720 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@33244.4]
  assign _T_723 = _T_720 & _T_482; // @[MemPrimitives.scala 82:228:@33246.4]
  assign _T_724 = io_wPort_1_en_0 & _T_723; // @[MemPrimitives.scala 83:102:@33247.4]
  assign _T_726 = io_wPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@33248.4]
  assign _T_729 = _T_726 & _T_488; // @[MemPrimitives.scala 82:228:@33250.4]
  assign _T_730 = io_wPort_3_en_0 & _T_729; // @[MemPrimitives.scala 83:102:@33251.4]
  assign _T_732 = {_T_724,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33253.4]
  assign _T_734 = {_T_730,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33255.4]
  assign _T_735 = _T_724 ? _T_732 : _T_734; // @[Mux.scala 31:69:@33256.4]
  assign _T_743 = _T_700 & _T_502; // @[MemPrimitives.scala 82:228:@33265.4]
  assign _T_744 = io_wPort_0_en_0 & _T_743; // @[MemPrimitives.scala 83:102:@33266.4]
  assign _T_749 = _T_706 & _T_508; // @[MemPrimitives.scala 82:228:@33269.4]
  assign _T_750 = io_wPort_2_en_0 & _T_749; // @[MemPrimitives.scala 83:102:@33270.4]
  assign _T_752 = {_T_744,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33272.4]
  assign _T_754 = {_T_750,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33274.4]
  assign _T_755 = _T_744 ? _T_752 : _T_754; // @[Mux.scala 31:69:@33275.4]
  assign _T_763 = _T_720 & _T_522; // @[MemPrimitives.scala 82:228:@33284.4]
  assign _T_764 = io_wPort_1_en_0 & _T_763; // @[MemPrimitives.scala 83:102:@33285.4]
  assign _T_769 = _T_726 & _T_528; // @[MemPrimitives.scala 82:228:@33288.4]
  assign _T_770 = io_wPort_3_en_0 & _T_769; // @[MemPrimitives.scala 83:102:@33289.4]
  assign _T_772 = {_T_764,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33291.4]
  assign _T_774 = {_T_770,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33293.4]
  assign _T_775 = _T_764 ? _T_772 : _T_774; // @[Mux.scala 31:69:@33294.4]
  assign _T_783 = _T_700 & _T_542; // @[MemPrimitives.scala 82:228:@33303.4]
  assign _T_784 = io_wPort_0_en_0 & _T_783; // @[MemPrimitives.scala 83:102:@33304.4]
  assign _T_789 = _T_706 & _T_548; // @[MemPrimitives.scala 82:228:@33307.4]
  assign _T_790 = io_wPort_2_en_0 & _T_789; // @[MemPrimitives.scala 83:102:@33308.4]
  assign _T_792 = {_T_784,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33310.4]
  assign _T_794 = {_T_790,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33312.4]
  assign _T_795 = _T_784 ? _T_792 : _T_794; // @[Mux.scala 31:69:@33313.4]
  assign _T_803 = _T_720 & _T_562; // @[MemPrimitives.scala 82:228:@33322.4]
  assign _T_804 = io_wPort_1_en_0 & _T_803; // @[MemPrimitives.scala 83:102:@33323.4]
  assign _T_809 = _T_726 & _T_568; // @[MemPrimitives.scala 82:228:@33326.4]
  assign _T_810 = io_wPort_3_en_0 & _T_809; // @[MemPrimitives.scala 83:102:@33327.4]
  assign _T_812 = {_T_804,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33329.4]
  assign _T_814 = {_T_810,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33331.4]
  assign _T_815 = _T_804 ? _T_812 : _T_814; // @[Mux.scala 31:69:@33332.4]
  assign _T_820 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@33339.4]
  assign _T_823 = _T_820 & _T_462; // @[MemPrimitives.scala 82:228:@33341.4]
  assign _T_824 = io_wPort_0_en_0 & _T_823; // @[MemPrimitives.scala 83:102:@33342.4]
  assign _T_826 = io_wPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@33343.4]
  assign _T_829 = _T_826 & _T_468; // @[MemPrimitives.scala 82:228:@33345.4]
  assign _T_830 = io_wPort_2_en_0 & _T_829; // @[MemPrimitives.scala 83:102:@33346.4]
  assign _T_832 = {_T_824,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33348.4]
  assign _T_834 = {_T_830,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33350.4]
  assign _T_835 = _T_824 ? _T_832 : _T_834; // @[Mux.scala 31:69:@33351.4]
  assign _T_840 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@33358.4]
  assign _T_843 = _T_840 & _T_482; // @[MemPrimitives.scala 82:228:@33360.4]
  assign _T_844 = io_wPort_1_en_0 & _T_843; // @[MemPrimitives.scala 83:102:@33361.4]
  assign _T_846 = io_wPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@33362.4]
  assign _T_849 = _T_846 & _T_488; // @[MemPrimitives.scala 82:228:@33364.4]
  assign _T_850 = io_wPort_3_en_0 & _T_849; // @[MemPrimitives.scala 83:102:@33365.4]
  assign _T_852 = {_T_844,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33367.4]
  assign _T_854 = {_T_850,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33369.4]
  assign _T_855 = _T_844 ? _T_852 : _T_854; // @[Mux.scala 31:69:@33370.4]
  assign _T_863 = _T_820 & _T_502; // @[MemPrimitives.scala 82:228:@33379.4]
  assign _T_864 = io_wPort_0_en_0 & _T_863; // @[MemPrimitives.scala 83:102:@33380.4]
  assign _T_869 = _T_826 & _T_508; // @[MemPrimitives.scala 82:228:@33383.4]
  assign _T_870 = io_wPort_2_en_0 & _T_869; // @[MemPrimitives.scala 83:102:@33384.4]
  assign _T_872 = {_T_864,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33386.4]
  assign _T_874 = {_T_870,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33388.4]
  assign _T_875 = _T_864 ? _T_872 : _T_874; // @[Mux.scala 31:69:@33389.4]
  assign _T_883 = _T_840 & _T_522; // @[MemPrimitives.scala 82:228:@33398.4]
  assign _T_884 = io_wPort_1_en_0 & _T_883; // @[MemPrimitives.scala 83:102:@33399.4]
  assign _T_889 = _T_846 & _T_528; // @[MemPrimitives.scala 82:228:@33402.4]
  assign _T_890 = io_wPort_3_en_0 & _T_889; // @[MemPrimitives.scala 83:102:@33403.4]
  assign _T_892 = {_T_884,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33405.4]
  assign _T_894 = {_T_890,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33407.4]
  assign _T_895 = _T_884 ? _T_892 : _T_894; // @[Mux.scala 31:69:@33408.4]
  assign _T_903 = _T_820 & _T_542; // @[MemPrimitives.scala 82:228:@33417.4]
  assign _T_904 = io_wPort_0_en_0 & _T_903; // @[MemPrimitives.scala 83:102:@33418.4]
  assign _T_909 = _T_826 & _T_548; // @[MemPrimitives.scala 82:228:@33421.4]
  assign _T_910 = io_wPort_2_en_0 & _T_909; // @[MemPrimitives.scala 83:102:@33422.4]
  assign _T_912 = {_T_904,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@33424.4]
  assign _T_914 = {_T_910,io_wPort_2_data_0,io_wPort_2_ofs_0}; // @[Cat.scala 30:58:@33426.4]
  assign _T_915 = _T_904 ? _T_912 : _T_914; // @[Mux.scala 31:69:@33427.4]
  assign _T_923 = _T_840 & _T_562; // @[MemPrimitives.scala 82:228:@33436.4]
  assign _T_924 = io_wPort_1_en_0 & _T_923; // @[MemPrimitives.scala 83:102:@33437.4]
  assign _T_929 = _T_846 & _T_568; // @[MemPrimitives.scala 82:228:@33440.4]
  assign _T_930 = io_wPort_3_en_0 & _T_929; // @[MemPrimitives.scala 83:102:@33441.4]
  assign _T_932 = {_T_924,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@33443.4]
  assign _T_934 = {_T_930,io_wPort_3_data_0,io_wPort_3_ofs_0}; // @[Cat.scala 30:58:@33445.4]
  assign _T_935 = _T_924 ? _T_932 : _T_934; // @[Mux.scala 31:69:@33446.4]
  assign _T_940 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33453.4]
  assign _T_942 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@33454.4]
  assign _T_943 = _T_940 & _T_942; // @[MemPrimitives.scala 110:228:@33455.4]
  assign _T_946 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33457.4]
  assign _T_948 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@33458.4]
  assign _T_949 = _T_946 & _T_948; // @[MemPrimitives.scala 110:228:@33459.4]
  assign _T_952 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33461.4]
  assign _T_954 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@33462.4]
  assign _T_955 = _T_952 & _T_954; // @[MemPrimitives.scala 110:228:@33463.4]
  assign _T_958 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33465.4]
  assign _T_960 = io_rPort_9_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@33466.4]
  assign _T_961 = _T_958 & _T_960; // @[MemPrimitives.scala 110:228:@33467.4]
  assign _T_963 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@33476.4]
  assign _T_964 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@33477.4]
  assign _T_965 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@33478.4]
  assign _T_966 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@33479.4]
  assign _T_968 = {_T_963,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@33481.4]
  assign _T_970 = {_T_964,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@33483.4]
  assign _T_972 = {_T_965,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@33485.4]
  assign _T_974 = {_T_966,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@33487.4]
  assign _T_975 = _T_965 ? _T_972 : _T_974; // @[Mux.scala 31:69:@33488.4]
  assign _T_976 = _T_964 ? _T_970 : _T_975; // @[Mux.scala 31:69:@33489.4]
  assign _T_977 = _T_963 ? _T_968 : _T_976; // @[Mux.scala 31:69:@33490.4]
  assign _T_982 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33497.4]
  assign _T_984 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@33498.4]
  assign _T_985 = _T_982 & _T_984; // @[MemPrimitives.scala 110:228:@33499.4]
  assign _T_988 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33501.4]
  assign _T_990 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@33502.4]
  assign _T_991 = _T_988 & _T_990; // @[MemPrimitives.scala 110:228:@33503.4]
  assign _T_994 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33505.4]
  assign _T_996 = io_rPort_2_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@33506.4]
  assign _T_997 = _T_994 & _T_996; // @[MemPrimitives.scala 110:228:@33507.4]
  assign _T_1000 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33509.4]
  assign _T_1002 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@33510.4]
  assign _T_1003 = _T_1000 & _T_1002; // @[MemPrimitives.scala 110:228:@33511.4]
  assign _T_1006 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33513.4]
  assign _T_1008 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@33514.4]
  assign _T_1009 = _T_1006 & _T_1008; // @[MemPrimitives.scala 110:228:@33515.4]
  assign _T_1012 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@33517.4]
  assign _T_1014 = io_rPort_8_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@33518.4]
  assign _T_1015 = _T_1012 & _T_1014; // @[MemPrimitives.scala 110:228:@33519.4]
  assign _T_1017 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@33530.4]
  assign _T_1018 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@33531.4]
  assign _T_1019 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@33532.4]
  assign _T_1020 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@33533.4]
  assign _T_1021 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@33534.4]
  assign _T_1022 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@33535.4]
  assign _T_1024 = {_T_1017,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@33537.4]
  assign _T_1026 = {_T_1018,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@33539.4]
  assign _T_1028 = {_T_1019,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@33541.4]
  assign _T_1030 = {_T_1020,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@33543.4]
  assign _T_1032 = {_T_1021,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@33545.4]
  assign _T_1034 = {_T_1022,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@33547.4]
  assign _T_1035 = _T_1021 ? _T_1032 : _T_1034; // @[Mux.scala 31:69:@33548.4]
  assign _T_1036 = _T_1020 ? _T_1030 : _T_1035; // @[Mux.scala 31:69:@33549.4]
  assign _T_1037 = _T_1019 ? _T_1028 : _T_1036; // @[Mux.scala 31:69:@33550.4]
  assign _T_1038 = _T_1018 ? _T_1026 : _T_1037; // @[Mux.scala 31:69:@33551.4]
  assign _T_1039 = _T_1017 ? _T_1024 : _T_1038; // @[Mux.scala 31:69:@33552.4]
  assign _T_1046 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@33560.4]
  assign _T_1047 = _T_940 & _T_1046; // @[MemPrimitives.scala 110:228:@33561.4]
  assign _T_1052 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@33564.4]
  assign _T_1053 = _T_946 & _T_1052; // @[MemPrimitives.scala 110:228:@33565.4]
  assign _T_1058 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@33568.4]
  assign _T_1059 = _T_952 & _T_1058; // @[MemPrimitives.scala 110:228:@33569.4]
  assign _T_1064 = io_rPort_9_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@33572.4]
  assign _T_1065 = _T_958 & _T_1064; // @[MemPrimitives.scala 110:228:@33573.4]
  assign _T_1067 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@33582.4]
  assign _T_1068 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@33583.4]
  assign _T_1069 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@33584.4]
  assign _T_1070 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@33585.4]
  assign _T_1072 = {_T_1067,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@33587.4]
  assign _T_1074 = {_T_1068,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@33589.4]
  assign _T_1076 = {_T_1069,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@33591.4]
  assign _T_1078 = {_T_1070,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@33593.4]
  assign _T_1079 = _T_1069 ? _T_1076 : _T_1078; // @[Mux.scala 31:69:@33594.4]
  assign _T_1080 = _T_1068 ? _T_1074 : _T_1079; // @[Mux.scala 31:69:@33595.4]
  assign _T_1081 = _T_1067 ? _T_1072 : _T_1080; // @[Mux.scala 31:69:@33596.4]
  assign _T_1088 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@33604.4]
  assign _T_1089 = _T_982 & _T_1088; // @[MemPrimitives.scala 110:228:@33605.4]
  assign _T_1094 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@33608.4]
  assign _T_1095 = _T_988 & _T_1094; // @[MemPrimitives.scala 110:228:@33609.4]
  assign _T_1100 = io_rPort_2_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@33612.4]
  assign _T_1101 = _T_994 & _T_1100; // @[MemPrimitives.scala 110:228:@33613.4]
  assign _T_1106 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@33616.4]
  assign _T_1107 = _T_1000 & _T_1106; // @[MemPrimitives.scala 110:228:@33617.4]
  assign _T_1112 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@33620.4]
  assign _T_1113 = _T_1006 & _T_1112; // @[MemPrimitives.scala 110:228:@33621.4]
  assign _T_1118 = io_rPort_8_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@33624.4]
  assign _T_1119 = _T_1012 & _T_1118; // @[MemPrimitives.scala 110:228:@33625.4]
  assign _T_1121 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@33636.4]
  assign _T_1122 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@33637.4]
  assign _T_1123 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@33638.4]
  assign _T_1124 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@33639.4]
  assign _T_1125 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@33640.4]
  assign _T_1126 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@33641.4]
  assign _T_1128 = {_T_1121,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@33643.4]
  assign _T_1130 = {_T_1122,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@33645.4]
  assign _T_1132 = {_T_1123,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@33647.4]
  assign _T_1134 = {_T_1124,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@33649.4]
  assign _T_1136 = {_T_1125,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@33651.4]
  assign _T_1138 = {_T_1126,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@33653.4]
  assign _T_1139 = _T_1125 ? _T_1136 : _T_1138; // @[Mux.scala 31:69:@33654.4]
  assign _T_1140 = _T_1124 ? _T_1134 : _T_1139; // @[Mux.scala 31:69:@33655.4]
  assign _T_1141 = _T_1123 ? _T_1132 : _T_1140; // @[Mux.scala 31:69:@33656.4]
  assign _T_1142 = _T_1122 ? _T_1130 : _T_1141; // @[Mux.scala 31:69:@33657.4]
  assign _T_1143 = _T_1121 ? _T_1128 : _T_1142; // @[Mux.scala 31:69:@33658.4]
  assign _T_1150 = io_rPort_4_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@33666.4]
  assign _T_1151 = _T_940 & _T_1150; // @[MemPrimitives.scala 110:228:@33667.4]
  assign _T_1156 = io_rPort_6_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@33670.4]
  assign _T_1157 = _T_946 & _T_1156; // @[MemPrimitives.scala 110:228:@33671.4]
  assign _T_1162 = io_rPort_7_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@33674.4]
  assign _T_1163 = _T_952 & _T_1162; // @[MemPrimitives.scala 110:228:@33675.4]
  assign _T_1168 = io_rPort_9_banks_1 == 3'h4; // @[MemPrimitives.scala 110:210:@33678.4]
  assign _T_1169 = _T_958 & _T_1168; // @[MemPrimitives.scala 110:228:@33679.4]
  assign _T_1171 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@33688.4]
  assign _T_1172 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@33689.4]
  assign _T_1173 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@33690.4]
  assign _T_1174 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@33691.4]
  assign _T_1176 = {_T_1171,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@33693.4]
  assign _T_1178 = {_T_1172,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@33695.4]
  assign _T_1180 = {_T_1173,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@33697.4]
  assign _T_1182 = {_T_1174,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@33699.4]
  assign _T_1183 = _T_1173 ? _T_1180 : _T_1182; // @[Mux.scala 31:69:@33700.4]
  assign _T_1184 = _T_1172 ? _T_1178 : _T_1183; // @[Mux.scala 31:69:@33701.4]
  assign _T_1185 = _T_1171 ? _T_1176 : _T_1184; // @[Mux.scala 31:69:@33702.4]
  assign _T_1192 = io_rPort_0_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@33710.4]
  assign _T_1193 = _T_982 & _T_1192; // @[MemPrimitives.scala 110:228:@33711.4]
  assign _T_1198 = io_rPort_1_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@33714.4]
  assign _T_1199 = _T_988 & _T_1198; // @[MemPrimitives.scala 110:228:@33715.4]
  assign _T_1204 = io_rPort_2_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@33718.4]
  assign _T_1205 = _T_994 & _T_1204; // @[MemPrimitives.scala 110:228:@33719.4]
  assign _T_1210 = io_rPort_3_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@33722.4]
  assign _T_1211 = _T_1000 & _T_1210; // @[MemPrimitives.scala 110:228:@33723.4]
  assign _T_1216 = io_rPort_5_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@33726.4]
  assign _T_1217 = _T_1006 & _T_1216; // @[MemPrimitives.scala 110:228:@33727.4]
  assign _T_1222 = io_rPort_8_banks_1 == 3'h5; // @[MemPrimitives.scala 110:210:@33730.4]
  assign _T_1223 = _T_1012 & _T_1222; // @[MemPrimitives.scala 110:228:@33731.4]
  assign _T_1225 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@33742.4]
  assign _T_1226 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@33743.4]
  assign _T_1227 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@33744.4]
  assign _T_1228 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@33745.4]
  assign _T_1229 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@33746.4]
  assign _T_1230 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@33747.4]
  assign _T_1232 = {_T_1225,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@33749.4]
  assign _T_1234 = {_T_1226,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@33751.4]
  assign _T_1236 = {_T_1227,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@33753.4]
  assign _T_1238 = {_T_1228,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@33755.4]
  assign _T_1240 = {_T_1229,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@33757.4]
  assign _T_1242 = {_T_1230,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@33759.4]
  assign _T_1243 = _T_1229 ? _T_1240 : _T_1242; // @[Mux.scala 31:69:@33760.4]
  assign _T_1244 = _T_1228 ? _T_1238 : _T_1243; // @[Mux.scala 31:69:@33761.4]
  assign _T_1245 = _T_1227 ? _T_1236 : _T_1244; // @[Mux.scala 31:69:@33762.4]
  assign _T_1246 = _T_1226 ? _T_1234 : _T_1245; // @[Mux.scala 31:69:@33763.4]
  assign _T_1247 = _T_1225 ? _T_1232 : _T_1246; // @[Mux.scala 31:69:@33764.4]
  assign _T_1252 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33771.4]
  assign _T_1255 = _T_1252 & _T_942; // @[MemPrimitives.scala 110:228:@33773.4]
  assign _T_1258 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33775.4]
  assign _T_1261 = _T_1258 & _T_948; // @[MemPrimitives.scala 110:228:@33777.4]
  assign _T_1264 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33779.4]
  assign _T_1267 = _T_1264 & _T_954; // @[MemPrimitives.scala 110:228:@33781.4]
  assign _T_1270 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33783.4]
  assign _T_1273 = _T_1270 & _T_960; // @[MemPrimitives.scala 110:228:@33785.4]
  assign _T_1275 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@33794.4]
  assign _T_1276 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@33795.4]
  assign _T_1277 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@33796.4]
  assign _T_1278 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@33797.4]
  assign _T_1280 = {_T_1275,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@33799.4]
  assign _T_1282 = {_T_1276,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@33801.4]
  assign _T_1284 = {_T_1277,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@33803.4]
  assign _T_1286 = {_T_1278,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@33805.4]
  assign _T_1287 = _T_1277 ? _T_1284 : _T_1286; // @[Mux.scala 31:69:@33806.4]
  assign _T_1288 = _T_1276 ? _T_1282 : _T_1287; // @[Mux.scala 31:69:@33807.4]
  assign _T_1289 = _T_1275 ? _T_1280 : _T_1288; // @[Mux.scala 31:69:@33808.4]
  assign _T_1294 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33815.4]
  assign _T_1297 = _T_1294 & _T_984; // @[MemPrimitives.scala 110:228:@33817.4]
  assign _T_1300 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33819.4]
  assign _T_1303 = _T_1300 & _T_990; // @[MemPrimitives.scala 110:228:@33821.4]
  assign _T_1306 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33823.4]
  assign _T_1309 = _T_1306 & _T_996; // @[MemPrimitives.scala 110:228:@33825.4]
  assign _T_1312 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33827.4]
  assign _T_1315 = _T_1312 & _T_1002; // @[MemPrimitives.scala 110:228:@33829.4]
  assign _T_1318 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33831.4]
  assign _T_1321 = _T_1318 & _T_1008; // @[MemPrimitives.scala 110:228:@33833.4]
  assign _T_1324 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@33835.4]
  assign _T_1327 = _T_1324 & _T_1014; // @[MemPrimitives.scala 110:228:@33837.4]
  assign _T_1329 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@33848.4]
  assign _T_1330 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@33849.4]
  assign _T_1331 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@33850.4]
  assign _T_1332 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@33851.4]
  assign _T_1333 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@33852.4]
  assign _T_1334 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@33853.4]
  assign _T_1336 = {_T_1329,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@33855.4]
  assign _T_1338 = {_T_1330,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@33857.4]
  assign _T_1340 = {_T_1331,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@33859.4]
  assign _T_1342 = {_T_1332,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@33861.4]
  assign _T_1344 = {_T_1333,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@33863.4]
  assign _T_1346 = {_T_1334,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@33865.4]
  assign _T_1347 = _T_1333 ? _T_1344 : _T_1346; // @[Mux.scala 31:69:@33866.4]
  assign _T_1348 = _T_1332 ? _T_1342 : _T_1347; // @[Mux.scala 31:69:@33867.4]
  assign _T_1349 = _T_1331 ? _T_1340 : _T_1348; // @[Mux.scala 31:69:@33868.4]
  assign _T_1350 = _T_1330 ? _T_1338 : _T_1349; // @[Mux.scala 31:69:@33869.4]
  assign _T_1351 = _T_1329 ? _T_1336 : _T_1350; // @[Mux.scala 31:69:@33870.4]
  assign _T_1359 = _T_1252 & _T_1046; // @[MemPrimitives.scala 110:228:@33879.4]
  assign _T_1365 = _T_1258 & _T_1052; // @[MemPrimitives.scala 110:228:@33883.4]
  assign _T_1371 = _T_1264 & _T_1058; // @[MemPrimitives.scala 110:228:@33887.4]
  assign _T_1377 = _T_1270 & _T_1064; // @[MemPrimitives.scala 110:228:@33891.4]
  assign _T_1379 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@33900.4]
  assign _T_1380 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@33901.4]
  assign _T_1381 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@33902.4]
  assign _T_1382 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@33903.4]
  assign _T_1384 = {_T_1379,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@33905.4]
  assign _T_1386 = {_T_1380,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@33907.4]
  assign _T_1388 = {_T_1381,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@33909.4]
  assign _T_1390 = {_T_1382,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@33911.4]
  assign _T_1391 = _T_1381 ? _T_1388 : _T_1390; // @[Mux.scala 31:69:@33912.4]
  assign _T_1392 = _T_1380 ? _T_1386 : _T_1391; // @[Mux.scala 31:69:@33913.4]
  assign _T_1393 = _T_1379 ? _T_1384 : _T_1392; // @[Mux.scala 31:69:@33914.4]
  assign _T_1401 = _T_1294 & _T_1088; // @[MemPrimitives.scala 110:228:@33923.4]
  assign _T_1407 = _T_1300 & _T_1094; // @[MemPrimitives.scala 110:228:@33927.4]
  assign _T_1413 = _T_1306 & _T_1100; // @[MemPrimitives.scala 110:228:@33931.4]
  assign _T_1419 = _T_1312 & _T_1106; // @[MemPrimitives.scala 110:228:@33935.4]
  assign _T_1425 = _T_1318 & _T_1112; // @[MemPrimitives.scala 110:228:@33939.4]
  assign _T_1431 = _T_1324 & _T_1118; // @[MemPrimitives.scala 110:228:@33943.4]
  assign _T_1433 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@33954.4]
  assign _T_1434 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@33955.4]
  assign _T_1435 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@33956.4]
  assign _T_1436 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@33957.4]
  assign _T_1437 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@33958.4]
  assign _T_1438 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@33959.4]
  assign _T_1440 = {_T_1433,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@33961.4]
  assign _T_1442 = {_T_1434,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@33963.4]
  assign _T_1444 = {_T_1435,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@33965.4]
  assign _T_1446 = {_T_1436,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@33967.4]
  assign _T_1448 = {_T_1437,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@33969.4]
  assign _T_1450 = {_T_1438,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@33971.4]
  assign _T_1451 = _T_1437 ? _T_1448 : _T_1450; // @[Mux.scala 31:69:@33972.4]
  assign _T_1452 = _T_1436 ? _T_1446 : _T_1451; // @[Mux.scala 31:69:@33973.4]
  assign _T_1453 = _T_1435 ? _T_1444 : _T_1452; // @[Mux.scala 31:69:@33974.4]
  assign _T_1454 = _T_1434 ? _T_1442 : _T_1453; // @[Mux.scala 31:69:@33975.4]
  assign _T_1455 = _T_1433 ? _T_1440 : _T_1454; // @[Mux.scala 31:69:@33976.4]
  assign _T_1463 = _T_1252 & _T_1150; // @[MemPrimitives.scala 110:228:@33985.4]
  assign _T_1469 = _T_1258 & _T_1156; // @[MemPrimitives.scala 110:228:@33989.4]
  assign _T_1475 = _T_1264 & _T_1162; // @[MemPrimitives.scala 110:228:@33993.4]
  assign _T_1481 = _T_1270 & _T_1168; // @[MemPrimitives.scala 110:228:@33997.4]
  assign _T_1483 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@34006.4]
  assign _T_1484 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@34007.4]
  assign _T_1485 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@34008.4]
  assign _T_1486 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@34009.4]
  assign _T_1488 = {_T_1483,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@34011.4]
  assign _T_1490 = {_T_1484,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@34013.4]
  assign _T_1492 = {_T_1485,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@34015.4]
  assign _T_1494 = {_T_1486,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@34017.4]
  assign _T_1495 = _T_1485 ? _T_1492 : _T_1494; // @[Mux.scala 31:69:@34018.4]
  assign _T_1496 = _T_1484 ? _T_1490 : _T_1495; // @[Mux.scala 31:69:@34019.4]
  assign _T_1497 = _T_1483 ? _T_1488 : _T_1496; // @[Mux.scala 31:69:@34020.4]
  assign _T_1505 = _T_1294 & _T_1192; // @[MemPrimitives.scala 110:228:@34029.4]
  assign _T_1511 = _T_1300 & _T_1198; // @[MemPrimitives.scala 110:228:@34033.4]
  assign _T_1517 = _T_1306 & _T_1204; // @[MemPrimitives.scala 110:228:@34037.4]
  assign _T_1523 = _T_1312 & _T_1210; // @[MemPrimitives.scala 110:228:@34041.4]
  assign _T_1529 = _T_1318 & _T_1216; // @[MemPrimitives.scala 110:228:@34045.4]
  assign _T_1535 = _T_1324 & _T_1222; // @[MemPrimitives.scala 110:228:@34049.4]
  assign _T_1537 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@34060.4]
  assign _T_1538 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@34061.4]
  assign _T_1539 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@34062.4]
  assign _T_1540 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@34063.4]
  assign _T_1541 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@34064.4]
  assign _T_1542 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@34065.4]
  assign _T_1544 = {_T_1537,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@34067.4]
  assign _T_1546 = {_T_1538,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@34069.4]
  assign _T_1548 = {_T_1539,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@34071.4]
  assign _T_1550 = {_T_1540,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@34073.4]
  assign _T_1552 = {_T_1541,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@34075.4]
  assign _T_1554 = {_T_1542,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@34077.4]
  assign _T_1555 = _T_1541 ? _T_1552 : _T_1554; // @[Mux.scala 31:69:@34078.4]
  assign _T_1556 = _T_1540 ? _T_1550 : _T_1555; // @[Mux.scala 31:69:@34079.4]
  assign _T_1557 = _T_1539 ? _T_1548 : _T_1556; // @[Mux.scala 31:69:@34080.4]
  assign _T_1558 = _T_1538 ? _T_1546 : _T_1557; // @[Mux.scala 31:69:@34081.4]
  assign _T_1559 = _T_1537 ? _T_1544 : _T_1558; // @[Mux.scala 31:69:@34082.4]
  assign _T_1564 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34089.4]
  assign _T_1567 = _T_1564 & _T_942; // @[MemPrimitives.scala 110:228:@34091.4]
  assign _T_1570 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34093.4]
  assign _T_1573 = _T_1570 & _T_948; // @[MemPrimitives.scala 110:228:@34095.4]
  assign _T_1576 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34097.4]
  assign _T_1579 = _T_1576 & _T_954; // @[MemPrimitives.scala 110:228:@34099.4]
  assign _T_1582 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34101.4]
  assign _T_1585 = _T_1582 & _T_960; // @[MemPrimitives.scala 110:228:@34103.4]
  assign _T_1587 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@34112.4]
  assign _T_1588 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@34113.4]
  assign _T_1589 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@34114.4]
  assign _T_1590 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@34115.4]
  assign _T_1592 = {_T_1587,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@34117.4]
  assign _T_1594 = {_T_1588,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@34119.4]
  assign _T_1596 = {_T_1589,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@34121.4]
  assign _T_1598 = {_T_1590,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@34123.4]
  assign _T_1599 = _T_1589 ? _T_1596 : _T_1598; // @[Mux.scala 31:69:@34124.4]
  assign _T_1600 = _T_1588 ? _T_1594 : _T_1599; // @[Mux.scala 31:69:@34125.4]
  assign _T_1601 = _T_1587 ? _T_1592 : _T_1600; // @[Mux.scala 31:69:@34126.4]
  assign _T_1606 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34133.4]
  assign _T_1609 = _T_1606 & _T_984; // @[MemPrimitives.scala 110:228:@34135.4]
  assign _T_1612 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34137.4]
  assign _T_1615 = _T_1612 & _T_990; // @[MemPrimitives.scala 110:228:@34139.4]
  assign _T_1618 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34141.4]
  assign _T_1621 = _T_1618 & _T_996; // @[MemPrimitives.scala 110:228:@34143.4]
  assign _T_1624 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34145.4]
  assign _T_1627 = _T_1624 & _T_1002; // @[MemPrimitives.scala 110:228:@34147.4]
  assign _T_1630 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34149.4]
  assign _T_1633 = _T_1630 & _T_1008; // @[MemPrimitives.scala 110:228:@34151.4]
  assign _T_1636 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@34153.4]
  assign _T_1639 = _T_1636 & _T_1014; // @[MemPrimitives.scala 110:228:@34155.4]
  assign _T_1641 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@34166.4]
  assign _T_1642 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@34167.4]
  assign _T_1643 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@34168.4]
  assign _T_1644 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@34169.4]
  assign _T_1645 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@34170.4]
  assign _T_1646 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@34171.4]
  assign _T_1648 = {_T_1641,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@34173.4]
  assign _T_1650 = {_T_1642,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@34175.4]
  assign _T_1652 = {_T_1643,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@34177.4]
  assign _T_1654 = {_T_1644,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@34179.4]
  assign _T_1656 = {_T_1645,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@34181.4]
  assign _T_1658 = {_T_1646,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@34183.4]
  assign _T_1659 = _T_1645 ? _T_1656 : _T_1658; // @[Mux.scala 31:69:@34184.4]
  assign _T_1660 = _T_1644 ? _T_1654 : _T_1659; // @[Mux.scala 31:69:@34185.4]
  assign _T_1661 = _T_1643 ? _T_1652 : _T_1660; // @[Mux.scala 31:69:@34186.4]
  assign _T_1662 = _T_1642 ? _T_1650 : _T_1661; // @[Mux.scala 31:69:@34187.4]
  assign _T_1663 = _T_1641 ? _T_1648 : _T_1662; // @[Mux.scala 31:69:@34188.4]
  assign _T_1671 = _T_1564 & _T_1046; // @[MemPrimitives.scala 110:228:@34197.4]
  assign _T_1677 = _T_1570 & _T_1052; // @[MemPrimitives.scala 110:228:@34201.4]
  assign _T_1683 = _T_1576 & _T_1058; // @[MemPrimitives.scala 110:228:@34205.4]
  assign _T_1689 = _T_1582 & _T_1064; // @[MemPrimitives.scala 110:228:@34209.4]
  assign _T_1691 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@34218.4]
  assign _T_1692 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@34219.4]
  assign _T_1693 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@34220.4]
  assign _T_1694 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@34221.4]
  assign _T_1696 = {_T_1691,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@34223.4]
  assign _T_1698 = {_T_1692,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@34225.4]
  assign _T_1700 = {_T_1693,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@34227.4]
  assign _T_1702 = {_T_1694,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@34229.4]
  assign _T_1703 = _T_1693 ? _T_1700 : _T_1702; // @[Mux.scala 31:69:@34230.4]
  assign _T_1704 = _T_1692 ? _T_1698 : _T_1703; // @[Mux.scala 31:69:@34231.4]
  assign _T_1705 = _T_1691 ? _T_1696 : _T_1704; // @[Mux.scala 31:69:@34232.4]
  assign _T_1713 = _T_1606 & _T_1088; // @[MemPrimitives.scala 110:228:@34241.4]
  assign _T_1719 = _T_1612 & _T_1094; // @[MemPrimitives.scala 110:228:@34245.4]
  assign _T_1725 = _T_1618 & _T_1100; // @[MemPrimitives.scala 110:228:@34249.4]
  assign _T_1731 = _T_1624 & _T_1106; // @[MemPrimitives.scala 110:228:@34253.4]
  assign _T_1737 = _T_1630 & _T_1112; // @[MemPrimitives.scala 110:228:@34257.4]
  assign _T_1743 = _T_1636 & _T_1118; // @[MemPrimitives.scala 110:228:@34261.4]
  assign _T_1745 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@34272.4]
  assign _T_1746 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@34273.4]
  assign _T_1747 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@34274.4]
  assign _T_1748 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@34275.4]
  assign _T_1749 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@34276.4]
  assign _T_1750 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@34277.4]
  assign _T_1752 = {_T_1745,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@34279.4]
  assign _T_1754 = {_T_1746,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@34281.4]
  assign _T_1756 = {_T_1747,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@34283.4]
  assign _T_1758 = {_T_1748,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@34285.4]
  assign _T_1760 = {_T_1749,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@34287.4]
  assign _T_1762 = {_T_1750,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@34289.4]
  assign _T_1763 = _T_1749 ? _T_1760 : _T_1762; // @[Mux.scala 31:69:@34290.4]
  assign _T_1764 = _T_1748 ? _T_1758 : _T_1763; // @[Mux.scala 31:69:@34291.4]
  assign _T_1765 = _T_1747 ? _T_1756 : _T_1764; // @[Mux.scala 31:69:@34292.4]
  assign _T_1766 = _T_1746 ? _T_1754 : _T_1765; // @[Mux.scala 31:69:@34293.4]
  assign _T_1767 = _T_1745 ? _T_1752 : _T_1766; // @[Mux.scala 31:69:@34294.4]
  assign _T_1775 = _T_1564 & _T_1150; // @[MemPrimitives.scala 110:228:@34303.4]
  assign _T_1781 = _T_1570 & _T_1156; // @[MemPrimitives.scala 110:228:@34307.4]
  assign _T_1787 = _T_1576 & _T_1162; // @[MemPrimitives.scala 110:228:@34311.4]
  assign _T_1793 = _T_1582 & _T_1168; // @[MemPrimitives.scala 110:228:@34315.4]
  assign _T_1795 = StickySelects_16_io_outs_0; // @[MemPrimitives.scala 126:35:@34324.4]
  assign _T_1796 = StickySelects_16_io_outs_1; // @[MemPrimitives.scala 126:35:@34325.4]
  assign _T_1797 = StickySelects_16_io_outs_2; // @[MemPrimitives.scala 126:35:@34326.4]
  assign _T_1798 = StickySelects_16_io_outs_3; // @[MemPrimitives.scala 126:35:@34327.4]
  assign _T_1800 = {_T_1795,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@34329.4]
  assign _T_1802 = {_T_1796,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@34331.4]
  assign _T_1804 = {_T_1797,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@34333.4]
  assign _T_1806 = {_T_1798,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@34335.4]
  assign _T_1807 = _T_1797 ? _T_1804 : _T_1806; // @[Mux.scala 31:69:@34336.4]
  assign _T_1808 = _T_1796 ? _T_1802 : _T_1807; // @[Mux.scala 31:69:@34337.4]
  assign _T_1809 = _T_1795 ? _T_1800 : _T_1808; // @[Mux.scala 31:69:@34338.4]
  assign _T_1817 = _T_1606 & _T_1192; // @[MemPrimitives.scala 110:228:@34347.4]
  assign _T_1823 = _T_1612 & _T_1198; // @[MemPrimitives.scala 110:228:@34351.4]
  assign _T_1829 = _T_1618 & _T_1204; // @[MemPrimitives.scala 110:228:@34355.4]
  assign _T_1835 = _T_1624 & _T_1210; // @[MemPrimitives.scala 110:228:@34359.4]
  assign _T_1841 = _T_1630 & _T_1216; // @[MemPrimitives.scala 110:228:@34363.4]
  assign _T_1847 = _T_1636 & _T_1222; // @[MemPrimitives.scala 110:228:@34367.4]
  assign _T_1849 = StickySelects_17_io_outs_0; // @[MemPrimitives.scala 126:35:@34378.4]
  assign _T_1850 = StickySelects_17_io_outs_1; // @[MemPrimitives.scala 126:35:@34379.4]
  assign _T_1851 = StickySelects_17_io_outs_2; // @[MemPrimitives.scala 126:35:@34380.4]
  assign _T_1852 = StickySelects_17_io_outs_3; // @[MemPrimitives.scala 126:35:@34381.4]
  assign _T_1853 = StickySelects_17_io_outs_4; // @[MemPrimitives.scala 126:35:@34382.4]
  assign _T_1854 = StickySelects_17_io_outs_5; // @[MemPrimitives.scala 126:35:@34383.4]
  assign _T_1856 = {_T_1849,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@34385.4]
  assign _T_1858 = {_T_1850,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@34387.4]
  assign _T_1860 = {_T_1851,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@34389.4]
  assign _T_1862 = {_T_1852,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@34391.4]
  assign _T_1864 = {_T_1853,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@34393.4]
  assign _T_1866 = {_T_1854,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@34395.4]
  assign _T_1867 = _T_1853 ? _T_1864 : _T_1866; // @[Mux.scala 31:69:@34396.4]
  assign _T_1868 = _T_1852 ? _T_1862 : _T_1867; // @[Mux.scala 31:69:@34397.4]
  assign _T_1869 = _T_1851 ? _T_1860 : _T_1868; // @[Mux.scala 31:69:@34398.4]
  assign _T_1870 = _T_1850 ? _T_1858 : _T_1869; // @[Mux.scala 31:69:@34399.4]
  assign _T_1871 = _T_1849 ? _T_1856 : _T_1870; // @[Mux.scala 31:69:@34400.4]
  assign _T_1876 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34407.4]
  assign _T_1879 = _T_1876 & _T_942; // @[MemPrimitives.scala 110:228:@34409.4]
  assign _T_1882 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34411.4]
  assign _T_1885 = _T_1882 & _T_948; // @[MemPrimitives.scala 110:228:@34413.4]
  assign _T_1888 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34415.4]
  assign _T_1891 = _T_1888 & _T_954; // @[MemPrimitives.scala 110:228:@34417.4]
  assign _T_1894 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34419.4]
  assign _T_1897 = _T_1894 & _T_960; // @[MemPrimitives.scala 110:228:@34421.4]
  assign _T_1899 = StickySelects_18_io_outs_0; // @[MemPrimitives.scala 126:35:@34430.4]
  assign _T_1900 = StickySelects_18_io_outs_1; // @[MemPrimitives.scala 126:35:@34431.4]
  assign _T_1901 = StickySelects_18_io_outs_2; // @[MemPrimitives.scala 126:35:@34432.4]
  assign _T_1902 = StickySelects_18_io_outs_3; // @[MemPrimitives.scala 126:35:@34433.4]
  assign _T_1904 = {_T_1899,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@34435.4]
  assign _T_1906 = {_T_1900,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@34437.4]
  assign _T_1908 = {_T_1901,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@34439.4]
  assign _T_1910 = {_T_1902,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@34441.4]
  assign _T_1911 = _T_1901 ? _T_1908 : _T_1910; // @[Mux.scala 31:69:@34442.4]
  assign _T_1912 = _T_1900 ? _T_1906 : _T_1911; // @[Mux.scala 31:69:@34443.4]
  assign _T_1913 = _T_1899 ? _T_1904 : _T_1912; // @[Mux.scala 31:69:@34444.4]
  assign _T_1918 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34451.4]
  assign _T_1921 = _T_1918 & _T_984; // @[MemPrimitives.scala 110:228:@34453.4]
  assign _T_1924 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34455.4]
  assign _T_1927 = _T_1924 & _T_990; // @[MemPrimitives.scala 110:228:@34457.4]
  assign _T_1930 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34459.4]
  assign _T_1933 = _T_1930 & _T_996; // @[MemPrimitives.scala 110:228:@34461.4]
  assign _T_1936 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34463.4]
  assign _T_1939 = _T_1936 & _T_1002; // @[MemPrimitives.scala 110:228:@34465.4]
  assign _T_1942 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34467.4]
  assign _T_1945 = _T_1942 & _T_1008; // @[MemPrimitives.scala 110:228:@34469.4]
  assign _T_1948 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@34471.4]
  assign _T_1951 = _T_1948 & _T_1014; // @[MemPrimitives.scala 110:228:@34473.4]
  assign _T_1953 = StickySelects_19_io_outs_0; // @[MemPrimitives.scala 126:35:@34484.4]
  assign _T_1954 = StickySelects_19_io_outs_1; // @[MemPrimitives.scala 126:35:@34485.4]
  assign _T_1955 = StickySelects_19_io_outs_2; // @[MemPrimitives.scala 126:35:@34486.4]
  assign _T_1956 = StickySelects_19_io_outs_3; // @[MemPrimitives.scala 126:35:@34487.4]
  assign _T_1957 = StickySelects_19_io_outs_4; // @[MemPrimitives.scala 126:35:@34488.4]
  assign _T_1958 = StickySelects_19_io_outs_5; // @[MemPrimitives.scala 126:35:@34489.4]
  assign _T_1960 = {_T_1953,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@34491.4]
  assign _T_1962 = {_T_1954,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@34493.4]
  assign _T_1964 = {_T_1955,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@34495.4]
  assign _T_1966 = {_T_1956,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@34497.4]
  assign _T_1968 = {_T_1957,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@34499.4]
  assign _T_1970 = {_T_1958,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@34501.4]
  assign _T_1971 = _T_1957 ? _T_1968 : _T_1970; // @[Mux.scala 31:69:@34502.4]
  assign _T_1972 = _T_1956 ? _T_1966 : _T_1971; // @[Mux.scala 31:69:@34503.4]
  assign _T_1973 = _T_1955 ? _T_1964 : _T_1972; // @[Mux.scala 31:69:@34504.4]
  assign _T_1974 = _T_1954 ? _T_1962 : _T_1973; // @[Mux.scala 31:69:@34505.4]
  assign _T_1975 = _T_1953 ? _T_1960 : _T_1974; // @[Mux.scala 31:69:@34506.4]
  assign _T_1983 = _T_1876 & _T_1046; // @[MemPrimitives.scala 110:228:@34515.4]
  assign _T_1989 = _T_1882 & _T_1052; // @[MemPrimitives.scala 110:228:@34519.4]
  assign _T_1995 = _T_1888 & _T_1058; // @[MemPrimitives.scala 110:228:@34523.4]
  assign _T_2001 = _T_1894 & _T_1064; // @[MemPrimitives.scala 110:228:@34527.4]
  assign _T_2003 = StickySelects_20_io_outs_0; // @[MemPrimitives.scala 126:35:@34536.4]
  assign _T_2004 = StickySelects_20_io_outs_1; // @[MemPrimitives.scala 126:35:@34537.4]
  assign _T_2005 = StickySelects_20_io_outs_2; // @[MemPrimitives.scala 126:35:@34538.4]
  assign _T_2006 = StickySelects_20_io_outs_3; // @[MemPrimitives.scala 126:35:@34539.4]
  assign _T_2008 = {_T_2003,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@34541.4]
  assign _T_2010 = {_T_2004,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@34543.4]
  assign _T_2012 = {_T_2005,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@34545.4]
  assign _T_2014 = {_T_2006,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@34547.4]
  assign _T_2015 = _T_2005 ? _T_2012 : _T_2014; // @[Mux.scala 31:69:@34548.4]
  assign _T_2016 = _T_2004 ? _T_2010 : _T_2015; // @[Mux.scala 31:69:@34549.4]
  assign _T_2017 = _T_2003 ? _T_2008 : _T_2016; // @[Mux.scala 31:69:@34550.4]
  assign _T_2025 = _T_1918 & _T_1088; // @[MemPrimitives.scala 110:228:@34559.4]
  assign _T_2031 = _T_1924 & _T_1094; // @[MemPrimitives.scala 110:228:@34563.4]
  assign _T_2037 = _T_1930 & _T_1100; // @[MemPrimitives.scala 110:228:@34567.4]
  assign _T_2043 = _T_1936 & _T_1106; // @[MemPrimitives.scala 110:228:@34571.4]
  assign _T_2049 = _T_1942 & _T_1112; // @[MemPrimitives.scala 110:228:@34575.4]
  assign _T_2055 = _T_1948 & _T_1118; // @[MemPrimitives.scala 110:228:@34579.4]
  assign _T_2057 = StickySelects_21_io_outs_0; // @[MemPrimitives.scala 126:35:@34590.4]
  assign _T_2058 = StickySelects_21_io_outs_1; // @[MemPrimitives.scala 126:35:@34591.4]
  assign _T_2059 = StickySelects_21_io_outs_2; // @[MemPrimitives.scala 126:35:@34592.4]
  assign _T_2060 = StickySelects_21_io_outs_3; // @[MemPrimitives.scala 126:35:@34593.4]
  assign _T_2061 = StickySelects_21_io_outs_4; // @[MemPrimitives.scala 126:35:@34594.4]
  assign _T_2062 = StickySelects_21_io_outs_5; // @[MemPrimitives.scala 126:35:@34595.4]
  assign _T_2064 = {_T_2057,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@34597.4]
  assign _T_2066 = {_T_2058,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@34599.4]
  assign _T_2068 = {_T_2059,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@34601.4]
  assign _T_2070 = {_T_2060,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@34603.4]
  assign _T_2072 = {_T_2061,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@34605.4]
  assign _T_2074 = {_T_2062,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@34607.4]
  assign _T_2075 = _T_2061 ? _T_2072 : _T_2074; // @[Mux.scala 31:69:@34608.4]
  assign _T_2076 = _T_2060 ? _T_2070 : _T_2075; // @[Mux.scala 31:69:@34609.4]
  assign _T_2077 = _T_2059 ? _T_2068 : _T_2076; // @[Mux.scala 31:69:@34610.4]
  assign _T_2078 = _T_2058 ? _T_2066 : _T_2077; // @[Mux.scala 31:69:@34611.4]
  assign _T_2079 = _T_2057 ? _T_2064 : _T_2078; // @[Mux.scala 31:69:@34612.4]
  assign _T_2087 = _T_1876 & _T_1150; // @[MemPrimitives.scala 110:228:@34621.4]
  assign _T_2093 = _T_1882 & _T_1156; // @[MemPrimitives.scala 110:228:@34625.4]
  assign _T_2099 = _T_1888 & _T_1162; // @[MemPrimitives.scala 110:228:@34629.4]
  assign _T_2105 = _T_1894 & _T_1168; // @[MemPrimitives.scala 110:228:@34633.4]
  assign _T_2107 = StickySelects_22_io_outs_0; // @[MemPrimitives.scala 126:35:@34642.4]
  assign _T_2108 = StickySelects_22_io_outs_1; // @[MemPrimitives.scala 126:35:@34643.4]
  assign _T_2109 = StickySelects_22_io_outs_2; // @[MemPrimitives.scala 126:35:@34644.4]
  assign _T_2110 = StickySelects_22_io_outs_3; // @[MemPrimitives.scala 126:35:@34645.4]
  assign _T_2112 = {_T_2107,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@34647.4]
  assign _T_2114 = {_T_2108,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@34649.4]
  assign _T_2116 = {_T_2109,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@34651.4]
  assign _T_2118 = {_T_2110,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@34653.4]
  assign _T_2119 = _T_2109 ? _T_2116 : _T_2118; // @[Mux.scala 31:69:@34654.4]
  assign _T_2120 = _T_2108 ? _T_2114 : _T_2119; // @[Mux.scala 31:69:@34655.4]
  assign _T_2121 = _T_2107 ? _T_2112 : _T_2120; // @[Mux.scala 31:69:@34656.4]
  assign _T_2129 = _T_1918 & _T_1192; // @[MemPrimitives.scala 110:228:@34665.4]
  assign _T_2135 = _T_1924 & _T_1198; // @[MemPrimitives.scala 110:228:@34669.4]
  assign _T_2141 = _T_1930 & _T_1204; // @[MemPrimitives.scala 110:228:@34673.4]
  assign _T_2147 = _T_1936 & _T_1210; // @[MemPrimitives.scala 110:228:@34677.4]
  assign _T_2153 = _T_1942 & _T_1216; // @[MemPrimitives.scala 110:228:@34681.4]
  assign _T_2159 = _T_1948 & _T_1222; // @[MemPrimitives.scala 110:228:@34685.4]
  assign _T_2161 = StickySelects_23_io_outs_0; // @[MemPrimitives.scala 126:35:@34696.4]
  assign _T_2162 = StickySelects_23_io_outs_1; // @[MemPrimitives.scala 126:35:@34697.4]
  assign _T_2163 = StickySelects_23_io_outs_2; // @[MemPrimitives.scala 126:35:@34698.4]
  assign _T_2164 = StickySelects_23_io_outs_3; // @[MemPrimitives.scala 126:35:@34699.4]
  assign _T_2165 = StickySelects_23_io_outs_4; // @[MemPrimitives.scala 126:35:@34700.4]
  assign _T_2166 = StickySelects_23_io_outs_5; // @[MemPrimitives.scala 126:35:@34701.4]
  assign _T_2168 = {_T_2161,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@34703.4]
  assign _T_2170 = {_T_2162,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@34705.4]
  assign _T_2172 = {_T_2163,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@34707.4]
  assign _T_2174 = {_T_2164,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@34709.4]
  assign _T_2176 = {_T_2165,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@34711.4]
  assign _T_2178 = {_T_2166,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@34713.4]
  assign _T_2179 = _T_2165 ? _T_2176 : _T_2178; // @[Mux.scala 31:69:@34714.4]
  assign _T_2180 = _T_2164 ? _T_2174 : _T_2179; // @[Mux.scala 31:69:@34715.4]
  assign _T_2181 = _T_2163 ? _T_2172 : _T_2180; // @[Mux.scala 31:69:@34716.4]
  assign _T_2182 = _T_2162 ? _T_2170 : _T_2181; // @[Mux.scala 31:69:@34717.4]
  assign _T_2183 = _T_2161 ? _T_2168 : _T_2182; // @[Mux.scala 31:69:@34718.4]
  assign _T_2279 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@34847.4 package.scala 96:25:@34848.4]
  assign _T_2283 = _T_2279 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@34857.4]
  assign _T_2276 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@34839.4 package.scala 96:25:@34840.4]
  assign _T_2284 = _T_2276 ? Mem1D_19_io_output : _T_2283; // @[Mux.scala 31:69:@34858.4]
  assign _T_2273 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@34831.4 package.scala 96:25:@34832.4]
  assign _T_2285 = _T_2273 ? Mem1D_17_io_output : _T_2284; // @[Mux.scala 31:69:@34859.4]
  assign _T_2270 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@34823.4 package.scala 96:25:@34824.4]
  assign _T_2286 = _T_2270 ? Mem1D_15_io_output : _T_2285; // @[Mux.scala 31:69:@34860.4]
  assign _T_2267 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@34815.4 package.scala 96:25:@34816.4]
  assign _T_2287 = _T_2267 ? Mem1D_13_io_output : _T_2286; // @[Mux.scala 31:69:@34861.4]
  assign _T_2264 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@34807.4 package.scala 96:25:@34808.4]
  assign _T_2288 = _T_2264 ? Mem1D_11_io_output : _T_2287; // @[Mux.scala 31:69:@34862.4]
  assign _T_2261 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@34799.4 package.scala 96:25:@34800.4]
  assign _T_2289 = _T_2261 ? Mem1D_9_io_output : _T_2288; // @[Mux.scala 31:69:@34863.4]
  assign _T_2258 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@34791.4 package.scala 96:25:@34792.4]
  assign _T_2290 = _T_2258 ? Mem1D_7_io_output : _T_2289; // @[Mux.scala 31:69:@34864.4]
  assign _T_2255 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@34783.4 package.scala 96:25:@34784.4]
  assign _T_2291 = _T_2255 ? Mem1D_5_io_output : _T_2290; // @[Mux.scala 31:69:@34865.4]
  assign _T_2252 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@34775.4 package.scala 96:25:@34776.4]
  assign _T_2292 = _T_2252 ? Mem1D_3_io_output : _T_2291; // @[Mux.scala 31:69:@34866.4]
  assign _T_2249 = RetimeWrapper_io_out; // @[package.scala 96:25:@34767.4 package.scala 96:25:@34768.4]
  assign _T_2386 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@34991.4 package.scala 96:25:@34992.4]
  assign _T_2390 = _T_2386 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@35001.4]
  assign _T_2383 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@34983.4 package.scala 96:25:@34984.4]
  assign _T_2391 = _T_2383 ? Mem1D_19_io_output : _T_2390; // @[Mux.scala 31:69:@35002.4]
  assign _T_2380 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@34975.4 package.scala 96:25:@34976.4]
  assign _T_2392 = _T_2380 ? Mem1D_17_io_output : _T_2391; // @[Mux.scala 31:69:@35003.4]
  assign _T_2377 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@34967.4 package.scala 96:25:@34968.4]
  assign _T_2393 = _T_2377 ? Mem1D_15_io_output : _T_2392; // @[Mux.scala 31:69:@35004.4]
  assign _T_2374 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@34959.4 package.scala 96:25:@34960.4]
  assign _T_2394 = _T_2374 ? Mem1D_13_io_output : _T_2393; // @[Mux.scala 31:69:@35005.4]
  assign _T_2371 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@34951.4 package.scala 96:25:@34952.4]
  assign _T_2395 = _T_2371 ? Mem1D_11_io_output : _T_2394; // @[Mux.scala 31:69:@35006.4]
  assign _T_2368 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@34943.4 package.scala 96:25:@34944.4]
  assign _T_2396 = _T_2368 ? Mem1D_9_io_output : _T_2395; // @[Mux.scala 31:69:@35007.4]
  assign _T_2365 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@34935.4 package.scala 96:25:@34936.4]
  assign _T_2397 = _T_2365 ? Mem1D_7_io_output : _T_2396; // @[Mux.scala 31:69:@35008.4]
  assign _T_2362 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@34927.4 package.scala 96:25:@34928.4]
  assign _T_2398 = _T_2362 ? Mem1D_5_io_output : _T_2397; // @[Mux.scala 31:69:@35009.4]
  assign _T_2359 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@34919.4 package.scala 96:25:@34920.4]
  assign _T_2399 = _T_2359 ? Mem1D_3_io_output : _T_2398; // @[Mux.scala 31:69:@35010.4]
  assign _T_2356 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@34911.4 package.scala 96:25:@34912.4]
  assign _T_2493 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@35135.4 package.scala 96:25:@35136.4]
  assign _T_2497 = _T_2493 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@35145.4]
  assign _T_2490 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@35127.4 package.scala 96:25:@35128.4]
  assign _T_2498 = _T_2490 ? Mem1D_19_io_output : _T_2497; // @[Mux.scala 31:69:@35146.4]
  assign _T_2487 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@35119.4 package.scala 96:25:@35120.4]
  assign _T_2499 = _T_2487 ? Mem1D_17_io_output : _T_2498; // @[Mux.scala 31:69:@35147.4]
  assign _T_2484 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@35111.4 package.scala 96:25:@35112.4]
  assign _T_2500 = _T_2484 ? Mem1D_15_io_output : _T_2499; // @[Mux.scala 31:69:@35148.4]
  assign _T_2481 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@35103.4 package.scala 96:25:@35104.4]
  assign _T_2501 = _T_2481 ? Mem1D_13_io_output : _T_2500; // @[Mux.scala 31:69:@35149.4]
  assign _T_2478 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@35095.4 package.scala 96:25:@35096.4]
  assign _T_2502 = _T_2478 ? Mem1D_11_io_output : _T_2501; // @[Mux.scala 31:69:@35150.4]
  assign _T_2475 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@35087.4 package.scala 96:25:@35088.4]
  assign _T_2503 = _T_2475 ? Mem1D_9_io_output : _T_2502; // @[Mux.scala 31:69:@35151.4]
  assign _T_2472 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@35079.4 package.scala 96:25:@35080.4]
  assign _T_2504 = _T_2472 ? Mem1D_7_io_output : _T_2503; // @[Mux.scala 31:69:@35152.4]
  assign _T_2469 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@35071.4 package.scala 96:25:@35072.4]
  assign _T_2505 = _T_2469 ? Mem1D_5_io_output : _T_2504; // @[Mux.scala 31:69:@35153.4]
  assign _T_2466 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@35063.4 package.scala 96:25:@35064.4]
  assign _T_2506 = _T_2466 ? Mem1D_3_io_output : _T_2505; // @[Mux.scala 31:69:@35154.4]
  assign _T_2463 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@35055.4 package.scala 96:25:@35056.4]
  assign _T_2600 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@35279.4 package.scala 96:25:@35280.4]
  assign _T_2604 = _T_2600 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@35289.4]
  assign _T_2597 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@35271.4 package.scala 96:25:@35272.4]
  assign _T_2605 = _T_2597 ? Mem1D_19_io_output : _T_2604; // @[Mux.scala 31:69:@35290.4]
  assign _T_2594 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@35263.4 package.scala 96:25:@35264.4]
  assign _T_2606 = _T_2594 ? Mem1D_17_io_output : _T_2605; // @[Mux.scala 31:69:@35291.4]
  assign _T_2591 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@35255.4 package.scala 96:25:@35256.4]
  assign _T_2607 = _T_2591 ? Mem1D_15_io_output : _T_2606; // @[Mux.scala 31:69:@35292.4]
  assign _T_2588 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@35247.4 package.scala 96:25:@35248.4]
  assign _T_2608 = _T_2588 ? Mem1D_13_io_output : _T_2607; // @[Mux.scala 31:69:@35293.4]
  assign _T_2585 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@35239.4 package.scala 96:25:@35240.4]
  assign _T_2609 = _T_2585 ? Mem1D_11_io_output : _T_2608; // @[Mux.scala 31:69:@35294.4]
  assign _T_2582 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@35231.4 package.scala 96:25:@35232.4]
  assign _T_2610 = _T_2582 ? Mem1D_9_io_output : _T_2609; // @[Mux.scala 31:69:@35295.4]
  assign _T_2579 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@35223.4 package.scala 96:25:@35224.4]
  assign _T_2611 = _T_2579 ? Mem1D_7_io_output : _T_2610; // @[Mux.scala 31:69:@35296.4]
  assign _T_2576 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@35215.4 package.scala 96:25:@35216.4]
  assign _T_2612 = _T_2576 ? Mem1D_5_io_output : _T_2611; // @[Mux.scala 31:69:@35297.4]
  assign _T_2573 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@35207.4 package.scala 96:25:@35208.4]
  assign _T_2613 = _T_2573 ? Mem1D_3_io_output : _T_2612; // @[Mux.scala 31:69:@35298.4]
  assign _T_2570 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@35199.4 package.scala 96:25:@35200.4]
  assign _T_2707 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@35423.4 package.scala 96:25:@35424.4]
  assign _T_2711 = _T_2707 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@35433.4]
  assign _T_2704 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@35415.4 package.scala 96:25:@35416.4]
  assign _T_2712 = _T_2704 ? Mem1D_18_io_output : _T_2711; // @[Mux.scala 31:69:@35434.4]
  assign _T_2701 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@35407.4 package.scala 96:25:@35408.4]
  assign _T_2713 = _T_2701 ? Mem1D_16_io_output : _T_2712; // @[Mux.scala 31:69:@35435.4]
  assign _T_2698 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@35399.4 package.scala 96:25:@35400.4]
  assign _T_2714 = _T_2698 ? Mem1D_14_io_output : _T_2713; // @[Mux.scala 31:69:@35436.4]
  assign _T_2695 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@35391.4 package.scala 96:25:@35392.4]
  assign _T_2715 = _T_2695 ? Mem1D_12_io_output : _T_2714; // @[Mux.scala 31:69:@35437.4]
  assign _T_2692 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@35383.4 package.scala 96:25:@35384.4]
  assign _T_2716 = _T_2692 ? Mem1D_10_io_output : _T_2715; // @[Mux.scala 31:69:@35438.4]
  assign _T_2689 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@35375.4 package.scala 96:25:@35376.4]
  assign _T_2717 = _T_2689 ? Mem1D_8_io_output : _T_2716; // @[Mux.scala 31:69:@35439.4]
  assign _T_2686 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@35367.4 package.scala 96:25:@35368.4]
  assign _T_2718 = _T_2686 ? Mem1D_6_io_output : _T_2717; // @[Mux.scala 31:69:@35440.4]
  assign _T_2683 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@35359.4 package.scala 96:25:@35360.4]
  assign _T_2719 = _T_2683 ? Mem1D_4_io_output : _T_2718; // @[Mux.scala 31:69:@35441.4]
  assign _T_2680 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@35351.4 package.scala 96:25:@35352.4]
  assign _T_2720 = _T_2680 ? Mem1D_2_io_output : _T_2719; // @[Mux.scala 31:69:@35442.4]
  assign _T_2677 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@35343.4 package.scala 96:25:@35344.4]
  assign _T_2814 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@35567.4 package.scala 96:25:@35568.4]
  assign _T_2818 = _T_2814 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@35577.4]
  assign _T_2811 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@35559.4 package.scala 96:25:@35560.4]
  assign _T_2819 = _T_2811 ? Mem1D_19_io_output : _T_2818; // @[Mux.scala 31:69:@35578.4]
  assign _T_2808 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@35551.4 package.scala 96:25:@35552.4]
  assign _T_2820 = _T_2808 ? Mem1D_17_io_output : _T_2819; // @[Mux.scala 31:69:@35579.4]
  assign _T_2805 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@35543.4 package.scala 96:25:@35544.4]
  assign _T_2821 = _T_2805 ? Mem1D_15_io_output : _T_2820; // @[Mux.scala 31:69:@35580.4]
  assign _T_2802 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@35535.4 package.scala 96:25:@35536.4]
  assign _T_2822 = _T_2802 ? Mem1D_13_io_output : _T_2821; // @[Mux.scala 31:69:@35581.4]
  assign _T_2799 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@35527.4 package.scala 96:25:@35528.4]
  assign _T_2823 = _T_2799 ? Mem1D_11_io_output : _T_2822; // @[Mux.scala 31:69:@35582.4]
  assign _T_2796 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@35519.4 package.scala 96:25:@35520.4]
  assign _T_2824 = _T_2796 ? Mem1D_9_io_output : _T_2823; // @[Mux.scala 31:69:@35583.4]
  assign _T_2793 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@35511.4 package.scala 96:25:@35512.4]
  assign _T_2825 = _T_2793 ? Mem1D_7_io_output : _T_2824; // @[Mux.scala 31:69:@35584.4]
  assign _T_2790 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@35503.4 package.scala 96:25:@35504.4]
  assign _T_2826 = _T_2790 ? Mem1D_5_io_output : _T_2825; // @[Mux.scala 31:69:@35585.4]
  assign _T_2787 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@35495.4 package.scala 96:25:@35496.4]
  assign _T_2827 = _T_2787 ? Mem1D_3_io_output : _T_2826; // @[Mux.scala 31:69:@35586.4]
  assign _T_2784 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@35487.4 package.scala 96:25:@35488.4]
  assign _T_2921 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@35711.4 package.scala 96:25:@35712.4]
  assign _T_2925 = _T_2921 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@35721.4]
  assign _T_2918 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@35703.4 package.scala 96:25:@35704.4]
  assign _T_2926 = _T_2918 ? Mem1D_18_io_output : _T_2925; // @[Mux.scala 31:69:@35722.4]
  assign _T_2915 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@35695.4 package.scala 96:25:@35696.4]
  assign _T_2927 = _T_2915 ? Mem1D_16_io_output : _T_2926; // @[Mux.scala 31:69:@35723.4]
  assign _T_2912 = RetimeWrapper_79_io_out; // @[package.scala 96:25:@35687.4 package.scala 96:25:@35688.4]
  assign _T_2928 = _T_2912 ? Mem1D_14_io_output : _T_2927; // @[Mux.scala 31:69:@35724.4]
  assign _T_2909 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@35679.4 package.scala 96:25:@35680.4]
  assign _T_2929 = _T_2909 ? Mem1D_12_io_output : _T_2928; // @[Mux.scala 31:69:@35725.4]
  assign _T_2906 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@35671.4 package.scala 96:25:@35672.4]
  assign _T_2930 = _T_2906 ? Mem1D_10_io_output : _T_2929; // @[Mux.scala 31:69:@35726.4]
  assign _T_2903 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@35663.4 package.scala 96:25:@35664.4]
  assign _T_2931 = _T_2903 ? Mem1D_8_io_output : _T_2930; // @[Mux.scala 31:69:@35727.4]
  assign _T_2900 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@35655.4 package.scala 96:25:@35656.4]
  assign _T_2932 = _T_2900 ? Mem1D_6_io_output : _T_2931; // @[Mux.scala 31:69:@35728.4]
  assign _T_2897 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@35647.4 package.scala 96:25:@35648.4]
  assign _T_2933 = _T_2897 ? Mem1D_4_io_output : _T_2932; // @[Mux.scala 31:69:@35729.4]
  assign _T_2894 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@35639.4 package.scala 96:25:@35640.4]
  assign _T_2934 = _T_2894 ? Mem1D_2_io_output : _T_2933; // @[Mux.scala 31:69:@35730.4]
  assign _T_2891 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@35631.4 package.scala 96:25:@35632.4]
  assign _T_3028 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@35855.4 package.scala 96:25:@35856.4]
  assign _T_3032 = _T_3028 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@35865.4]
  assign _T_3025 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@35847.4 package.scala 96:25:@35848.4]
  assign _T_3033 = _T_3025 ? Mem1D_18_io_output : _T_3032; // @[Mux.scala 31:69:@35866.4]
  assign _T_3022 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@35839.4 package.scala 96:25:@35840.4]
  assign _T_3034 = _T_3022 ? Mem1D_16_io_output : _T_3033; // @[Mux.scala 31:69:@35867.4]
  assign _T_3019 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@35831.4 package.scala 96:25:@35832.4]
  assign _T_3035 = _T_3019 ? Mem1D_14_io_output : _T_3034; // @[Mux.scala 31:69:@35868.4]
  assign _T_3016 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@35823.4 package.scala 96:25:@35824.4]
  assign _T_3036 = _T_3016 ? Mem1D_12_io_output : _T_3035; // @[Mux.scala 31:69:@35869.4]
  assign _T_3013 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@35815.4 package.scala 96:25:@35816.4]
  assign _T_3037 = _T_3013 ? Mem1D_10_io_output : _T_3036; // @[Mux.scala 31:69:@35870.4]
  assign _T_3010 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@35807.4 package.scala 96:25:@35808.4]
  assign _T_3038 = _T_3010 ? Mem1D_8_io_output : _T_3037; // @[Mux.scala 31:69:@35871.4]
  assign _T_3007 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@35799.4 package.scala 96:25:@35800.4]
  assign _T_3039 = _T_3007 ? Mem1D_6_io_output : _T_3038; // @[Mux.scala 31:69:@35872.4]
  assign _T_3004 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@35791.4 package.scala 96:25:@35792.4]
  assign _T_3040 = _T_3004 ? Mem1D_4_io_output : _T_3039; // @[Mux.scala 31:69:@35873.4]
  assign _T_3001 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@35783.4 package.scala 96:25:@35784.4]
  assign _T_3041 = _T_3001 ? Mem1D_2_io_output : _T_3040; // @[Mux.scala 31:69:@35874.4]
  assign _T_2998 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@35775.4 package.scala 96:25:@35776.4]
  assign _T_3135 = RetimeWrapper_106_io_out; // @[package.scala 96:25:@35999.4 package.scala 96:25:@36000.4]
  assign _T_3139 = _T_3135 ? Mem1D_21_io_output : Mem1D_23_io_output; // @[Mux.scala 31:69:@36009.4]
  assign _T_3132 = RetimeWrapper_105_io_out; // @[package.scala 96:25:@35991.4 package.scala 96:25:@35992.4]
  assign _T_3140 = _T_3132 ? Mem1D_19_io_output : _T_3139; // @[Mux.scala 31:69:@36010.4]
  assign _T_3129 = RetimeWrapper_104_io_out; // @[package.scala 96:25:@35983.4 package.scala 96:25:@35984.4]
  assign _T_3141 = _T_3129 ? Mem1D_17_io_output : _T_3140; // @[Mux.scala 31:69:@36011.4]
  assign _T_3126 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@35975.4 package.scala 96:25:@35976.4]
  assign _T_3142 = _T_3126 ? Mem1D_15_io_output : _T_3141; // @[Mux.scala 31:69:@36012.4]
  assign _T_3123 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@35967.4 package.scala 96:25:@35968.4]
  assign _T_3143 = _T_3123 ? Mem1D_13_io_output : _T_3142; // @[Mux.scala 31:69:@36013.4]
  assign _T_3120 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@35959.4 package.scala 96:25:@35960.4]
  assign _T_3144 = _T_3120 ? Mem1D_11_io_output : _T_3143; // @[Mux.scala 31:69:@36014.4]
  assign _T_3117 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@35951.4 package.scala 96:25:@35952.4]
  assign _T_3145 = _T_3117 ? Mem1D_9_io_output : _T_3144; // @[Mux.scala 31:69:@36015.4]
  assign _T_3114 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@35943.4 package.scala 96:25:@35944.4]
  assign _T_3146 = _T_3114 ? Mem1D_7_io_output : _T_3145; // @[Mux.scala 31:69:@36016.4]
  assign _T_3111 = RetimeWrapper_98_io_out; // @[package.scala 96:25:@35935.4 package.scala 96:25:@35936.4]
  assign _T_3147 = _T_3111 ? Mem1D_5_io_output : _T_3146; // @[Mux.scala 31:69:@36017.4]
  assign _T_3108 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@35927.4 package.scala 96:25:@35928.4]
  assign _T_3148 = _T_3108 ? Mem1D_3_io_output : _T_3147; // @[Mux.scala 31:69:@36018.4]
  assign _T_3105 = RetimeWrapper_96_io_out; // @[package.scala 96:25:@35919.4 package.scala 96:25:@35920.4]
  assign _T_3242 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@36143.4 package.scala 96:25:@36144.4]
  assign _T_3246 = _T_3242 ? Mem1D_20_io_output : Mem1D_22_io_output; // @[Mux.scala 31:69:@36153.4]
  assign _T_3239 = RetimeWrapper_117_io_out; // @[package.scala 96:25:@36135.4 package.scala 96:25:@36136.4]
  assign _T_3247 = _T_3239 ? Mem1D_18_io_output : _T_3246; // @[Mux.scala 31:69:@36154.4]
  assign _T_3236 = RetimeWrapper_116_io_out; // @[package.scala 96:25:@36127.4 package.scala 96:25:@36128.4]
  assign _T_3248 = _T_3236 ? Mem1D_16_io_output : _T_3247; // @[Mux.scala 31:69:@36155.4]
  assign _T_3233 = RetimeWrapper_115_io_out; // @[package.scala 96:25:@36119.4 package.scala 96:25:@36120.4]
  assign _T_3249 = _T_3233 ? Mem1D_14_io_output : _T_3248; // @[Mux.scala 31:69:@36156.4]
  assign _T_3230 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@36111.4 package.scala 96:25:@36112.4]
  assign _T_3250 = _T_3230 ? Mem1D_12_io_output : _T_3249; // @[Mux.scala 31:69:@36157.4]
  assign _T_3227 = RetimeWrapper_113_io_out; // @[package.scala 96:25:@36103.4 package.scala 96:25:@36104.4]
  assign _T_3251 = _T_3227 ? Mem1D_10_io_output : _T_3250; // @[Mux.scala 31:69:@36158.4]
  assign _T_3224 = RetimeWrapper_112_io_out; // @[package.scala 96:25:@36095.4 package.scala 96:25:@36096.4]
  assign _T_3252 = _T_3224 ? Mem1D_8_io_output : _T_3251; // @[Mux.scala 31:69:@36159.4]
  assign _T_3221 = RetimeWrapper_111_io_out; // @[package.scala 96:25:@36087.4 package.scala 96:25:@36088.4]
  assign _T_3253 = _T_3221 ? Mem1D_6_io_output : _T_3252; // @[Mux.scala 31:69:@36160.4]
  assign _T_3218 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@36079.4 package.scala 96:25:@36080.4]
  assign _T_3254 = _T_3218 ? Mem1D_4_io_output : _T_3253; // @[Mux.scala 31:69:@36161.4]
  assign _T_3215 = RetimeWrapper_109_io_out; // @[package.scala 96:25:@36071.4 package.scala 96:25:@36072.4]
  assign _T_3255 = _T_3215 ? Mem1D_2_io_output : _T_3254; // @[Mux.scala 31:69:@36162.4]
  assign _T_3212 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@36063.4 package.scala 96:25:@36064.4]
  assign io_rPort_9_output_0 = _T_3212 ? Mem1D_io_output : _T_3255; // @[MemPrimitives.scala 152:13:@36164.4]
  assign io_rPort_8_output_0 = _T_3105 ? Mem1D_1_io_output : _T_3148; // @[MemPrimitives.scala 152:13:@36020.4]
  assign io_rPort_7_output_0 = _T_2998 ? Mem1D_io_output : _T_3041; // @[MemPrimitives.scala 152:13:@35876.4]
  assign io_rPort_6_output_0 = _T_2891 ? Mem1D_io_output : _T_2934; // @[MemPrimitives.scala 152:13:@35732.4]
  assign io_rPort_5_output_0 = _T_2784 ? Mem1D_1_io_output : _T_2827; // @[MemPrimitives.scala 152:13:@35588.4]
  assign io_rPort_4_output_0 = _T_2677 ? Mem1D_io_output : _T_2720; // @[MemPrimitives.scala 152:13:@35444.4]
  assign io_rPort_3_output_0 = _T_2570 ? Mem1D_1_io_output : _T_2613; // @[MemPrimitives.scala 152:13:@35300.4]
  assign io_rPort_2_output_0 = _T_2463 ? Mem1D_1_io_output : _T_2506; // @[MemPrimitives.scala 152:13:@35156.4]
  assign io_rPort_1_output_0 = _T_2356 ? Mem1D_1_io_output : _T_2399; // @[MemPrimitives.scala 152:13:@35012.4]
  assign io_rPort_0_output_0 = _T_2249 ? Mem1D_1_io_output : _T_2292; // @[MemPrimitives.scala 152:13:@34868.4]
  assign Mem1D_clock = clock; // @[:@32614.4]
  assign Mem1D_reset = reset; // @[:@32615.4]
  assign Mem1D_io_r_ofs_0 = _T_977[8:0]; // @[MemPrimitives.scala 131:28:@33494.4]
  assign Mem1D_io_r_backpressure = _T_977[9]; // @[MemPrimitives.scala 132:32:@33495.4]
  assign Mem1D_io_w_ofs_0 = _T_475[8:0]; // @[MemPrimitives.scala 94:28:@33013.4]
  assign Mem1D_io_w_data_0 = _T_475[40:9]; // @[MemPrimitives.scala 95:29:@33014.4]
  assign Mem1D_io_w_en_0 = _T_475[41]; // @[MemPrimitives.scala 96:27:@33015.4]
  assign Mem1D_1_clock = clock; // @[:@32630.4]
  assign Mem1D_1_reset = reset; // @[:@32631.4]
  assign Mem1D_1_io_r_ofs_0 = _T_1039[8:0]; // @[MemPrimitives.scala 131:28:@33556.4]
  assign Mem1D_1_io_r_backpressure = _T_1039[9]; // @[MemPrimitives.scala 132:32:@33557.4]
  assign Mem1D_1_io_w_ofs_0 = _T_495[8:0]; // @[MemPrimitives.scala 94:28:@33032.4]
  assign Mem1D_1_io_w_data_0 = _T_495[40:9]; // @[MemPrimitives.scala 95:29:@33033.4]
  assign Mem1D_1_io_w_en_0 = _T_495[41]; // @[MemPrimitives.scala 96:27:@33034.4]
  assign Mem1D_2_clock = clock; // @[:@32646.4]
  assign Mem1D_2_reset = reset; // @[:@32647.4]
  assign Mem1D_2_io_r_ofs_0 = _T_1081[8:0]; // @[MemPrimitives.scala 131:28:@33600.4]
  assign Mem1D_2_io_r_backpressure = _T_1081[9]; // @[MemPrimitives.scala 132:32:@33601.4]
  assign Mem1D_2_io_w_ofs_0 = _T_515[8:0]; // @[MemPrimitives.scala 94:28:@33051.4]
  assign Mem1D_2_io_w_data_0 = _T_515[40:9]; // @[MemPrimitives.scala 95:29:@33052.4]
  assign Mem1D_2_io_w_en_0 = _T_515[41]; // @[MemPrimitives.scala 96:27:@33053.4]
  assign Mem1D_3_clock = clock; // @[:@32662.4]
  assign Mem1D_3_reset = reset; // @[:@32663.4]
  assign Mem1D_3_io_r_ofs_0 = _T_1143[8:0]; // @[MemPrimitives.scala 131:28:@33662.4]
  assign Mem1D_3_io_r_backpressure = _T_1143[9]; // @[MemPrimitives.scala 132:32:@33663.4]
  assign Mem1D_3_io_w_ofs_0 = _T_535[8:0]; // @[MemPrimitives.scala 94:28:@33070.4]
  assign Mem1D_3_io_w_data_0 = _T_535[40:9]; // @[MemPrimitives.scala 95:29:@33071.4]
  assign Mem1D_3_io_w_en_0 = _T_535[41]; // @[MemPrimitives.scala 96:27:@33072.4]
  assign Mem1D_4_clock = clock; // @[:@32678.4]
  assign Mem1D_4_reset = reset; // @[:@32679.4]
  assign Mem1D_4_io_r_ofs_0 = _T_1185[8:0]; // @[MemPrimitives.scala 131:28:@33706.4]
  assign Mem1D_4_io_r_backpressure = _T_1185[9]; // @[MemPrimitives.scala 132:32:@33707.4]
  assign Mem1D_4_io_w_ofs_0 = _T_555[8:0]; // @[MemPrimitives.scala 94:28:@33089.4]
  assign Mem1D_4_io_w_data_0 = _T_555[40:9]; // @[MemPrimitives.scala 95:29:@33090.4]
  assign Mem1D_4_io_w_en_0 = _T_555[41]; // @[MemPrimitives.scala 96:27:@33091.4]
  assign Mem1D_5_clock = clock; // @[:@32694.4]
  assign Mem1D_5_reset = reset; // @[:@32695.4]
  assign Mem1D_5_io_r_ofs_0 = _T_1247[8:0]; // @[MemPrimitives.scala 131:28:@33768.4]
  assign Mem1D_5_io_r_backpressure = _T_1247[9]; // @[MemPrimitives.scala 132:32:@33769.4]
  assign Mem1D_5_io_w_ofs_0 = _T_575[8:0]; // @[MemPrimitives.scala 94:28:@33108.4]
  assign Mem1D_5_io_w_data_0 = _T_575[40:9]; // @[MemPrimitives.scala 95:29:@33109.4]
  assign Mem1D_5_io_w_en_0 = _T_575[41]; // @[MemPrimitives.scala 96:27:@33110.4]
  assign Mem1D_6_clock = clock; // @[:@32710.4]
  assign Mem1D_6_reset = reset; // @[:@32711.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1289[8:0]; // @[MemPrimitives.scala 131:28:@33812.4]
  assign Mem1D_6_io_r_backpressure = _T_1289[9]; // @[MemPrimitives.scala 132:32:@33813.4]
  assign Mem1D_6_io_w_ofs_0 = _T_595[8:0]; // @[MemPrimitives.scala 94:28:@33127.4]
  assign Mem1D_6_io_w_data_0 = _T_595[40:9]; // @[MemPrimitives.scala 95:29:@33128.4]
  assign Mem1D_6_io_w_en_0 = _T_595[41]; // @[MemPrimitives.scala 96:27:@33129.4]
  assign Mem1D_7_clock = clock; // @[:@32726.4]
  assign Mem1D_7_reset = reset; // @[:@32727.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1351[8:0]; // @[MemPrimitives.scala 131:28:@33874.4]
  assign Mem1D_7_io_r_backpressure = _T_1351[9]; // @[MemPrimitives.scala 132:32:@33875.4]
  assign Mem1D_7_io_w_ofs_0 = _T_615[8:0]; // @[MemPrimitives.scala 94:28:@33146.4]
  assign Mem1D_7_io_w_data_0 = _T_615[40:9]; // @[MemPrimitives.scala 95:29:@33147.4]
  assign Mem1D_7_io_w_en_0 = _T_615[41]; // @[MemPrimitives.scala 96:27:@33148.4]
  assign Mem1D_8_clock = clock; // @[:@32742.4]
  assign Mem1D_8_reset = reset; // @[:@32743.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1393[8:0]; // @[MemPrimitives.scala 131:28:@33918.4]
  assign Mem1D_8_io_r_backpressure = _T_1393[9]; // @[MemPrimitives.scala 132:32:@33919.4]
  assign Mem1D_8_io_w_ofs_0 = _T_635[8:0]; // @[MemPrimitives.scala 94:28:@33165.4]
  assign Mem1D_8_io_w_data_0 = _T_635[40:9]; // @[MemPrimitives.scala 95:29:@33166.4]
  assign Mem1D_8_io_w_en_0 = _T_635[41]; // @[MemPrimitives.scala 96:27:@33167.4]
  assign Mem1D_9_clock = clock; // @[:@32758.4]
  assign Mem1D_9_reset = reset; // @[:@32759.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1455[8:0]; // @[MemPrimitives.scala 131:28:@33980.4]
  assign Mem1D_9_io_r_backpressure = _T_1455[9]; // @[MemPrimitives.scala 132:32:@33981.4]
  assign Mem1D_9_io_w_ofs_0 = _T_655[8:0]; // @[MemPrimitives.scala 94:28:@33184.4]
  assign Mem1D_9_io_w_data_0 = _T_655[40:9]; // @[MemPrimitives.scala 95:29:@33185.4]
  assign Mem1D_9_io_w_en_0 = _T_655[41]; // @[MemPrimitives.scala 96:27:@33186.4]
  assign Mem1D_10_clock = clock; // @[:@32774.4]
  assign Mem1D_10_reset = reset; // @[:@32775.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1497[8:0]; // @[MemPrimitives.scala 131:28:@34024.4]
  assign Mem1D_10_io_r_backpressure = _T_1497[9]; // @[MemPrimitives.scala 132:32:@34025.4]
  assign Mem1D_10_io_w_ofs_0 = _T_675[8:0]; // @[MemPrimitives.scala 94:28:@33203.4]
  assign Mem1D_10_io_w_data_0 = _T_675[40:9]; // @[MemPrimitives.scala 95:29:@33204.4]
  assign Mem1D_10_io_w_en_0 = _T_675[41]; // @[MemPrimitives.scala 96:27:@33205.4]
  assign Mem1D_11_clock = clock; // @[:@32790.4]
  assign Mem1D_11_reset = reset; // @[:@32791.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1559[8:0]; // @[MemPrimitives.scala 131:28:@34086.4]
  assign Mem1D_11_io_r_backpressure = _T_1559[9]; // @[MemPrimitives.scala 132:32:@34087.4]
  assign Mem1D_11_io_w_ofs_0 = _T_695[8:0]; // @[MemPrimitives.scala 94:28:@33222.4]
  assign Mem1D_11_io_w_data_0 = _T_695[40:9]; // @[MemPrimitives.scala 95:29:@33223.4]
  assign Mem1D_11_io_w_en_0 = _T_695[41]; // @[MemPrimitives.scala 96:27:@33224.4]
  assign Mem1D_12_clock = clock; // @[:@32806.4]
  assign Mem1D_12_reset = reset; // @[:@32807.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1601[8:0]; // @[MemPrimitives.scala 131:28:@34130.4]
  assign Mem1D_12_io_r_backpressure = _T_1601[9]; // @[MemPrimitives.scala 132:32:@34131.4]
  assign Mem1D_12_io_w_ofs_0 = _T_715[8:0]; // @[MemPrimitives.scala 94:28:@33241.4]
  assign Mem1D_12_io_w_data_0 = _T_715[40:9]; // @[MemPrimitives.scala 95:29:@33242.4]
  assign Mem1D_12_io_w_en_0 = _T_715[41]; // @[MemPrimitives.scala 96:27:@33243.4]
  assign Mem1D_13_clock = clock; // @[:@32822.4]
  assign Mem1D_13_reset = reset; // @[:@32823.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1663[8:0]; // @[MemPrimitives.scala 131:28:@34192.4]
  assign Mem1D_13_io_r_backpressure = _T_1663[9]; // @[MemPrimitives.scala 132:32:@34193.4]
  assign Mem1D_13_io_w_ofs_0 = _T_735[8:0]; // @[MemPrimitives.scala 94:28:@33260.4]
  assign Mem1D_13_io_w_data_0 = _T_735[40:9]; // @[MemPrimitives.scala 95:29:@33261.4]
  assign Mem1D_13_io_w_en_0 = _T_735[41]; // @[MemPrimitives.scala 96:27:@33262.4]
  assign Mem1D_14_clock = clock; // @[:@32838.4]
  assign Mem1D_14_reset = reset; // @[:@32839.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1705[8:0]; // @[MemPrimitives.scala 131:28:@34236.4]
  assign Mem1D_14_io_r_backpressure = _T_1705[9]; // @[MemPrimitives.scala 132:32:@34237.4]
  assign Mem1D_14_io_w_ofs_0 = _T_755[8:0]; // @[MemPrimitives.scala 94:28:@33279.4]
  assign Mem1D_14_io_w_data_0 = _T_755[40:9]; // @[MemPrimitives.scala 95:29:@33280.4]
  assign Mem1D_14_io_w_en_0 = _T_755[41]; // @[MemPrimitives.scala 96:27:@33281.4]
  assign Mem1D_15_clock = clock; // @[:@32854.4]
  assign Mem1D_15_reset = reset; // @[:@32855.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1767[8:0]; // @[MemPrimitives.scala 131:28:@34298.4]
  assign Mem1D_15_io_r_backpressure = _T_1767[9]; // @[MemPrimitives.scala 132:32:@34299.4]
  assign Mem1D_15_io_w_ofs_0 = _T_775[8:0]; // @[MemPrimitives.scala 94:28:@33298.4]
  assign Mem1D_15_io_w_data_0 = _T_775[40:9]; // @[MemPrimitives.scala 95:29:@33299.4]
  assign Mem1D_15_io_w_en_0 = _T_775[41]; // @[MemPrimitives.scala 96:27:@33300.4]
  assign Mem1D_16_clock = clock; // @[:@32870.4]
  assign Mem1D_16_reset = reset; // @[:@32871.4]
  assign Mem1D_16_io_r_ofs_0 = _T_1809[8:0]; // @[MemPrimitives.scala 131:28:@34342.4]
  assign Mem1D_16_io_r_backpressure = _T_1809[9]; // @[MemPrimitives.scala 132:32:@34343.4]
  assign Mem1D_16_io_w_ofs_0 = _T_795[8:0]; // @[MemPrimitives.scala 94:28:@33317.4]
  assign Mem1D_16_io_w_data_0 = _T_795[40:9]; // @[MemPrimitives.scala 95:29:@33318.4]
  assign Mem1D_16_io_w_en_0 = _T_795[41]; // @[MemPrimitives.scala 96:27:@33319.4]
  assign Mem1D_17_clock = clock; // @[:@32886.4]
  assign Mem1D_17_reset = reset; // @[:@32887.4]
  assign Mem1D_17_io_r_ofs_0 = _T_1871[8:0]; // @[MemPrimitives.scala 131:28:@34404.4]
  assign Mem1D_17_io_r_backpressure = _T_1871[9]; // @[MemPrimitives.scala 132:32:@34405.4]
  assign Mem1D_17_io_w_ofs_0 = _T_815[8:0]; // @[MemPrimitives.scala 94:28:@33336.4]
  assign Mem1D_17_io_w_data_0 = _T_815[40:9]; // @[MemPrimitives.scala 95:29:@33337.4]
  assign Mem1D_17_io_w_en_0 = _T_815[41]; // @[MemPrimitives.scala 96:27:@33338.4]
  assign Mem1D_18_clock = clock; // @[:@32902.4]
  assign Mem1D_18_reset = reset; // @[:@32903.4]
  assign Mem1D_18_io_r_ofs_0 = _T_1913[8:0]; // @[MemPrimitives.scala 131:28:@34448.4]
  assign Mem1D_18_io_r_backpressure = _T_1913[9]; // @[MemPrimitives.scala 132:32:@34449.4]
  assign Mem1D_18_io_w_ofs_0 = _T_835[8:0]; // @[MemPrimitives.scala 94:28:@33355.4]
  assign Mem1D_18_io_w_data_0 = _T_835[40:9]; // @[MemPrimitives.scala 95:29:@33356.4]
  assign Mem1D_18_io_w_en_0 = _T_835[41]; // @[MemPrimitives.scala 96:27:@33357.4]
  assign Mem1D_19_clock = clock; // @[:@32918.4]
  assign Mem1D_19_reset = reset; // @[:@32919.4]
  assign Mem1D_19_io_r_ofs_0 = _T_1975[8:0]; // @[MemPrimitives.scala 131:28:@34510.4]
  assign Mem1D_19_io_r_backpressure = _T_1975[9]; // @[MemPrimitives.scala 132:32:@34511.4]
  assign Mem1D_19_io_w_ofs_0 = _T_855[8:0]; // @[MemPrimitives.scala 94:28:@33374.4]
  assign Mem1D_19_io_w_data_0 = _T_855[40:9]; // @[MemPrimitives.scala 95:29:@33375.4]
  assign Mem1D_19_io_w_en_0 = _T_855[41]; // @[MemPrimitives.scala 96:27:@33376.4]
  assign Mem1D_20_clock = clock; // @[:@32934.4]
  assign Mem1D_20_reset = reset; // @[:@32935.4]
  assign Mem1D_20_io_r_ofs_0 = _T_2017[8:0]; // @[MemPrimitives.scala 131:28:@34554.4]
  assign Mem1D_20_io_r_backpressure = _T_2017[9]; // @[MemPrimitives.scala 132:32:@34555.4]
  assign Mem1D_20_io_w_ofs_0 = _T_875[8:0]; // @[MemPrimitives.scala 94:28:@33393.4]
  assign Mem1D_20_io_w_data_0 = _T_875[40:9]; // @[MemPrimitives.scala 95:29:@33394.4]
  assign Mem1D_20_io_w_en_0 = _T_875[41]; // @[MemPrimitives.scala 96:27:@33395.4]
  assign Mem1D_21_clock = clock; // @[:@32950.4]
  assign Mem1D_21_reset = reset; // @[:@32951.4]
  assign Mem1D_21_io_r_ofs_0 = _T_2079[8:0]; // @[MemPrimitives.scala 131:28:@34616.4]
  assign Mem1D_21_io_r_backpressure = _T_2079[9]; // @[MemPrimitives.scala 132:32:@34617.4]
  assign Mem1D_21_io_w_ofs_0 = _T_895[8:0]; // @[MemPrimitives.scala 94:28:@33412.4]
  assign Mem1D_21_io_w_data_0 = _T_895[40:9]; // @[MemPrimitives.scala 95:29:@33413.4]
  assign Mem1D_21_io_w_en_0 = _T_895[41]; // @[MemPrimitives.scala 96:27:@33414.4]
  assign Mem1D_22_clock = clock; // @[:@32966.4]
  assign Mem1D_22_reset = reset; // @[:@32967.4]
  assign Mem1D_22_io_r_ofs_0 = _T_2121[8:0]; // @[MemPrimitives.scala 131:28:@34660.4]
  assign Mem1D_22_io_r_backpressure = _T_2121[9]; // @[MemPrimitives.scala 132:32:@34661.4]
  assign Mem1D_22_io_w_ofs_0 = _T_915[8:0]; // @[MemPrimitives.scala 94:28:@33431.4]
  assign Mem1D_22_io_w_data_0 = _T_915[40:9]; // @[MemPrimitives.scala 95:29:@33432.4]
  assign Mem1D_22_io_w_en_0 = _T_915[41]; // @[MemPrimitives.scala 96:27:@33433.4]
  assign Mem1D_23_clock = clock; // @[:@32982.4]
  assign Mem1D_23_reset = reset; // @[:@32983.4]
  assign Mem1D_23_io_r_ofs_0 = _T_2183[8:0]; // @[MemPrimitives.scala 131:28:@34722.4]
  assign Mem1D_23_io_r_backpressure = _T_2183[9]; // @[MemPrimitives.scala 132:32:@34723.4]
  assign Mem1D_23_io_w_ofs_0 = _T_935[8:0]; // @[MemPrimitives.scala 94:28:@33450.4]
  assign Mem1D_23_io_w_data_0 = _T_935[40:9]; // @[MemPrimitives.scala 95:29:@33451.4]
  assign Mem1D_23_io_w_en_0 = _T_935[41]; // @[MemPrimitives.scala 96:27:@33452.4]
  assign StickySelects_clock = clock; // @[:@33470.4]
  assign StickySelects_reset = reset; // @[:@33471.4]
  assign StickySelects_io_ins_0 = io_rPort_4_en_0 & _T_943; // @[MemPrimitives.scala 125:64:@33472.4]
  assign StickySelects_io_ins_1 = io_rPort_6_en_0 & _T_949; // @[MemPrimitives.scala 125:64:@33473.4]
  assign StickySelects_io_ins_2 = io_rPort_7_en_0 & _T_955; // @[MemPrimitives.scala 125:64:@33474.4]
  assign StickySelects_io_ins_3 = io_rPort_9_en_0 & _T_961; // @[MemPrimitives.scala 125:64:@33475.4]
  assign StickySelects_1_clock = clock; // @[:@33522.4]
  assign StickySelects_1_reset = reset; // @[:@33523.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_985; // @[MemPrimitives.scala 125:64:@33524.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_991; // @[MemPrimitives.scala 125:64:@33525.4]
  assign StickySelects_1_io_ins_2 = io_rPort_2_en_0 & _T_997; // @[MemPrimitives.scala 125:64:@33526.4]
  assign StickySelects_1_io_ins_3 = io_rPort_3_en_0 & _T_1003; // @[MemPrimitives.scala 125:64:@33527.4]
  assign StickySelects_1_io_ins_4 = io_rPort_5_en_0 & _T_1009; // @[MemPrimitives.scala 125:64:@33528.4]
  assign StickySelects_1_io_ins_5 = io_rPort_8_en_0 & _T_1015; // @[MemPrimitives.scala 125:64:@33529.4]
  assign StickySelects_2_clock = clock; // @[:@33576.4]
  assign StickySelects_2_reset = reset; // @[:@33577.4]
  assign StickySelects_2_io_ins_0 = io_rPort_4_en_0 & _T_1047; // @[MemPrimitives.scala 125:64:@33578.4]
  assign StickySelects_2_io_ins_1 = io_rPort_6_en_0 & _T_1053; // @[MemPrimitives.scala 125:64:@33579.4]
  assign StickySelects_2_io_ins_2 = io_rPort_7_en_0 & _T_1059; // @[MemPrimitives.scala 125:64:@33580.4]
  assign StickySelects_2_io_ins_3 = io_rPort_9_en_0 & _T_1065; // @[MemPrimitives.scala 125:64:@33581.4]
  assign StickySelects_3_clock = clock; // @[:@33628.4]
  assign StickySelects_3_reset = reset; // @[:@33629.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_1089; // @[MemPrimitives.scala 125:64:@33630.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_1095; // @[MemPrimitives.scala 125:64:@33631.4]
  assign StickySelects_3_io_ins_2 = io_rPort_2_en_0 & _T_1101; // @[MemPrimitives.scala 125:64:@33632.4]
  assign StickySelects_3_io_ins_3 = io_rPort_3_en_0 & _T_1107; // @[MemPrimitives.scala 125:64:@33633.4]
  assign StickySelects_3_io_ins_4 = io_rPort_5_en_0 & _T_1113; // @[MemPrimitives.scala 125:64:@33634.4]
  assign StickySelects_3_io_ins_5 = io_rPort_8_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@33635.4]
  assign StickySelects_4_clock = clock; // @[:@33682.4]
  assign StickySelects_4_reset = reset; // @[:@33683.4]
  assign StickySelects_4_io_ins_0 = io_rPort_4_en_0 & _T_1151; // @[MemPrimitives.scala 125:64:@33684.4]
  assign StickySelects_4_io_ins_1 = io_rPort_6_en_0 & _T_1157; // @[MemPrimitives.scala 125:64:@33685.4]
  assign StickySelects_4_io_ins_2 = io_rPort_7_en_0 & _T_1163; // @[MemPrimitives.scala 125:64:@33686.4]
  assign StickySelects_4_io_ins_3 = io_rPort_9_en_0 & _T_1169; // @[MemPrimitives.scala 125:64:@33687.4]
  assign StickySelects_5_clock = clock; // @[:@33734.4]
  assign StickySelects_5_reset = reset; // @[:@33735.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@33736.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@33737.4]
  assign StickySelects_5_io_ins_2 = io_rPort_2_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@33738.4]
  assign StickySelects_5_io_ins_3 = io_rPort_3_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@33739.4]
  assign StickySelects_5_io_ins_4 = io_rPort_5_en_0 & _T_1217; // @[MemPrimitives.scala 125:64:@33740.4]
  assign StickySelects_5_io_ins_5 = io_rPort_8_en_0 & _T_1223; // @[MemPrimitives.scala 125:64:@33741.4]
  assign StickySelects_6_clock = clock; // @[:@33788.4]
  assign StickySelects_6_reset = reset; // @[:@33789.4]
  assign StickySelects_6_io_ins_0 = io_rPort_4_en_0 & _T_1255; // @[MemPrimitives.scala 125:64:@33790.4]
  assign StickySelects_6_io_ins_1 = io_rPort_6_en_0 & _T_1261; // @[MemPrimitives.scala 125:64:@33791.4]
  assign StickySelects_6_io_ins_2 = io_rPort_7_en_0 & _T_1267; // @[MemPrimitives.scala 125:64:@33792.4]
  assign StickySelects_6_io_ins_3 = io_rPort_9_en_0 & _T_1273; // @[MemPrimitives.scala 125:64:@33793.4]
  assign StickySelects_7_clock = clock; // @[:@33840.4]
  assign StickySelects_7_reset = reset; // @[:@33841.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1297; // @[MemPrimitives.scala 125:64:@33842.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1303; // @[MemPrimitives.scala 125:64:@33843.4]
  assign StickySelects_7_io_ins_2 = io_rPort_2_en_0 & _T_1309; // @[MemPrimitives.scala 125:64:@33844.4]
  assign StickySelects_7_io_ins_3 = io_rPort_3_en_0 & _T_1315; // @[MemPrimitives.scala 125:64:@33845.4]
  assign StickySelects_7_io_ins_4 = io_rPort_5_en_0 & _T_1321; // @[MemPrimitives.scala 125:64:@33846.4]
  assign StickySelects_7_io_ins_5 = io_rPort_8_en_0 & _T_1327; // @[MemPrimitives.scala 125:64:@33847.4]
  assign StickySelects_8_clock = clock; // @[:@33894.4]
  assign StickySelects_8_reset = reset; // @[:@33895.4]
  assign StickySelects_8_io_ins_0 = io_rPort_4_en_0 & _T_1359; // @[MemPrimitives.scala 125:64:@33896.4]
  assign StickySelects_8_io_ins_1 = io_rPort_6_en_0 & _T_1365; // @[MemPrimitives.scala 125:64:@33897.4]
  assign StickySelects_8_io_ins_2 = io_rPort_7_en_0 & _T_1371; // @[MemPrimitives.scala 125:64:@33898.4]
  assign StickySelects_8_io_ins_3 = io_rPort_9_en_0 & _T_1377; // @[MemPrimitives.scala 125:64:@33899.4]
  assign StickySelects_9_clock = clock; // @[:@33946.4]
  assign StickySelects_9_reset = reset; // @[:@33947.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1401; // @[MemPrimitives.scala 125:64:@33948.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1407; // @[MemPrimitives.scala 125:64:@33949.4]
  assign StickySelects_9_io_ins_2 = io_rPort_2_en_0 & _T_1413; // @[MemPrimitives.scala 125:64:@33950.4]
  assign StickySelects_9_io_ins_3 = io_rPort_3_en_0 & _T_1419; // @[MemPrimitives.scala 125:64:@33951.4]
  assign StickySelects_9_io_ins_4 = io_rPort_5_en_0 & _T_1425; // @[MemPrimitives.scala 125:64:@33952.4]
  assign StickySelects_9_io_ins_5 = io_rPort_8_en_0 & _T_1431; // @[MemPrimitives.scala 125:64:@33953.4]
  assign StickySelects_10_clock = clock; // @[:@34000.4]
  assign StickySelects_10_reset = reset; // @[:@34001.4]
  assign StickySelects_10_io_ins_0 = io_rPort_4_en_0 & _T_1463; // @[MemPrimitives.scala 125:64:@34002.4]
  assign StickySelects_10_io_ins_1 = io_rPort_6_en_0 & _T_1469; // @[MemPrimitives.scala 125:64:@34003.4]
  assign StickySelects_10_io_ins_2 = io_rPort_7_en_0 & _T_1475; // @[MemPrimitives.scala 125:64:@34004.4]
  assign StickySelects_10_io_ins_3 = io_rPort_9_en_0 & _T_1481; // @[MemPrimitives.scala 125:64:@34005.4]
  assign StickySelects_11_clock = clock; // @[:@34052.4]
  assign StickySelects_11_reset = reset; // @[:@34053.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1505; // @[MemPrimitives.scala 125:64:@34054.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1511; // @[MemPrimitives.scala 125:64:@34055.4]
  assign StickySelects_11_io_ins_2 = io_rPort_2_en_0 & _T_1517; // @[MemPrimitives.scala 125:64:@34056.4]
  assign StickySelects_11_io_ins_3 = io_rPort_3_en_0 & _T_1523; // @[MemPrimitives.scala 125:64:@34057.4]
  assign StickySelects_11_io_ins_4 = io_rPort_5_en_0 & _T_1529; // @[MemPrimitives.scala 125:64:@34058.4]
  assign StickySelects_11_io_ins_5 = io_rPort_8_en_0 & _T_1535; // @[MemPrimitives.scala 125:64:@34059.4]
  assign StickySelects_12_clock = clock; // @[:@34106.4]
  assign StickySelects_12_reset = reset; // @[:@34107.4]
  assign StickySelects_12_io_ins_0 = io_rPort_4_en_0 & _T_1567; // @[MemPrimitives.scala 125:64:@34108.4]
  assign StickySelects_12_io_ins_1 = io_rPort_6_en_0 & _T_1573; // @[MemPrimitives.scala 125:64:@34109.4]
  assign StickySelects_12_io_ins_2 = io_rPort_7_en_0 & _T_1579; // @[MemPrimitives.scala 125:64:@34110.4]
  assign StickySelects_12_io_ins_3 = io_rPort_9_en_0 & _T_1585; // @[MemPrimitives.scala 125:64:@34111.4]
  assign StickySelects_13_clock = clock; // @[:@34158.4]
  assign StickySelects_13_reset = reset; // @[:@34159.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_1609; // @[MemPrimitives.scala 125:64:@34160.4]
  assign StickySelects_13_io_ins_1 = io_rPort_1_en_0 & _T_1615; // @[MemPrimitives.scala 125:64:@34161.4]
  assign StickySelects_13_io_ins_2 = io_rPort_2_en_0 & _T_1621; // @[MemPrimitives.scala 125:64:@34162.4]
  assign StickySelects_13_io_ins_3 = io_rPort_3_en_0 & _T_1627; // @[MemPrimitives.scala 125:64:@34163.4]
  assign StickySelects_13_io_ins_4 = io_rPort_5_en_0 & _T_1633; // @[MemPrimitives.scala 125:64:@34164.4]
  assign StickySelects_13_io_ins_5 = io_rPort_8_en_0 & _T_1639; // @[MemPrimitives.scala 125:64:@34165.4]
  assign StickySelects_14_clock = clock; // @[:@34212.4]
  assign StickySelects_14_reset = reset; // @[:@34213.4]
  assign StickySelects_14_io_ins_0 = io_rPort_4_en_0 & _T_1671; // @[MemPrimitives.scala 125:64:@34214.4]
  assign StickySelects_14_io_ins_1 = io_rPort_6_en_0 & _T_1677; // @[MemPrimitives.scala 125:64:@34215.4]
  assign StickySelects_14_io_ins_2 = io_rPort_7_en_0 & _T_1683; // @[MemPrimitives.scala 125:64:@34216.4]
  assign StickySelects_14_io_ins_3 = io_rPort_9_en_0 & _T_1689; // @[MemPrimitives.scala 125:64:@34217.4]
  assign StickySelects_15_clock = clock; // @[:@34264.4]
  assign StickySelects_15_reset = reset; // @[:@34265.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_1713; // @[MemPrimitives.scala 125:64:@34266.4]
  assign StickySelects_15_io_ins_1 = io_rPort_1_en_0 & _T_1719; // @[MemPrimitives.scala 125:64:@34267.4]
  assign StickySelects_15_io_ins_2 = io_rPort_2_en_0 & _T_1725; // @[MemPrimitives.scala 125:64:@34268.4]
  assign StickySelects_15_io_ins_3 = io_rPort_3_en_0 & _T_1731; // @[MemPrimitives.scala 125:64:@34269.4]
  assign StickySelects_15_io_ins_4 = io_rPort_5_en_0 & _T_1737; // @[MemPrimitives.scala 125:64:@34270.4]
  assign StickySelects_15_io_ins_5 = io_rPort_8_en_0 & _T_1743; // @[MemPrimitives.scala 125:64:@34271.4]
  assign StickySelects_16_clock = clock; // @[:@34318.4]
  assign StickySelects_16_reset = reset; // @[:@34319.4]
  assign StickySelects_16_io_ins_0 = io_rPort_4_en_0 & _T_1775; // @[MemPrimitives.scala 125:64:@34320.4]
  assign StickySelects_16_io_ins_1 = io_rPort_6_en_0 & _T_1781; // @[MemPrimitives.scala 125:64:@34321.4]
  assign StickySelects_16_io_ins_2 = io_rPort_7_en_0 & _T_1787; // @[MemPrimitives.scala 125:64:@34322.4]
  assign StickySelects_16_io_ins_3 = io_rPort_9_en_0 & _T_1793; // @[MemPrimitives.scala 125:64:@34323.4]
  assign StickySelects_17_clock = clock; // @[:@34370.4]
  assign StickySelects_17_reset = reset; // @[:@34371.4]
  assign StickySelects_17_io_ins_0 = io_rPort_0_en_0 & _T_1817; // @[MemPrimitives.scala 125:64:@34372.4]
  assign StickySelects_17_io_ins_1 = io_rPort_1_en_0 & _T_1823; // @[MemPrimitives.scala 125:64:@34373.4]
  assign StickySelects_17_io_ins_2 = io_rPort_2_en_0 & _T_1829; // @[MemPrimitives.scala 125:64:@34374.4]
  assign StickySelects_17_io_ins_3 = io_rPort_3_en_0 & _T_1835; // @[MemPrimitives.scala 125:64:@34375.4]
  assign StickySelects_17_io_ins_4 = io_rPort_5_en_0 & _T_1841; // @[MemPrimitives.scala 125:64:@34376.4]
  assign StickySelects_17_io_ins_5 = io_rPort_8_en_0 & _T_1847; // @[MemPrimitives.scala 125:64:@34377.4]
  assign StickySelects_18_clock = clock; // @[:@34424.4]
  assign StickySelects_18_reset = reset; // @[:@34425.4]
  assign StickySelects_18_io_ins_0 = io_rPort_4_en_0 & _T_1879; // @[MemPrimitives.scala 125:64:@34426.4]
  assign StickySelects_18_io_ins_1 = io_rPort_6_en_0 & _T_1885; // @[MemPrimitives.scala 125:64:@34427.4]
  assign StickySelects_18_io_ins_2 = io_rPort_7_en_0 & _T_1891; // @[MemPrimitives.scala 125:64:@34428.4]
  assign StickySelects_18_io_ins_3 = io_rPort_9_en_0 & _T_1897; // @[MemPrimitives.scala 125:64:@34429.4]
  assign StickySelects_19_clock = clock; // @[:@34476.4]
  assign StickySelects_19_reset = reset; // @[:@34477.4]
  assign StickySelects_19_io_ins_0 = io_rPort_0_en_0 & _T_1921; // @[MemPrimitives.scala 125:64:@34478.4]
  assign StickySelects_19_io_ins_1 = io_rPort_1_en_0 & _T_1927; // @[MemPrimitives.scala 125:64:@34479.4]
  assign StickySelects_19_io_ins_2 = io_rPort_2_en_0 & _T_1933; // @[MemPrimitives.scala 125:64:@34480.4]
  assign StickySelects_19_io_ins_3 = io_rPort_3_en_0 & _T_1939; // @[MemPrimitives.scala 125:64:@34481.4]
  assign StickySelects_19_io_ins_4 = io_rPort_5_en_0 & _T_1945; // @[MemPrimitives.scala 125:64:@34482.4]
  assign StickySelects_19_io_ins_5 = io_rPort_8_en_0 & _T_1951; // @[MemPrimitives.scala 125:64:@34483.4]
  assign StickySelects_20_clock = clock; // @[:@34530.4]
  assign StickySelects_20_reset = reset; // @[:@34531.4]
  assign StickySelects_20_io_ins_0 = io_rPort_4_en_0 & _T_1983; // @[MemPrimitives.scala 125:64:@34532.4]
  assign StickySelects_20_io_ins_1 = io_rPort_6_en_0 & _T_1989; // @[MemPrimitives.scala 125:64:@34533.4]
  assign StickySelects_20_io_ins_2 = io_rPort_7_en_0 & _T_1995; // @[MemPrimitives.scala 125:64:@34534.4]
  assign StickySelects_20_io_ins_3 = io_rPort_9_en_0 & _T_2001; // @[MemPrimitives.scala 125:64:@34535.4]
  assign StickySelects_21_clock = clock; // @[:@34582.4]
  assign StickySelects_21_reset = reset; // @[:@34583.4]
  assign StickySelects_21_io_ins_0 = io_rPort_0_en_0 & _T_2025; // @[MemPrimitives.scala 125:64:@34584.4]
  assign StickySelects_21_io_ins_1 = io_rPort_1_en_0 & _T_2031; // @[MemPrimitives.scala 125:64:@34585.4]
  assign StickySelects_21_io_ins_2 = io_rPort_2_en_0 & _T_2037; // @[MemPrimitives.scala 125:64:@34586.4]
  assign StickySelects_21_io_ins_3 = io_rPort_3_en_0 & _T_2043; // @[MemPrimitives.scala 125:64:@34587.4]
  assign StickySelects_21_io_ins_4 = io_rPort_5_en_0 & _T_2049; // @[MemPrimitives.scala 125:64:@34588.4]
  assign StickySelects_21_io_ins_5 = io_rPort_8_en_0 & _T_2055; // @[MemPrimitives.scala 125:64:@34589.4]
  assign StickySelects_22_clock = clock; // @[:@34636.4]
  assign StickySelects_22_reset = reset; // @[:@34637.4]
  assign StickySelects_22_io_ins_0 = io_rPort_4_en_0 & _T_2087; // @[MemPrimitives.scala 125:64:@34638.4]
  assign StickySelects_22_io_ins_1 = io_rPort_6_en_0 & _T_2093; // @[MemPrimitives.scala 125:64:@34639.4]
  assign StickySelects_22_io_ins_2 = io_rPort_7_en_0 & _T_2099; // @[MemPrimitives.scala 125:64:@34640.4]
  assign StickySelects_22_io_ins_3 = io_rPort_9_en_0 & _T_2105; // @[MemPrimitives.scala 125:64:@34641.4]
  assign StickySelects_23_clock = clock; // @[:@34688.4]
  assign StickySelects_23_reset = reset; // @[:@34689.4]
  assign StickySelects_23_io_ins_0 = io_rPort_0_en_0 & _T_2129; // @[MemPrimitives.scala 125:64:@34690.4]
  assign StickySelects_23_io_ins_1 = io_rPort_1_en_0 & _T_2135; // @[MemPrimitives.scala 125:64:@34691.4]
  assign StickySelects_23_io_ins_2 = io_rPort_2_en_0 & _T_2141; // @[MemPrimitives.scala 125:64:@34692.4]
  assign StickySelects_23_io_ins_3 = io_rPort_3_en_0 & _T_2147; // @[MemPrimitives.scala 125:64:@34693.4]
  assign StickySelects_23_io_ins_4 = io_rPort_5_en_0 & _T_2153; // @[MemPrimitives.scala 125:64:@34694.4]
  assign StickySelects_23_io_ins_5 = io_rPort_8_en_0 & _T_2159; // @[MemPrimitives.scala 125:64:@34695.4]
  assign RetimeWrapper_clock = clock; // @[:@34763.4]
  assign RetimeWrapper_reset = reset; // @[:@34764.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34766.4]
  assign RetimeWrapper_io_in = _T_985 & io_rPort_0_en_0; // @[package.scala 94:16:@34765.4]
  assign RetimeWrapper_1_clock = clock; // @[:@34771.4]
  assign RetimeWrapper_1_reset = reset; // @[:@34772.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34774.4]
  assign RetimeWrapper_1_io_in = _T_1089 & io_rPort_0_en_0; // @[package.scala 94:16:@34773.4]
  assign RetimeWrapper_2_clock = clock; // @[:@34779.4]
  assign RetimeWrapper_2_reset = reset; // @[:@34780.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34782.4]
  assign RetimeWrapper_2_io_in = _T_1193 & io_rPort_0_en_0; // @[package.scala 94:16:@34781.4]
  assign RetimeWrapper_3_clock = clock; // @[:@34787.4]
  assign RetimeWrapper_3_reset = reset; // @[:@34788.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34790.4]
  assign RetimeWrapper_3_io_in = _T_1297 & io_rPort_0_en_0; // @[package.scala 94:16:@34789.4]
  assign RetimeWrapper_4_clock = clock; // @[:@34795.4]
  assign RetimeWrapper_4_reset = reset; // @[:@34796.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34798.4]
  assign RetimeWrapper_4_io_in = _T_1401 & io_rPort_0_en_0; // @[package.scala 94:16:@34797.4]
  assign RetimeWrapper_5_clock = clock; // @[:@34803.4]
  assign RetimeWrapper_5_reset = reset; // @[:@34804.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34806.4]
  assign RetimeWrapper_5_io_in = _T_1505 & io_rPort_0_en_0; // @[package.scala 94:16:@34805.4]
  assign RetimeWrapper_6_clock = clock; // @[:@34811.4]
  assign RetimeWrapper_6_reset = reset; // @[:@34812.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34814.4]
  assign RetimeWrapper_6_io_in = _T_1609 & io_rPort_0_en_0; // @[package.scala 94:16:@34813.4]
  assign RetimeWrapper_7_clock = clock; // @[:@34819.4]
  assign RetimeWrapper_7_reset = reset; // @[:@34820.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34822.4]
  assign RetimeWrapper_7_io_in = _T_1713 & io_rPort_0_en_0; // @[package.scala 94:16:@34821.4]
  assign RetimeWrapper_8_clock = clock; // @[:@34827.4]
  assign RetimeWrapper_8_reset = reset; // @[:@34828.4]
  assign RetimeWrapper_8_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34830.4]
  assign RetimeWrapper_8_io_in = _T_1817 & io_rPort_0_en_0; // @[package.scala 94:16:@34829.4]
  assign RetimeWrapper_9_clock = clock; // @[:@34835.4]
  assign RetimeWrapper_9_reset = reset; // @[:@34836.4]
  assign RetimeWrapper_9_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34838.4]
  assign RetimeWrapper_9_io_in = _T_1921 & io_rPort_0_en_0; // @[package.scala 94:16:@34837.4]
  assign RetimeWrapper_10_clock = clock; // @[:@34843.4]
  assign RetimeWrapper_10_reset = reset; // @[:@34844.4]
  assign RetimeWrapper_10_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34846.4]
  assign RetimeWrapper_10_io_in = _T_2025 & io_rPort_0_en_0; // @[package.scala 94:16:@34845.4]
  assign RetimeWrapper_11_clock = clock; // @[:@34851.4]
  assign RetimeWrapper_11_reset = reset; // @[:@34852.4]
  assign RetimeWrapper_11_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@34854.4]
  assign RetimeWrapper_11_io_in = _T_2129 & io_rPort_0_en_0; // @[package.scala 94:16:@34853.4]
  assign RetimeWrapper_12_clock = clock; // @[:@34907.4]
  assign RetimeWrapper_12_reset = reset; // @[:@34908.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34910.4]
  assign RetimeWrapper_12_io_in = _T_991 & io_rPort_1_en_0; // @[package.scala 94:16:@34909.4]
  assign RetimeWrapper_13_clock = clock; // @[:@34915.4]
  assign RetimeWrapper_13_reset = reset; // @[:@34916.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34918.4]
  assign RetimeWrapper_13_io_in = _T_1095 & io_rPort_1_en_0; // @[package.scala 94:16:@34917.4]
  assign RetimeWrapper_14_clock = clock; // @[:@34923.4]
  assign RetimeWrapper_14_reset = reset; // @[:@34924.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34926.4]
  assign RetimeWrapper_14_io_in = _T_1199 & io_rPort_1_en_0; // @[package.scala 94:16:@34925.4]
  assign RetimeWrapper_15_clock = clock; // @[:@34931.4]
  assign RetimeWrapper_15_reset = reset; // @[:@34932.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34934.4]
  assign RetimeWrapper_15_io_in = _T_1303 & io_rPort_1_en_0; // @[package.scala 94:16:@34933.4]
  assign RetimeWrapper_16_clock = clock; // @[:@34939.4]
  assign RetimeWrapper_16_reset = reset; // @[:@34940.4]
  assign RetimeWrapper_16_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34942.4]
  assign RetimeWrapper_16_io_in = _T_1407 & io_rPort_1_en_0; // @[package.scala 94:16:@34941.4]
  assign RetimeWrapper_17_clock = clock; // @[:@34947.4]
  assign RetimeWrapper_17_reset = reset; // @[:@34948.4]
  assign RetimeWrapper_17_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34950.4]
  assign RetimeWrapper_17_io_in = _T_1511 & io_rPort_1_en_0; // @[package.scala 94:16:@34949.4]
  assign RetimeWrapper_18_clock = clock; // @[:@34955.4]
  assign RetimeWrapper_18_reset = reset; // @[:@34956.4]
  assign RetimeWrapper_18_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34958.4]
  assign RetimeWrapper_18_io_in = _T_1615 & io_rPort_1_en_0; // @[package.scala 94:16:@34957.4]
  assign RetimeWrapper_19_clock = clock; // @[:@34963.4]
  assign RetimeWrapper_19_reset = reset; // @[:@34964.4]
  assign RetimeWrapper_19_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34966.4]
  assign RetimeWrapper_19_io_in = _T_1719 & io_rPort_1_en_0; // @[package.scala 94:16:@34965.4]
  assign RetimeWrapper_20_clock = clock; // @[:@34971.4]
  assign RetimeWrapper_20_reset = reset; // @[:@34972.4]
  assign RetimeWrapper_20_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34974.4]
  assign RetimeWrapper_20_io_in = _T_1823 & io_rPort_1_en_0; // @[package.scala 94:16:@34973.4]
  assign RetimeWrapper_21_clock = clock; // @[:@34979.4]
  assign RetimeWrapper_21_reset = reset; // @[:@34980.4]
  assign RetimeWrapper_21_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34982.4]
  assign RetimeWrapper_21_io_in = _T_1927 & io_rPort_1_en_0; // @[package.scala 94:16:@34981.4]
  assign RetimeWrapper_22_clock = clock; // @[:@34987.4]
  assign RetimeWrapper_22_reset = reset; // @[:@34988.4]
  assign RetimeWrapper_22_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34990.4]
  assign RetimeWrapper_22_io_in = _T_2031 & io_rPort_1_en_0; // @[package.scala 94:16:@34989.4]
  assign RetimeWrapper_23_clock = clock; // @[:@34995.4]
  assign RetimeWrapper_23_reset = reset; // @[:@34996.4]
  assign RetimeWrapper_23_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@34998.4]
  assign RetimeWrapper_23_io_in = _T_2135 & io_rPort_1_en_0; // @[package.scala 94:16:@34997.4]
  assign RetimeWrapper_24_clock = clock; // @[:@35051.4]
  assign RetimeWrapper_24_reset = reset; // @[:@35052.4]
  assign RetimeWrapper_24_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35054.4]
  assign RetimeWrapper_24_io_in = _T_997 & io_rPort_2_en_0; // @[package.scala 94:16:@35053.4]
  assign RetimeWrapper_25_clock = clock; // @[:@35059.4]
  assign RetimeWrapper_25_reset = reset; // @[:@35060.4]
  assign RetimeWrapper_25_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35062.4]
  assign RetimeWrapper_25_io_in = _T_1101 & io_rPort_2_en_0; // @[package.scala 94:16:@35061.4]
  assign RetimeWrapper_26_clock = clock; // @[:@35067.4]
  assign RetimeWrapper_26_reset = reset; // @[:@35068.4]
  assign RetimeWrapper_26_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35070.4]
  assign RetimeWrapper_26_io_in = _T_1205 & io_rPort_2_en_0; // @[package.scala 94:16:@35069.4]
  assign RetimeWrapper_27_clock = clock; // @[:@35075.4]
  assign RetimeWrapper_27_reset = reset; // @[:@35076.4]
  assign RetimeWrapper_27_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35078.4]
  assign RetimeWrapper_27_io_in = _T_1309 & io_rPort_2_en_0; // @[package.scala 94:16:@35077.4]
  assign RetimeWrapper_28_clock = clock; // @[:@35083.4]
  assign RetimeWrapper_28_reset = reset; // @[:@35084.4]
  assign RetimeWrapper_28_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35086.4]
  assign RetimeWrapper_28_io_in = _T_1413 & io_rPort_2_en_0; // @[package.scala 94:16:@35085.4]
  assign RetimeWrapper_29_clock = clock; // @[:@35091.4]
  assign RetimeWrapper_29_reset = reset; // @[:@35092.4]
  assign RetimeWrapper_29_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35094.4]
  assign RetimeWrapper_29_io_in = _T_1517 & io_rPort_2_en_0; // @[package.scala 94:16:@35093.4]
  assign RetimeWrapper_30_clock = clock; // @[:@35099.4]
  assign RetimeWrapper_30_reset = reset; // @[:@35100.4]
  assign RetimeWrapper_30_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35102.4]
  assign RetimeWrapper_30_io_in = _T_1621 & io_rPort_2_en_0; // @[package.scala 94:16:@35101.4]
  assign RetimeWrapper_31_clock = clock; // @[:@35107.4]
  assign RetimeWrapper_31_reset = reset; // @[:@35108.4]
  assign RetimeWrapper_31_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35110.4]
  assign RetimeWrapper_31_io_in = _T_1725 & io_rPort_2_en_0; // @[package.scala 94:16:@35109.4]
  assign RetimeWrapper_32_clock = clock; // @[:@35115.4]
  assign RetimeWrapper_32_reset = reset; // @[:@35116.4]
  assign RetimeWrapper_32_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35118.4]
  assign RetimeWrapper_32_io_in = _T_1829 & io_rPort_2_en_0; // @[package.scala 94:16:@35117.4]
  assign RetimeWrapper_33_clock = clock; // @[:@35123.4]
  assign RetimeWrapper_33_reset = reset; // @[:@35124.4]
  assign RetimeWrapper_33_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35126.4]
  assign RetimeWrapper_33_io_in = _T_1933 & io_rPort_2_en_0; // @[package.scala 94:16:@35125.4]
  assign RetimeWrapper_34_clock = clock; // @[:@35131.4]
  assign RetimeWrapper_34_reset = reset; // @[:@35132.4]
  assign RetimeWrapper_34_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35134.4]
  assign RetimeWrapper_34_io_in = _T_2037 & io_rPort_2_en_0; // @[package.scala 94:16:@35133.4]
  assign RetimeWrapper_35_clock = clock; // @[:@35139.4]
  assign RetimeWrapper_35_reset = reset; // @[:@35140.4]
  assign RetimeWrapper_35_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@35142.4]
  assign RetimeWrapper_35_io_in = _T_2141 & io_rPort_2_en_0; // @[package.scala 94:16:@35141.4]
  assign RetimeWrapper_36_clock = clock; // @[:@35195.4]
  assign RetimeWrapper_36_reset = reset; // @[:@35196.4]
  assign RetimeWrapper_36_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35198.4]
  assign RetimeWrapper_36_io_in = _T_1003 & io_rPort_3_en_0; // @[package.scala 94:16:@35197.4]
  assign RetimeWrapper_37_clock = clock; // @[:@35203.4]
  assign RetimeWrapper_37_reset = reset; // @[:@35204.4]
  assign RetimeWrapper_37_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35206.4]
  assign RetimeWrapper_37_io_in = _T_1107 & io_rPort_3_en_0; // @[package.scala 94:16:@35205.4]
  assign RetimeWrapper_38_clock = clock; // @[:@35211.4]
  assign RetimeWrapper_38_reset = reset; // @[:@35212.4]
  assign RetimeWrapper_38_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35214.4]
  assign RetimeWrapper_38_io_in = _T_1211 & io_rPort_3_en_0; // @[package.scala 94:16:@35213.4]
  assign RetimeWrapper_39_clock = clock; // @[:@35219.4]
  assign RetimeWrapper_39_reset = reset; // @[:@35220.4]
  assign RetimeWrapper_39_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35222.4]
  assign RetimeWrapper_39_io_in = _T_1315 & io_rPort_3_en_0; // @[package.scala 94:16:@35221.4]
  assign RetimeWrapper_40_clock = clock; // @[:@35227.4]
  assign RetimeWrapper_40_reset = reset; // @[:@35228.4]
  assign RetimeWrapper_40_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35230.4]
  assign RetimeWrapper_40_io_in = _T_1419 & io_rPort_3_en_0; // @[package.scala 94:16:@35229.4]
  assign RetimeWrapper_41_clock = clock; // @[:@35235.4]
  assign RetimeWrapper_41_reset = reset; // @[:@35236.4]
  assign RetimeWrapper_41_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35238.4]
  assign RetimeWrapper_41_io_in = _T_1523 & io_rPort_3_en_0; // @[package.scala 94:16:@35237.4]
  assign RetimeWrapper_42_clock = clock; // @[:@35243.4]
  assign RetimeWrapper_42_reset = reset; // @[:@35244.4]
  assign RetimeWrapper_42_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35246.4]
  assign RetimeWrapper_42_io_in = _T_1627 & io_rPort_3_en_0; // @[package.scala 94:16:@35245.4]
  assign RetimeWrapper_43_clock = clock; // @[:@35251.4]
  assign RetimeWrapper_43_reset = reset; // @[:@35252.4]
  assign RetimeWrapper_43_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35254.4]
  assign RetimeWrapper_43_io_in = _T_1731 & io_rPort_3_en_0; // @[package.scala 94:16:@35253.4]
  assign RetimeWrapper_44_clock = clock; // @[:@35259.4]
  assign RetimeWrapper_44_reset = reset; // @[:@35260.4]
  assign RetimeWrapper_44_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35262.4]
  assign RetimeWrapper_44_io_in = _T_1835 & io_rPort_3_en_0; // @[package.scala 94:16:@35261.4]
  assign RetimeWrapper_45_clock = clock; // @[:@35267.4]
  assign RetimeWrapper_45_reset = reset; // @[:@35268.4]
  assign RetimeWrapper_45_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35270.4]
  assign RetimeWrapper_45_io_in = _T_1939 & io_rPort_3_en_0; // @[package.scala 94:16:@35269.4]
  assign RetimeWrapper_46_clock = clock; // @[:@35275.4]
  assign RetimeWrapper_46_reset = reset; // @[:@35276.4]
  assign RetimeWrapper_46_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35278.4]
  assign RetimeWrapper_46_io_in = _T_2043 & io_rPort_3_en_0; // @[package.scala 94:16:@35277.4]
  assign RetimeWrapper_47_clock = clock; // @[:@35283.4]
  assign RetimeWrapper_47_reset = reset; // @[:@35284.4]
  assign RetimeWrapper_47_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@35286.4]
  assign RetimeWrapper_47_io_in = _T_2147 & io_rPort_3_en_0; // @[package.scala 94:16:@35285.4]
  assign RetimeWrapper_48_clock = clock; // @[:@35339.4]
  assign RetimeWrapper_48_reset = reset; // @[:@35340.4]
  assign RetimeWrapper_48_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35342.4]
  assign RetimeWrapper_48_io_in = _T_943 & io_rPort_4_en_0; // @[package.scala 94:16:@35341.4]
  assign RetimeWrapper_49_clock = clock; // @[:@35347.4]
  assign RetimeWrapper_49_reset = reset; // @[:@35348.4]
  assign RetimeWrapper_49_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35350.4]
  assign RetimeWrapper_49_io_in = _T_1047 & io_rPort_4_en_0; // @[package.scala 94:16:@35349.4]
  assign RetimeWrapper_50_clock = clock; // @[:@35355.4]
  assign RetimeWrapper_50_reset = reset; // @[:@35356.4]
  assign RetimeWrapper_50_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35358.4]
  assign RetimeWrapper_50_io_in = _T_1151 & io_rPort_4_en_0; // @[package.scala 94:16:@35357.4]
  assign RetimeWrapper_51_clock = clock; // @[:@35363.4]
  assign RetimeWrapper_51_reset = reset; // @[:@35364.4]
  assign RetimeWrapper_51_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35366.4]
  assign RetimeWrapper_51_io_in = _T_1255 & io_rPort_4_en_0; // @[package.scala 94:16:@35365.4]
  assign RetimeWrapper_52_clock = clock; // @[:@35371.4]
  assign RetimeWrapper_52_reset = reset; // @[:@35372.4]
  assign RetimeWrapper_52_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35374.4]
  assign RetimeWrapper_52_io_in = _T_1359 & io_rPort_4_en_0; // @[package.scala 94:16:@35373.4]
  assign RetimeWrapper_53_clock = clock; // @[:@35379.4]
  assign RetimeWrapper_53_reset = reset; // @[:@35380.4]
  assign RetimeWrapper_53_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35382.4]
  assign RetimeWrapper_53_io_in = _T_1463 & io_rPort_4_en_0; // @[package.scala 94:16:@35381.4]
  assign RetimeWrapper_54_clock = clock; // @[:@35387.4]
  assign RetimeWrapper_54_reset = reset; // @[:@35388.4]
  assign RetimeWrapper_54_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35390.4]
  assign RetimeWrapper_54_io_in = _T_1567 & io_rPort_4_en_0; // @[package.scala 94:16:@35389.4]
  assign RetimeWrapper_55_clock = clock; // @[:@35395.4]
  assign RetimeWrapper_55_reset = reset; // @[:@35396.4]
  assign RetimeWrapper_55_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35398.4]
  assign RetimeWrapper_55_io_in = _T_1671 & io_rPort_4_en_0; // @[package.scala 94:16:@35397.4]
  assign RetimeWrapper_56_clock = clock; // @[:@35403.4]
  assign RetimeWrapper_56_reset = reset; // @[:@35404.4]
  assign RetimeWrapper_56_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35406.4]
  assign RetimeWrapper_56_io_in = _T_1775 & io_rPort_4_en_0; // @[package.scala 94:16:@35405.4]
  assign RetimeWrapper_57_clock = clock; // @[:@35411.4]
  assign RetimeWrapper_57_reset = reset; // @[:@35412.4]
  assign RetimeWrapper_57_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35414.4]
  assign RetimeWrapper_57_io_in = _T_1879 & io_rPort_4_en_0; // @[package.scala 94:16:@35413.4]
  assign RetimeWrapper_58_clock = clock; // @[:@35419.4]
  assign RetimeWrapper_58_reset = reset; // @[:@35420.4]
  assign RetimeWrapper_58_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35422.4]
  assign RetimeWrapper_58_io_in = _T_1983 & io_rPort_4_en_0; // @[package.scala 94:16:@35421.4]
  assign RetimeWrapper_59_clock = clock; // @[:@35427.4]
  assign RetimeWrapper_59_reset = reset; // @[:@35428.4]
  assign RetimeWrapper_59_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@35430.4]
  assign RetimeWrapper_59_io_in = _T_2087 & io_rPort_4_en_0; // @[package.scala 94:16:@35429.4]
  assign RetimeWrapper_60_clock = clock; // @[:@35483.4]
  assign RetimeWrapper_60_reset = reset; // @[:@35484.4]
  assign RetimeWrapper_60_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35486.4]
  assign RetimeWrapper_60_io_in = _T_1009 & io_rPort_5_en_0; // @[package.scala 94:16:@35485.4]
  assign RetimeWrapper_61_clock = clock; // @[:@35491.4]
  assign RetimeWrapper_61_reset = reset; // @[:@35492.4]
  assign RetimeWrapper_61_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35494.4]
  assign RetimeWrapper_61_io_in = _T_1113 & io_rPort_5_en_0; // @[package.scala 94:16:@35493.4]
  assign RetimeWrapper_62_clock = clock; // @[:@35499.4]
  assign RetimeWrapper_62_reset = reset; // @[:@35500.4]
  assign RetimeWrapper_62_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35502.4]
  assign RetimeWrapper_62_io_in = _T_1217 & io_rPort_5_en_0; // @[package.scala 94:16:@35501.4]
  assign RetimeWrapper_63_clock = clock; // @[:@35507.4]
  assign RetimeWrapper_63_reset = reset; // @[:@35508.4]
  assign RetimeWrapper_63_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35510.4]
  assign RetimeWrapper_63_io_in = _T_1321 & io_rPort_5_en_0; // @[package.scala 94:16:@35509.4]
  assign RetimeWrapper_64_clock = clock; // @[:@35515.4]
  assign RetimeWrapper_64_reset = reset; // @[:@35516.4]
  assign RetimeWrapper_64_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35518.4]
  assign RetimeWrapper_64_io_in = _T_1425 & io_rPort_5_en_0; // @[package.scala 94:16:@35517.4]
  assign RetimeWrapper_65_clock = clock; // @[:@35523.4]
  assign RetimeWrapper_65_reset = reset; // @[:@35524.4]
  assign RetimeWrapper_65_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35526.4]
  assign RetimeWrapper_65_io_in = _T_1529 & io_rPort_5_en_0; // @[package.scala 94:16:@35525.4]
  assign RetimeWrapper_66_clock = clock; // @[:@35531.4]
  assign RetimeWrapper_66_reset = reset; // @[:@35532.4]
  assign RetimeWrapper_66_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35534.4]
  assign RetimeWrapper_66_io_in = _T_1633 & io_rPort_5_en_0; // @[package.scala 94:16:@35533.4]
  assign RetimeWrapper_67_clock = clock; // @[:@35539.4]
  assign RetimeWrapper_67_reset = reset; // @[:@35540.4]
  assign RetimeWrapper_67_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35542.4]
  assign RetimeWrapper_67_io_in = _T_1737 & io_rPort_5_en_0; // @[package.scala 94:16:@35541.4]
  assign RetimeWrapper_68_clock = clock; // @[:@35547.4]
  assign RetimeWrapper_68_reset = reset; // @[:@35548.4]
  assign RetimeWrapper_68_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35550.4]
  assign RetimeWrapper_68_io_in = _T_1841 & io_rPort_5_en_0; // @[package.scala 94:16:@35549.4]
  assign RetimeWrapper_69_clock = clock; // @[:@35555.4]
  assign RetimeWrapper_69_reset = reset; // @[:@35556.4]
  assign RetimeWrapper_69_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35558.4]
  assign RetimeWrapper_69_io_in = _T_1945 & io_rPort_5_en_0; // @[package.scala 94:16:@35557.4]
  assign RetimeWrapper_70_clock = clock; // @[:@35563.4]
  assign RetimeWrapper_70_reset = reset; // @[:@35564.4]
  assign RetimeWrapper_70_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35566.4]
  assign RetimeWrapper_70_io_in = _T_2049 & io_rPort_5_en_0; // @[package.scala 94:16:@35565.4]
  assign RetimeWrapper_71_clock = clock; // @[:@35571.4]
  assign RetimeWrapper_71_reset = reset; // @[:@35572.4]
  assign RetimeWrapper_71_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@35574.4]
  assign RetimeWrapper_71_io_in = _T_2153 & io_rPort_5_en_0; // @[package.scala 94:16:@35573.4]
  assign RetimeWrapper_72_clock = clock; // @[:@35627.4]
  assign RetimeWrapper_72_reset = reset; // @[:@35628.4]
  assign RetimeWrapper_72_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35630.4]
  assign RetimeWrapper_72_io_in = _T_949 & io_rPort_6_en_0; // @[package.scala 94:16:@35629.4]
  assign RetimeWrapper_73_clock = clock; // @[:@35635.4]
  assign RetimeWrapper_73_reset = reset; // @[:@35636.4]
  assign RetimeWrapper_73_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35638.4]
  assign RetimeWrapper_73_io_in = _T_1053 & io_rPort_6_en_0; // @[package.scala 94:16:@35637.4]
  assign RetimeWrapper_74_clock = clock; // @[:@35643.4]
  assign RetimeWrapper_74_reset = reset; // @[:@35644.4]
  assign RetimeWrapper_74_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35646.4]
  assign RetimeWrapper_74_io_in = _T_1157 & io_rPort_6_en_0; // @[package.scala 94:16:@35645.4]
  assign RetimeWrapper_75_clock = clock; // @[:@35651.4]
  assign RetimeWrapper_75_reset = reset; // @[:@35652.4]
  assign RetimeWrapper_75_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35654.4]
  assign RetimeWrapper_75_io_in = _T_1261 & io_rPort_6_en_0; // @[package.scala 94:16:@35653.4]
  assign RetimeWrapper_76_clock = clock; // @[:@35659.4]
  assign RetimeWrapper_76_reset = reset; // @[:@35660.4]
  assign RetimeWrapper_76_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35662.4]
  assign RetimeWrapper_76_io_in = _T_1365 & io_rPort_6_en_0; // @[package.scala 94:16:@35661.4]
  assign RetimeWrapper_77_clock = clock; // @[:@35667.4]
  assign RetimeWrapper_77_reset = reset; // @[:@35668.4]
  assign RetimeWrapper_77_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35670.4]
  assign RetimeWrapper_77_io_in = _T_1469 & io_rPort_6_en_0; // @[package.scala 94:16:@35669.4]
  assign RetimeWrapper_78_clock = clock; // @[:@35675.4]
  assign RetimeWrapper_78_reset = reset; // @[:@35676.4]
  assign RetimeWrapper_78_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35678.4]
  assign RetimeWrapper_78_io_in = _T_1573 & io_rPort_6_en_0; // @[package.scala 94:16:@35677.4]
  assign RetimeWrapper_79_clock = clock; // @[:@35683.4]
  assign RetimeWrapper_79_reset = reset; // @[:@35684.4]
  assign RetimeWrapper_79_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35686.4]
  assign RetimeWrapper_79_io_in = _T_1677 & io_rPort_6_en_0; // @[package.scala 94:16:@35685.4]
  assign RetimeWrapper_80_clock = clock; // @[:@35691.4]
  assign RetimeWrapper_80_reset = reset; // @[:@35692.4]
  assign RetimeWrapper_80_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35694.4]
  assign RetimeWrapper_80_io_in = _T_1781 & io_rPort_6_en_0; // @[package.scala 94:16:@35693.4]
  assign RetimeWrapper_81_clock = clock; // @[:@35699.4]
  assign RetimeWrapper_81_reset = reset; // @[:@35700.4]
  assign RetimeWrapper_81_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35702.4]
  assign RetimeWrapper_81_io_in = _T_1885 & io_rPort_6_en_0; // @[package.scala 94:16:@35701.4]
  assign RetimeWrapper_82_clock = clock; // @[:@35707.4]
  assign RetimeWrapper_82_reset = reset; // @[:@35708.4]
  assign RetimeWrapper_82_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35710.4]
  assign RetimeWrapper_82_io_in = _T_1989 & io_rPort_6_en_0; // @[package.scala 94:16:@35709.4]
  assign RetimeWrapper_83_clock = clock; // @[:@35715.4]
  assign RetimeWrapper_83_reset = reset; // @[:@35716.4]
  assign RetimeWrapper_83_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@35718.4]
  assign RetimeWrapper_83_io_in = _T_2093 & io_rPort_6_en_0; // @[package.scala 94:16:@35717.4]
  assign RetimeWrapper_84_clock = clock; // @[:@35771.4]
  assign RetimeWrapper_84_reset = reset; // @[:@35772.4]
  assign RetimeWrapper_84_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35774.4]
  assign RetimeWrapper_84_io_in = _T_955 & io_rPort_7_en_0; // @[package.scala 94:16:@35773.4]
  assign RetimeWrapper_85_clock = clock; // @[:@35779.4]
  assign RetimeWrapper_85_reset = reset; // @[:@35780.4]
  assign RetimeWrapper_85_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35782.4]
  assign RetimeWrapper_85_io_in = _T_1059 & io_rPort_7_en_0; // @[package.scala 94:16:@35781.4]
  assign RetimeWrapper_86_clock = clock; // @[:@35787.4]
  assign RetimeWrapper_86_reset = reset; // @[:@35788.4]
  assign RetimeWrapper_86_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35790.4]
  assign RetimeWrapper_86_io_in = _T_1163 & io_rPort_7_en_0; // @[package.scala 94:16:@35789.4]
  assign RetimeWrapper_87_clock = clock; // @[:@35795.4]
  assign RetimeWrapper_87_reset = reset; // @[:@35796.4]
  assign RetimeWrapper_87_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35798.4]
  assign RetimeWrapper_87_io_in = _T_1267 & io_rPort_7_en_0; // @[package.scala 94:16:@35797.4]
  assign RetimeWrapper_88_clock = clock; // @[:@35803.4]
  assign RetimeWrapper_88_reset = reset; // @[:@35804.4]
  assign RetimeWrapper_88_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35806.4]
  assign RetimeWrapper_88_io_in = _T_1371 & io_rPort_7_en_0; // @[package.scala 94:16:@35805.4]
  assign RetimeWrapper_89_clock = clock; // @[:@35811.4]
  assign RetimeWrapper_89_reset = reset; // @[:@35812.4]
  assign RetimeWrapper_89_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35814.4]
  assign RetimeWrapper_89_io_in = _T_1475 & io_rPort_7_en_0; // @[package.scala 94:16:@35813.4]
  assign RetimeWrapper_90_clock = clock; // @[:@35819.4]
  assign RetimeWrapper_90_reset = reset; // @[:@35820.4]
  assign RetimeWrapper_90_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35822.4]
  assign RetimeWrapper_90_io_in = _T_1579 & io_rPort_7_en_0; // @[package.scala 94:16:@35821.4]
  assign RetimeWrapper_91_clock = clock; // @[:@35827.4]
  assign RetimeWrapper_91_reset = reset; // @[:@35828.4]
  assign RetimeWrapper_91_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35830.4]
  assign RetimeWrapper_91_io_in = _T_1683 & io_rPort_7_en_0; // @[package.scala 94:16:@35829.4]
  assign RetimeWrapper_92_clock = clock; // @[:@35835.4]
  assign RetimeWrapper_92_reset = reset; // @[:@35836.4]
  assign RetimeWrapper_92_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35838.4]
  assign RetimeWrapper_92_io_in = _T_1787 & io_rPort_7_en_0; // @[package.scala 94:16:@35837.4]
  assign RetimeWrapper_93_clock = clock; // @[:@35843.4]
  assign RetimeWrapper_93_reset = reset; // @[:@35844.4]
  assign RetimeWrapper_93_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35846.4]
  assign RetimeWrapper_93_io_in = _T_1891 & io_rPort_7_en_0; // @[package.scala 94:16:@35845.4]
  assign RetimeWrapper_94_clock = clock; // @[:@35851.4]
  assign RetimeWrapper_94_reset = reset; // @[:@35852.4]
  assign RetimeWrapper_94_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35854.4]
  assign RetimeWrapper_94_io_in = _T_1995 & io_rPort_7_en_0; // @[package.scala 94:16:@35853.4]
  assign RetimeWrapper_95_clock = clock; // @[:@35859.4]
  assign RetimeWrapper_95_reset = reset; // @[:@35860.4]
  assign RetimeWrapper_95_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@35862.4]
  assign RetimeWrapper_95_io_in = _T_2099 & io_rPort_7_en_0; // @[package.scala 94:16:@35861.4]
  assign RetimeWrapper_96_clock = clock; // @[:@35915.4]
  assign RetimeWrapper_96_reset = reset; // @[:@35916.4]
  assign RetimeWrapper_96_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35918.4]
  assign RetimeWrapper_96_io_in = _T_1015 & io_rPort_8_en_0; // @[package.scala 94:16:@35917.4]
  assign RetimeWrapper_97_clock = clock; // @[:@35923.4]
  assign RetimeWrapper_97_reset = reset; // @[:@35924.4]
  assign RetimeWrapper_97_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35926.4]
  assign RetimeWrapper_97_io_in = _T_1119 & io_rPort_8_en_0; // @[package.scala 94:16:@35925.4]
  assign RetimeWrapper_98_clock = clock; // @[:@35931.4]
  assign RetimeWrapper_98_reset = reset; // @[:@35932.4]
  assign RetimeWrapper_98_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35934.4]
  assign RetimeWrapper_98_io_in = _T_1223 & io_rPort_8_en_0; // @[package.scala 94:16:@35933.4]
  assign RetimeWrapper_99_clock = clock; // @[:@35939.4]
  assign RetimeWrapper_99_reset = reset; // @[:@35940.4]
  assign RetimeWrapper_99_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35942.4]
  assign RetimeWrapper_99_io_in = _T_1327 & io_rPort_8_en_0; // @[package.scala 94:16:@35941.4]
  assign RetimeWrapper_100_clock = clock; // @[:@35947.4]
  assign RetimeWrapper_100_reset = reset; // @[:@35948.4]
  assign RetimeWrapper_100_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35950.4]
  assign RetimeWrapper_100_io_in = _T_1431 & io_rPort_8_en_0; // @[package.scala 94:16:@35949.4]
  assign RetimeWrapper_101_clock = clock; // @[:@35955.4]
  assign RetimeWrapper_101_reset = reset; // @[:@35956.4]
  assign RetimeWrapper_101_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35958.4]
  assign RetimeWrapper_101_io_in = _T_1535 & io_rPort_8_en_0; // @[package.scala 94:16:@35957.4]
  assign RetimeWrapper_102_clock = clock; // @[:@35963.4]
  assign RetimeWrapper_102_reset = reset; // @[:@35964.4]
  assign RetimeWrapper_102_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35966.4]
  assign RetimeWrapper_102_io_in = _T_1639 & io_rPort_8_en_0; // @[package.scala 94:16:@35965.4]
  assign RetimeWrapper_103_clock = clock; // @[:@35971.4]
  assign RetimeWrapper_103_reset = reset; // @[:@35972.4]
  assign RetimeWrapper_103_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35974.4]
  assign RetimeWrapper_103_io_in = _T_1743 & io_rPort_8_en_0; // @[package.scala 94:16:@35973.4]
  assign RetimeWrapper_104_clock = clock; // @[:@35979.4]
  assign RetimeWrapper_104_reset = reset; // @[:@35980.4]
  assign RetimeWrapper_104_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35982.4]
  assign RetimeWrapper_104_io_in = _T_1847 & io_rPort_8_en_0; // @[package.scala 94:16:@35981.4]
  assign RetimeWrapper_105_clock = clock; // @[:@35987.4]
  assign RetimeWrapper_105_reset = reset; // @[:@35988.4]
  assign RetimeWrapper_105_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35990.4]
  assign RetimeWrapper_105_io_in = _T_1951 & io_rPort_8_en_0; // @[package.scala 94:16:@35989.4]
  assign RetimeWrapper_106_clock = clock; // @[:@35995.4]
  assign RetimeWrapper_106_reset = reset; // @[:@35996.4]
  assign RetimeWrapper_106_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@35998.4]
  assign RetimeWrapper_106_io_in = _T_2055 & io_rPort_8_en_0; // @[package.scala 94:16:@35997.4]
  assign RetimeWrapper_107_clock = clock; // @[:@36003.4]
  assign RetimeWrapper_107_reset = reset; // @[:@36004.4]
  assign RetimeWrapper_107_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@36006.4]
  assign RetimeWrapper_107_io_in = _T_2159 & io_rPort_8_en_0; // @[package.scala 94:16:@36005.4]
  assign RetimeWrapper_108_clock = clock; // @[:@36059.4]
  assign RetimeWrapper_108_reset = reset; // @[:@36060.4]
  assign RetimeWrapper_108_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36062.4]
  assign RetimeWrapper_108_io_in = _T_961 & io_rPort_9_en_0; // @[package.scala 94:16:@36061.4]
  assign RetimeWrapper_109_clock = clock; // @[:@36067.4]
  assign RetimeWrapper_109_reset = reset; // @[:@36068.4]
  assign RetimeWrapper_109_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36070.4]
  assign RetimeWrapper_109_io_in = _T_1065 & io_rPort_9_en_0; // @[package.scala 94:16:@36069.4]
  assign RetimeWrapper_110_clock = clock; // @[:@36075.4]
  assign RetimeWrapper_110_reset = reset; // @[:@36076.4]
  assign RetimeWrapper_110_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36078.4]
  assign RetimeWrapper_110_io_in = _T_1169 & io_rPort_9_en_0; // @[package.scala 94:16:@36077.4]
  assign RetimeWrapper_111_clock = clock; // @[:@36083.4]
  assign RetimeWrapper_111_reset = reset; // @[:@36084.4]
  assign RetimeWrapper_111_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36086.4]
  assign RetimeWrapper_111_io_in = _T_1273 & io_rPort_9_en_0; // @[package.scala 94:16:@36085.4]
  assign RetimeWrapper_112_clock = clock; // @[:@36091.4]
  assign RetimeWrapper_112_reset = reset; // @[:@36092.4]
  assign RetimeWrapper_112_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36094.4]
  assign RetimeWrapper_112_io_in = _T_1377 & io_rPort_9_en_0; // @[package.scala 94:16:@36093.4]
  assign RetimeWrapper_113_clock = clock; // @[:@36099.4]
  assign RetimeWrapper_113_reset = reset; // @[:@36100.4]
  assign RetimeWrapper_113_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36102.4]
  assign RetimeWrapper_113_io_in = _T_1481 & io_rPort_9_en_0; // @[package.scala 94:16:@36101.4]
  assign RetimeWrapper_114_clock = clock; // @[:@36107.4]
  assign RetimeWrapper_114_reset = reset; // @[:@36108.4]
  assign RetimeWrapper_114_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36110.4]
  assign RetimeWrapper_114_io_in = _T_1585 & io_rPort_9_en_0; // @[package.scala 94:16:@36109.4]
  assign RetimeWrapper_115_clock = clock; // @[:@36115.4]
  assign RetimeWrapper_115_reset = reset; // @[:@36116.4]
  assign RetimeWrapper_115_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36118.4]
  assign RetimeWrapper_115_io_in = _T_1689 & io_rPort_9_en_0; // @[package.scala 94:16:@36117.4]
  assign RetimeWrapper_116_clock = clock; // @[:@36123.4]
  assign RetimeWrapper_116_reset = reset; // @[:@36124.4]
  assign RetimeWrapper_116_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36126.4]
  assign RetimeWrapper_116_io_in = _T_1793 & io_rPort_9_en_0; // @[package.scala 94:16:@36125.4]
  assign RetimeWrapper_117_clock = clock; // @[:@36131.4]
  assign RetimeWrapper_117_reset = reset; // @[:@36132.4]
  assign RetimeWrapper_117_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36134.4]
  assign RetimeWrapper_117_io_in = _T_1897 & io_rPort_9_en_0; // @[package.scala 94:16:@36133.4]
  assign RetimeWrapper_118_clock = clock; // @[:@36139.4]
  assign RetimeWrapper_118_reset = reset; // @[:@36140.4]
  assign RetimeWrapper_118_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36142.4]
  assign RetimeWrapper_118_io_in = _T_2001 & io_rPort_9_en_0; // @[package.scala 94:16:@36141.4]
  assign RetimeWrapper_119_clock = clock; // @[:@36147.4]
  assign RetimeWrapper_119_reset = reset; // @[:@36148.4]
  assign RetimeWrapper_119_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@36150.4]
  assign RetimeWrapper_119_io_in = _T_2105 & io_rPort_9_en_0; // @[package.scala 94:16:@36149.4]
endmodule
module Modulo( // @[:@36179.2]
  input         clock, // @[:@36180.4]
  input         io_flow, // @[:@36182.4]
  input  [31:0] io_dividend, // @[:@36182.4]
  input  [31:0] io_divisor, // @[:@36182.4]
  output [31:0] io_out // @[:@36182.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 48:19:@36184.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 48:19:@36184.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 48:19:@36184.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 48:19:@36184.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 48:19:@36184.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 48:19:@36184.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 48:19:@36184.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 48:19:@36184.4]
  div_32_32_16_Unsigned_Remainder m ( // @[ZynqBlackBoxes.scala 48:19:@36184.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign io_out = m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 56:12:@36200.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 54:31:@36198.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 53:32:@36197.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 52:32:@36196.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 51:33:@36195.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 50:17:@36194.4 ZynqBlackBoxes.scala 55:17:@36199.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 49:15:@36193.4]
endmodule
module fix2fixBox_26( // @[:@36202.2]
  input  [63:0] io_a, // @[:@36205.4]
  output [31:0] io_b // @[:@36205.4]
);
  assign io_b = io_a[31:0]; // @[Converter.scala 95:38:@36218.4]
endmodule
module x389( // @[:@36220.2]
  input         clock, // @[:@36221.4]
  input  [31:0] io_a, // @[:@36223.4]
  input         io_flow, // @[:@36223.4]
  output [31:0] io_result // @[:@36223.4]
);
  wire  x389_clock; // @[BigIPZynq.scala 35:21:@36231.4]
  wire  x389_io_flow; // @[BigIPZynq.scala 35:21:@36231.4]
  wire [31:0] x389_io_dividend; // @[BigIPZynq.scala 35:21:@36231.4]
  wire [31:0] x389_io_divisor; // @[BigIPZynq.scala 35:21:@36231.4]
  wire [31:0] x389_io_out; // @[BigIPZynq.scala 35:21:@36231.4]
  wire [63:0] fix2fixBox_io_a; // @[Math.scala 357:30:@36238.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 357:30:@36238.4]
  Modulo x389 ( // @[BigIPZynq.scala 35:21:@36231.4]
    .clock(x389_clock),
    .io_flow(x389_io_flow),
    .io_dividend(x389_io_dividend),
    .io_divisor(x389_io_divisor),
    .io_out(x389_io_out)
  );
  fix2fixBox_26 fix2fixBox ( // @[Math.scala 357:30:@36238.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 363:17:@36246.4]
  assign x389_clock = clock; // @[:@36232.4]
  assign x389_io_flow = io_flow; // @[BigIPZynq.scala 38:17:@36236.4]
  assign x389_io_dividend = io_a; // @[BigIPZynq.scala 36:21:@36234.4]
  assign x389_io_divisor = 32'h6; // @[BigIPZynq.scala 37:20:@36235.4]
  assign fix2fixBox_io_a = {{32'd0}, x389_io_out}; // @[Math.scala 358:23:@36241.4]
endmodule
module Divider( // @[:@36440.2]
  input         clock, // @[:@36441.4]
  input         io_flow, // @[:@36443.4]
  input  [31:0] io_dividend, // @[:@36443.4]
  input  [31:0] io_divisor, // @[:@36443.4]
  output [31:0] io_out // @[:@36443.4]
);
  wire [31:0] m_m_axis_dout_tdata; // @[ZynqBlackBoxes.scala 26:19:@36445.4]
  wire  m_m_axis_dout_tvalid; // @[ZynqBlackBoxes.scala 26:19:@36445.4]
  wire [31:0] m_s_axis_divisor_tdata; // @[ZynqBlackBoxes.scala 26:19:@36445.4]
  wire  m_s_axis_divisor_tvalid; // @[ZynqBlackBoxes.scala 26:19:@36445.4]
  wire [31:0] m_s_axis_dividend_tdata; // @[ZynqBlackBoxes.scala 26:19:@36445.4]
  wire  m_s_axis_dividend_tvalid; // @[ZynqBlackBoxes.scala 26:19:@36445.4]
  wire  m_aclken; // @[ZynqBlackBoxes.scala 26:19:@36445.4]
  wire  m_aclk; // @[ZynqBlackBoxes.scala 26:19:@36445.4]
  wire [29:0] _T_15; // @[ZynqBlackBoxes.scala 34:37:@36461.4]
  div_32_32_20_Signed_Fractional m ( // @[ZynqBlackBoxes.scala 26:19:@36445.4]
    .m_axis_dout_tdata(m_m_axis_dout_tdata),
    .m_axis_dout_tvalid(m_m_axis_dout_tvalid),
    .s_axis_divisor_tdata(m_s_axis_divisor_tdata),
    .s_axis_divisor_tvalid(m_s_axis_divisor_tvalid),
    .s_axis_dividend_tdata(m_s_axis_dividend_tdata),
    .s_axis_dividend_tvalid(m_s_axis_dividend_tvalid),
    .aclken(m_aclken),
    .aclk(m_aclk)
  );
  assign _T_15 = m_m_axis_dout_tdata[31:2]; // @[ZynqBlackBoxes.scala 34:37:@36461.4]
  assign io_out = {{2'd0}, _T_15}; // @[ZynqBlackBoxes.scala 34:12:@36462.4]
  assign m_s_axis_divisor_tdata = io_divisor; // @[ZynqBlackBoxes.scala 32:31:@36459.4]
  assign m_s_axis_divisor_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 31:32:@36458.4]
  assign m_s_axis_dividend_tdata = io_dividend; // @[ZynqBlackBoxes.scala 30:32:@36457.4]
  assign m_s_axis_dividend_tvalid = 1'h1; // @[ZynqBlackBoxes.scala 29:33:@36456.4]
  assign m_aclken = io_flow; // @[ZynqBlackBoxes.scala 28:17:@36455.4 ZynqBlackBoxes.scala 33:17:@36460.4]
  assign m_aclk = clock; // @[ZynqBlackBoxes.scala 27:15:@36454.4]
endmodule
module x392_div( // @[:@36500.2]
  input         clock, // @[:@36501.4]
  input  [31:0] io_a, // @[:@36503.4]
  input         io_flow, // @[:@36503.4]
  output [31:0] io_result // @[:@36503.4]
);
  wire  x392_div_clock; // @[BigIPZynq.scala 25:21:@36511.4]
  wire  x392_div_io_flow; // @[BigIPZynq.scala 25:21:@36511.4]
  wire [31:0] x392_div_io_dividend; // @[BigIPZynq.scala 25:21:@36511.4]
  wire [31:0] x392_div_io_divisor; // @[BigIPZynq.scala 25:21:@36511.4]
  wire [31:0] x392_div_io_out; // @[BigIPZynq.scala 25:21:@36511.4]
  wire [31:0] __io_b; // @[Math.scala 720:24:@36524.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@36524.4]
  wire [31:0] _T_15; // @[FixedPoint.scala 24:59:@36509.4]
  wire [31:0] _T_19; // @[BigIPZynq.scala 29:16:@36519.4]
  Divider x392_div ( // @[BigIPZynq.scala 25:21:@36511.4]
    .clock(x392_div_clock),
    .io_flow(x392_div_io_flow),
    .io_dividend(x392_div_io_dividend),
    .io_divisor(x392_div_io_divisor),
    .io_out(x392_div_io_out)
  );
  _ _ ( // @[Math.scala 720:24:@36524.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  assign _T_15 = $signed(io_a); // @[FixedPoint.scala 24:59:@36509.4]
  assign _T_19 = $signed(x392_div_io_out); // @[BigIPZynq.scala 29:16:@36519.4]
  assign io_result = __io_result; // @[Math.scala 290:34:@36532.4]
  assign x392_div_clock = clock; // @[:@36512.4]
  assign x392_div_io_flow = io_flow; // @[BigIPZynq.scala 28:17:@36518.4]
  assign x392_div_io_dividend = $unsigned(_T_15); // @[BigIPZynq.scala 26:21:@36515.4]
  assign x392_div_io_divisor = 32'h6; // @[BigIPZynq.scala 27:20:@36517.4]
  assign __io_b = $unsigned(_T_19); // @[Math.scala 721:17:@36527.4]
endmodule
module RetimeWrapper_438( // @[:@36546.2]
  input         clock, // @[:@36547.4]
  input         reset, // @[:@36548.4]
  input         io_flow, // @[:@36549.4]
  input  [31:0] io_in, // @[:@36549.4]
  output [31:0] io_out // @[:@36549.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36551.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36551.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36551.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36551.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36551.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36551.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(19)) sr ( // @[RetimeShiftRegister.scala 15:20:@36551.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36564.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36563.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@36562.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36561.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36560.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36558.4]
endmodule
module RetimeWrapper_440( // @[:@36757.2]
  input   clock, // @[:@36758.4]
  input   reset, // @[:@36759.4]
  input   io_flow, // @[:@36760.4]
  input   io_in, // @[:@36760.4]
  output  io_out // @[:@36760.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@36762.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@36762.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@36762.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36762.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36762.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36762.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@36762.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36775.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36774.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@36773.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36772.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36771.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36769.4]
endmodule
module RetimeWrapper_441( // @[:@36789.2]
  input         clock, // @[:@36790.4]
  input         reset, // @[:@36791.4]
  input         io_flow, // @[:@36792.4]
  input  [31:0] io_in, // @[:@36792.4]
  output [31:0] io_out // @[:@36792.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36794.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36794.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36794.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36794.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36794.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36794.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@36794.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36807.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36806.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@36805.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36804.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36803.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36801.4]
endmodule
module RetimeWrapper_443( // @[:@36853.2]
  input         clock, // @[:@36854.4]
  input         reset, // @[:@36855.4]
  input         io_flow, // @[:@36856.4]
  input  [31:0] io_in, // @[:@36856.4]
  output [31:0] io_out // @[:@36856.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36858.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36858.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36858.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36858.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36858.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36858.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@36858.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36871.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36870.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@36869.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36868.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36867.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36865.4]
endmodule
module RetimeWrapper_444( // @[:@36885.2]
  input         clock, // @[:@36886.4]
  input         reset, // @[:@36887.4]
  input         io_flow, // @[:@36888.4]
  input  [31:0] io_in, // @[:@36888.4]
  output [31:0] io_out // @[:@36888.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36890.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36890.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36890.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36890.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36890.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36890.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(23)) sr ( // @[RetimeShiftRegister.scala 15:20:@36890.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36903.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36902.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@36901.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36900.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36899.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36897.4]
endmodule
module RetimeWrapper_445( // @[:@36917.2]
  input         clock, // @[:@36918.4]
  input         reset, // @[:@36919.4]
  input         io_flow, // @[:@36920.4]
  input  [31:0] io_in, // @[:@36920.4]
  output [31:0] io_out // @[:@36920.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@36922.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@36922.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@36922.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@36922.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@36922.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@36922.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(24)) sr ( // @[RetimeShiftRegister.scala 15:20:@36922.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@36935.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@36934.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@36933.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@36932.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@36931.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@36929.4]
endmodule
module RetimeWrapper_448( // @[:@37349.2]
  input         clock, // @[:@37350.4]
  input         reset, // @[:@37351.4]
  input         io_flow, // @[:@37352.4]
  input  [31:0] io_in, // @[:@37352.4]
  output [31:0] io_out // @[:@37352.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@37354.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@37354.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@37354.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@37354.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@37354.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@37354.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@37354.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@37367.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@37366.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@37365.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@37364.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@37363.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@37361.4]
endmodule
module RetimeWrapper_450( // @[:@37560.2]
  input         clock, // @[:@37561.4]
  input         reset, // @[:@37562.4]
  input         io_flow, // @[:@37563.4]
  input  [31:0] io_in, // @[:@37563.4]
  output [31:0] io_out // @[:@37563.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@37565.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@37565.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@37565.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@37565.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@37565.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@37565.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@37565.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@37578.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@37577.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@37576.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@37575.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@37574.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@37572.4]
endmodule
module RetimeWrapper_452( // @[:@37624.2]
  input         clock, // @[:@37625.4]
  input         reset, // @[:@37626.4]
  input         io_flow, // @[:@37627.4]
  input  [31:0] io_in, // @[:@37627.4]
  output [31:0] io_out // @[:@37627.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@37629.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@37629.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@37629.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@37629.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@37629.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@37629.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@37629.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@37642.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@37641.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@37640.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@37639.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@37638.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@37636.4]
endmodule
module RetimeWrapper_466( // @[:@39038.2]
  input         clock, // @[:@39039.4]
  input         reset, // @[:@39040.4]
  input         io_flow, // @[:@39041.4]
  input  [31:0] io_in, // @[:@39041.4]
  output [31:0] io_out // @[:@39041.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@39043.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@39043.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@39043.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39043.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39043.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39043.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(26)) sr ( // @[RetimeShiftRegister.scala 15:20:@39043.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39056.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39055.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@39054.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39053.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39052.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39050.4]
endmodule
module RetimeWrapper_471( // @[:@39198.2]
  input   clock, // @[:@39199.4]
  input   reset, // @[:@39200.4]
  input   io_flow, // @[:@39201.4]
  input   io_in, // @[:@39201.4]
  output  io_out // @[:@39201.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@39203.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@39203.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@39203.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39203.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39203.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39203.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(48)) sr ( // @[RetimeShiftRegister.scala 15:20:@39203.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39216.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39215.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@39214.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39213.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39212.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39210.4]
endmodule
module RetimeWrapper_472( // @[:@39230.2]
  input   clock, // @[:@39231.4]
  input   reset, // @[:@39232.4]
  input   io_flow, // @[:@39233.4]
  input   io_in, // @[:@39233.4]
  output  io_out // @[:@39233.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@39235.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@39235.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@39235.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39235.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39235.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39235.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(20)) sr ( // @[RetimeShiftRegister.scala 15:20:@39235.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39248.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39247.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@39246.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39245.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39244.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39242.4]
endmodule
module RetimeWrapper_475( // @[:@39326.2]
  input         clock, // @[:@39327.4]
  input         reset, // @[:@39328.4]
  input         io_flow, // @[:@39329.4]
  input  [31:0] io_in, // @[:@39329.4]
  output [31:0] io_out // @[:@39329.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@39331.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@39331.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@39331.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39331.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39331.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39331.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(48)) sr ( // @[RetimeShiftRegister.scala 15:20:@39331.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39344.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39343.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@39342.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39341.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39340.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39338.4]
endmodule
module RetimeWrapper_476( // @[:@39358.2]
  input         clock, // @[:@39359.4]
  input         reset, // @[:@39360.4]
  input         io_flow, // @[:@39361.4]
  input  [31:0] io_in, // @[:@39361.4]
  output [31:0] io_out // @[:@39361.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@39363.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@39363.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@39363.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39363.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39363.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39363.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(31)) sr ( // @[RetimeShiftRegister.scala 15:20:@39363.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39376.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39375.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@39374.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39373.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39372.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39370.4]
endmodule
module RetimeWrapper_492( // @[:@39870.2]
  input         clock, // @[:@39871.4]
  input         reset, // @[:@39872.4]
  input         io_flow, // @[:@39873.4]
  input  [31:0] io_in, // @[:@39873.4]
  output [31:0] io_out // @[:@39873.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@39875.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@39875.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@39875.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39875.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39875.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39875.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(32)) sr ( // @[RetimeShiftRegister.scala 15:20:@39875.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39888.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39887.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@39886.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39885.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39884.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39882.4]
endmodule
module RetimeWrapper_493( // @[:@39902.2]
  input         clock, // @[:@39903.4]
  input         reset, // @[:@39904.4]
  input         io_flow, // @[:@39905.4]
  input  [31:0] io_in, // @[:@39905.4]
  output [31:0] io_out // @[:@39905.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@39907.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@39907.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@39907.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39907.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39907.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39907.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(27)) sr ( // @[RetimeShiftRegister.scala 15:20:@39907.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39920.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39919.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@39918.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39917.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39916.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39914.4]
endmodule
module RetimeWrapper_494( // @[:@39934.2]
  input   clock, // @[:@39935.4]
  input   reset, // @[:@39936.4]
  input   io_flow, // @[:@39937.4]
  input   io_in, // @[:@39937.4]
  output  io_out // @[:@39937.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@39939.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@39939.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@39939.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@39939.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@39939.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@39939.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@39939.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@39952.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@39951.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@39950.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@39949.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@39948.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@39946.4]
endmodule
module RetimeWrapper_498( // @[:@40398.2]
  input         clock, // @[:@40399.4]
  input         reset, // @[:@40400.4]
  input         io_flow, // @[:@40401.4]
  input  [31:0] io_in, // @[:@40401.4]
  output [31:0] io_out // @[:@40401.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@40403.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@40403.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@40403.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@40403.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@40403.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@40403.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(46)) sr ( // @[RetimeShiftRegister.scala 15:20:@40403.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@40416.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@40415.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@40414.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@40413.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@40412.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@40410.4]
endmodule
module RetimeWrapper_500( // @[:@40609.2]
  input         clock, // @[:@40610.4]
  input         reset, // @[:@40611.4]
  input         io_flow, // @[:@40612.4]
  input  [31:0] io_in, // @[:@40612.4]
  output [31:0] io_out // @[:@40612.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@40614.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@40614.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@40614.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@40614.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@40614.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@40614.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@40614.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@40627.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@40626.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@40625.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@40624.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@40623.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@40621.4]
endmodule
module RetimeWrapper_515( // @[:@41867.2]
  input         clock, // @[:@41868.4]
  input         reset, // @[:@41869.4]
  input         io_flow, // @[:@41870.4]
  input  [31:0] io_in, // @[:@41870.4]
  output [31:0] io_out // @[:@41870.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@41872.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@41872.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@41872.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@41872.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@41872.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@41872.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(18)) sr ( // @[RetimeShiftRegister.scala 15:20:@41872.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@41885.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@41884.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@41883.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@41882.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@41881.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@41879.4]
endmodule
module RetimeWrapper_530( // @[:@42788.2]
  input         clock, // @[:@42789.4]
  input         reset, // @[:@42790.4]
  input         io_flow, // @[:@42791.4]
  input  [31:0] io_in, // @[:@42791.4]
  output [31:0] io_out // @[:@42791.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@42793.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@42793.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@42793.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@42793.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@42793.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@42793.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(17)) sr ( // @[RetimeShiftRegister.scala 15:20:@42793.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@42806.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@42805.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@42804.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@42803.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@42802.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@42800.4]
endmodule
module Multiplier( // @[:@45620.2]
  input         clock, // @[:@45621.4]
  input         io_flow, // @[:@45623.4]
  input  [31:0] io_a, // @[:@45623.4]
  input  [31:0] io_b, // @[:@45623.4]
  output [31:0] io_out // @[:@45623.4]
);
  wire [31:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@45625.4]
  wire [31:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@45625.4]
  wire [31:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@45625.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@45625.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@45625.4]
  mul_32_32_32_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@45625.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@45635.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@45633.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@45632.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@45634.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@45631.4]
endmodule
module x525( // @[:@45655.2]
  input         clock, // @[:@45656.4]
  input  [31:0] io_a, // @[:@45658.4]
  input  [31:0] io_b, // @[:@45658.4]
  input         io_flow, // @[:@45658.4]
  output [31:0] io_result // @[:@45658.4]
);
  wire  x525_clock; // @[BigIPZynq.scala 63:21:@45665.4]
  wire  x525_io_flow; // @[BigIPZynq.scala 63:21:@45665.4]
  wire [31:0] x525_io_a; // @[BigIPZynq.scala 63:21:@45665.4]
  wire [31:0] x525_io_b; // @[BigIPZynq.scala 63:21:@45665.4]
  wire [31:0] x525_io_out; // @[BigIPZynq.scala 63:21:@45665.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@45674.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@45674.4]
  Multiplier x525 ( // @[BigIPZynq.scala 63:21:@45665.4]
    .clock(x525_clock),
    .io_flow(x525_io_flow),
    .io_a(x525_io_a),
    .io_b(x525_io_b),
    .io_out(x525_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 253:30:@45674.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@45682.4]
  assign x525_clock = clock; // @[:@45666.4]
  assign x525_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@45670.4]
  assign x525_io_a = io_a; // @[BigIPZynq.scala 64:14:@45668.4]
  assign x525_io_b = io_b; // @[BigIPZynq.scala 65:14:@45669.4]
  assign fix2fixBox_io_a = x525_io_out; // @[Math.scala 254:23:@45677.4]
endmodule
module fix2fixBox_131( // @[:@46276.2]
  input  [31:0] io_a, // @[:@46279.4]
  output [32:0] io_b // @[:@46279.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@46293.4]
endmodule
module __78( // @[:@46295.2]
  input  [31:0] io_b, // @[:@46298.4]
  output [32:0] io_result // @[:@46298.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@46303.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@46303.4]
  fix2fixBox_131 fix2fixBox ( // @[BigIPZynq.scala 219:30:@46303.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@46311.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@46306.4]
endmodule
module x534_x7( // @[:@46407.2]
  input         clock, // @[:@46408.4]
  input         reset, // @[:@46409.4]
  input  [31:0] io_a, // @[:@46410.4]
  input  [31:0] io_b, // @[:@46410.4]
  input         io_flow, // @[:@46410.4]
  output [31:0] io_result // @[:@46410.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@46418.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@46418.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@46425.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@46425.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@46435.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@46435.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@46435.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@46435.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@46435.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@46423.4 Math.scala 724:14:@46424.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@46430.4 Math.scala 724:14:@46431.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@46432.4]
  __78 _ ( // @[Math.scala 720:24:@46418.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __78 __1 ( // @[Math.scala 720:24:@46425.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@46435.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@46423.4 Math.scala 724:14:@46424.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@46430.4 Math.scala 724:14:@46431.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@46432.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@46443.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@46421.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@46428.4]
  assign fix2fixBox_clock = clock; // @[:@46436.4]
  assign fix2fixBox_reset = reset; // @[:@46437.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@46438.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@46441.4]
endmodule
module fix2fixBox_155( // @[:@47660.2]
  input  [31:0] io_a, // @[:@47663.4]
  output [31:0] io_b // @[:@47663.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@47673.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@47673.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@47676.4]
endmodule
module x542( // @[:@47678.2]
  input  [31:0] io_b, // @[:@47681.4]
  output [31:0] io_result // @[:@47681.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@47686.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@47686.4]
  fix2fixBox_155 fix2fixBox ( // @[BigIPZynq.scala 219:30:@47686.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@47694.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@47689.4]
endmodule
module Multiplier_9( // @[:@47706.2]
  input         clock, // @[:@47707.4]
  input         io_flow, // @[:@47709.4]
  input  [38:0] io_a, // @[:@47709.4]
  input  [38:0] io_b, // @[:@47709.4]
  output [38:0] io_out // @[:@47709.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@47711.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@47711.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@47711.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@47711.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@47711.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@47711.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@47721.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@47719.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@47718.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@47720.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@47717.4]
endmodule
module fix2fixBox_156( // @[:@47723.2]
  input  [38:0] io_a, // @[:@47726.4]
  output [31:0] io_b // @[:@47726.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@47734.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@47737.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@47734.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@47737.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@47740.4]
endmodule
module x543_mul( // @[:@47742.2]
  input         clock, // @[:@47743.4]
  input  [31:0] io_a, // @[:@47745.4]
  input  [31:0] io_b, // @[:@47745.4]
  input         io_flow, // @[:@47745.4]
  output [31:0] io_result // @[:@47745.4]
);
  wire  x543_mul_clock; // @[BigIPZynq.scala 63:21:@47760.4]
  wire  x543_mul_io_flow; // @[BigIPZynq.scala 63:21:@47760.4]
  wire [38:0] x543_mul_io_a; // @[BigIPZynq.scala 63:21:@47760.4]
  wire [38:0] x543_mul_io_b; // @[BigIPZynq.scala 63:21:@47760.4]
  wire [38:0] x543_mul_io_out; // @[BigIPZynq.scala 63:21:@47760.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@47768.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@47768.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@47752.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@47754.4]
  wire  _T_22; // @[FixedPoint.scala 50:25:@47756.4]
  wire [6:0] _T_26; // @[Bitwise.scala 72:12:@47758.4]
  Multiplier_9 x543_mul ( // @[BigIPZynq.scala 63:21:@47760.4]
    .clock(x543_mul_clock),
    .io_flow(x543_mul_io_flow),
    .io_a(x543_mul_io_a),
    .io_b(x543_mul_io_b),
    .io_out(x543_mul_io_out)
  );
  fix2fixBox_156 fix2fixBox ( // @[Math.scala 253:30:@47768.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@47752.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@47754.4]
  assign _T_22 = io_b[31]; // @[FixedPoint.scala 50:25:@47756.4]
  assign _T_26 = _T_22 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@47758.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@47776.4]
  assign x543_mul_clock = clock; // @[:@47761.4]
  assign x543_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@47765.4]
  assign x543_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@47763.4]
  assign x543_mul_io_b = {_T_26,io_b}; // @[BigIPZynq.scala 65:14:@47764.4]
  assign fix2fixBox_io_a = x543_mul_io_out; // @[Math.scala 254:23:@47771.4]
endmodule
module fix2fixBox_157( // @[:@47778.2]
  input  [31:0] io_a, // @[:@47781.4]
  output [31:0] io_b // @[:@47781.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@47793.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@47793.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@47796.4]
endmodule
module x544( // @[:@47798.2]
  input  [31:0] io_b, // @[:@47801.4]
  output [31:0] io_result // @[:@47801.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@47806.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@47806.4]
  fix2fixBox_157 fix2fixBox ( // @[BigIPZynq.scala 219:30:@47806.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@47814.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@47809.4]
endmodule
module RetimeWrapper_604( // @[:@54002.2]
  input   clock, // @[:@54003.4]
  input   reset, // @[:@54004.4]
  input   io_flow, // @[:@54005.4]
  input   io_in, // @[:@54005.4]
  output  io_out // @[:@54005.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@54007.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@54007.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@54007.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54007.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54007.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54007.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(67)) sr ( // @[RetimeShiftRegister.scala 15:20:@54007.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54020.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54019.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@54018.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54017.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54016.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54014.4]
endmodule
module RetimeWrapper_605( // @[:@54034.2]
  input         clock, // @[:@54035.4]
  input         reset, // @[:@54036.4]
  input         io_flow, // @[:@54037.4]
  input  [31:0] io_in, // @[:@54037.4]
  output [31:0] io_out // @[:@54037.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@54039.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@54039.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@54039.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54039.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54039.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54039.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(51)) sr ( // @[RetimeShiftRegister.scala 15:20:@54039.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54052.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54051.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@54050.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54049.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54048.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54046.4]
endmodule
module RetimeWrapper_609( // @[:@54162.2]
  input         clock, // @[:@54163.4]
  input         reset, // @[:@54164.4]
  input         io_flow, // @[:@54165.4]
  input  [31:0] io_in, // @[:@54165.4]
  output [31:0] io_out // @[:@54165.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@54167.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@54167.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@54167.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54167.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54167.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54167.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(67)) sr ( // @[RetimeShiftRegister.scala 15:20:@54167.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54180.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54179.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@54178.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54177.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54176.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54174.4]
endmodule
module RetimeWrapper_611( // @[:@54226.2]
  input         clock, // @[:@54227.4]
  input         reset, // @[:@54228.4]
  input         io_flow, // @[:@54229.4]
  input  [31:0] io_in, // @[:@54229.4]
  output [31:0] io_out // @[:@54229.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@54231.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@54231.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@54231.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54231.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54231.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54231.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(50)) sr ( // @[RetimeShiftRegister.scala 15:20:@54231.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54244.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54243.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@54242.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54241.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54240.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54238.4]
endmodule
module RetimeWrapper_612( // @[:@54258.2]
  input         clock, // @[:@54259.4]
  input         reset, // @[:@54260.4]
  input         io_flow, // @[:@54261.4]
  input  [31:0] io_in, // @[:@54261.4]
  output [31:0] io_out // @[:@54261.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@54263.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@54263.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@54263.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54263.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54263.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54263.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(45)) sr ( // @[RetimeShiftRegister.scala 15:20:@54263.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54276.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54275.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@54274.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54273.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54272.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54270.4]
endmodule
module RetimeWrapper_623( // @[:@54610.2]
  input   clock, // @[:@54611.4]
  input   reset, // @[:@54612.4]
  input   io_flow, // @[:@54613.4]
  input   io_in, // @[:@54613.4]
  output  io_out // @[:@54613.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@54615.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@54615.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@54615.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54615.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54615.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54615.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(68)) sr ( // @[RetimeShiftRegister.scala 15:20:@54615.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54628.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54627.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@54626.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54625.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54624.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54622.4]
endmodule
module RetimeWrapper_624( // @[:@54642.2]
  input   clock, // @[:@54643.4]
  input   reset, // @[:@54644.4]
  input   io_flow, // @[:@54645.4]
  input   io_in, // @[:@54645.4]
  output  io_out // @[:@54645.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@54647.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@54647.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@54647.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54647.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54647.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54647.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(40)) sr ( // @[RetimeShiftRegister.scala 15:20:@54647.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54660.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54659.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@54658.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54657.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54656.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54654.4]
endmodule
module RetimeWrapper_627( // @[:@54738.2]
  input         clock, // @[:@54739.4]
  input         reset, // @[:@54740.4]
  input         io_flow, // @[:@54741.4]
  input  [31:0] io_in, // @[:@54741.4]
  output [31:0] io_out // @[:@54741.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@54743.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@54743.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@54743.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@54743.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@54743.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@54743.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(68)) sr ( // @[RetimeShiftRegister.scala 15:20:@54743.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@54756.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@54755.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@54754.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@54753.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@54752.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@54750.4]
endmodule
module RetimeWrapper_638( // @[:@55090.2]
  input         clock, // @[:@55091.4]
  input         reset, // @[:@55092.4]
  input         io_flow, // @[:@55093.4]
  input  [31:0] io_in, // @[:@55093.4]
  output [31:0] io_out // @[:@55093.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55095.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55095.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55095.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55095.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55095.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55095.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(52)) sr ( // @[RetimeShiftRegister.scala 15:20:@55095.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55108.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55107.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55106.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@55105.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55104.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55102.4]
endmodule
module RetimeWrapper_639( // @[:@55122.2]
  input         clock, // @[:@55123.4]
  input         reset, // @[:@55124.4]
  input         io_flow, // @[:@55125.4]
  input  [31:0] io_in, // @[:@55125.4]
  output [31:0] io_out // @[:@55125.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55127.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55127.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55127.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55127.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55127.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55127.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(47)) sr ( // @[RetimeShiftRegister.scala 15:20:@55127.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55140.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55139.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55138.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@55137.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55136.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55134.4]
endmodule
module RetimeWrapper_640( // @[:@55154.2]
  input   clock, // @[:@55155.4]
  input   reset, // @[:@55156.4]
  input   io_flow, // @[:@55157.4]
  input   io_in, // @[:@55157.4]
  output  io_out // @[:@55157.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@55159.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@55159.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@55159.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55159.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55159.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55159.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(41)) sr ( // @[RetimeShiftRegister.scala 15:20:@55159.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55172.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55171.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@55170.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@55169.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55168.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55166.4]
endmodule
module RetimeWrapper_642( // @[:@55218.2]
  input         clock, // @[:@55219.4]
  input         reset, // @[:@55220.4]
  input         io_flow, // @[:@55221.4]
  input  [31:0] io_in, // @[:@55221.4]
  output [31:0] io_out // @[:@55221.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55223.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55223.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55223.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55223.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55223.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55223.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(25)) sr ( // @[RetimeShiftRegister.scala 15:20:@55223.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55236.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55235.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55234.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@55233.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55232.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55230.4]
endmodule
module RetimeWrapper_648( // @[:@55410.2]
  input         clock, // @[:@55411.4]
  input         reset, // @[:@55412.4]
  input         io_flow, // @[:@55413.4]
  input  [31:0] io_in, // @[:@55413.4]
  output [31:0] io_out // @[:@55413.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55415.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55415.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55415.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55415.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55415.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55415.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(40)) sr ( // @[RetimeShiftRegister.scala 15:20:@55415.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55428.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55427.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55426.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@55425.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55424.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55422.4]
endmodule
module RetimeWrapper_657( // @[:@55698.2]
  input         clock, // @[:@55699.4]
  input         reset, // @[:@55700.4]
  input         io_flow, // @[:@55701.4]
  input  [31:0] io_in, // @[:@55701.4]
  output [31:0] io_out // @[:@55701.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@55703.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@55703.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@55703.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@55703.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@55703.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@55703.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(21)) sr ( // @[RetimeShiftRegister.scala 15:20:@55703.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@55716.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@55715.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@55714.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@55713.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@55712.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@55710.4]
endmodule
module RetimeWrapper_674( // @[:@59694.2]
  input          clock, // @[:@59695.4]
  input          reset, // @[:@59696.4]
  input          io_flow, // @[:@59697.4]
  input  [127:0] io_in, // @[:@59697.4]
  output [127:0] io_out // @[:@59697.4]
);
  wire [127:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@59699.4]
  wire [127:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@59699.4]
  wire [127:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@59699.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59699.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59699.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59699.4]
  RetimeShiftRegister #(.WIDTH(128), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@59699.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59712.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59711.4]
  assign sr_init = 128'h0; // @[RetimeShiftRegister.scala 19:16:@59710.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59709.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59708.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59706.4]
endmodule
module RetimeWrapper_675( // @[:@59726.2]
  input   clock, // @[:@59727.4]
  input   reset, // @[:@59728.4]
  input   io_flow, // @[:@59729.4]
  input   io_in, // @[:@59729.4]
  output  io_out // @[:@59729.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@59731.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@59731.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@59731.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@59731.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@59731.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@59731.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(87)) sr ( // @[RetimeShiftRegister.scala 15:20:@59731.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@59744.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@59743.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@59742.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@59741.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@59740.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@59738.4]
endmodule
module x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@59810.2]
  input          clock, // @[:@59811.4]
  input          reset, // @[:@59812.4]
  output         io_in_x343_TVALID, // @[:@59813.4]
  input          io_in_x343_TREADY, // @[:@59813.4]
  output [255:0] io_in_x343_TDATA, // @[:@59813.4]
  output         io_in_x342_TREADY, // @[:@59813.4]
  input  [255:0] io_in_x342_TDATA, // @[:@59813.4]
  input  [7:0]   io_in_x342_TID, // @[:@59813.4]
  input  [7:0]   io_in_x342_TDEST, // @[:@59813.4]
  input          io_sigsIn_backpressure, // @[:@59813.4]
  input          io_sigsIn_datapathEn, // @[:@59813.4]
  input          io_sigsIn_break, // @[:@59813.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@59813.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@59813.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@59813.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@59813.4]
  input          io_rr // @[:@59813.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@59827.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@59827.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@59839.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@59839.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@59862.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@59862.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@59862.4]
  wire [127:0] RetimeWrapper_io_in; // @[package.scala 93:22:@59862.4]
  wire [127:0] RetimeWrapper_io_out; // @[package.scala 93:22:@59862.4]
  wire  x383_lb_0_clock; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_reset; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_17_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_17_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_17_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_17_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_17_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_17_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_16_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_16_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_16_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_16_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_16_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_16_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_15_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_15_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_15_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_15_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_15_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_15_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_14_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_14_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_14_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_14_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_14_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_14_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_13_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_13_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_13_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_13_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_13_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_13_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_12_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_12_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_12_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_12_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_12_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_12_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_11_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_11_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_11_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_11_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_11_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_11_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_10_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_10_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_10_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_10_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_10_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_10_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_9_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_9_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_9_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_9_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_9_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_9_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_8_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_8_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_8_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_8_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_8_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_8_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_7_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_7_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_7_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_7_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_7_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_7_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_6_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_6_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_6_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_6_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_6_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_6_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_5_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_5_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_5_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_5_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_5_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_5_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_4_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_4_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_4_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_4_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_4_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_4_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_3_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_3_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_3_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_3_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_3_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_3_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_2_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_2_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_2_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_2_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_2_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_2_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_1_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_1_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_1_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_1_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_1_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_1_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_0_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_rPort_0_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_rPort_0_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_0_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_rPort_0_backpressure; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_rPort_0_output_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_wPort_3_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_wPort_3_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_wPort_3_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_wPort_3_data_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_wPort_3_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_wPort_2_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_wPort_2_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_wPort_2_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_wPort_2_data_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_wPort_2_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_wPort_1_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_wPort_1_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_wPort_1_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_wPort_1_data_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_wPort_1_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_wPort_0_banks_1; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [2:0] x383_lb_0_io_wPort_0_banks_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [8:0] x383_lb_0_io_wPort_0_ofs_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire [31:0] x383_lb_0_io_wPort_0_data_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x383_lb_0_io_wPort_0_en_0; // @[m_x383_lb_0.scala 47:17:@59872.4]
  wire  x384_lb2_0_clock; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_reset; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_9_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_9_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_9_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_9_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_9_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_9_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_8_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_8_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_8_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_8_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_8_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_8_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_7_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_7_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_7_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_7_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_7_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_7_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_6_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_6_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_6_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_6_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_6_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_6_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_5_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_5_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_5_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_5_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_5_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_5_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_4_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_4_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_4_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_4_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_4_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_4_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_3_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_3_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_3_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_3_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_3_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_3_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_2_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_2_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_2_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_2_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_2_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_2_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_1_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_1_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_1_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_1_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_1_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_1_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_0_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_rPort_0_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_rPort_0_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_0_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_rPort_0_backpressure; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_rPort_0_output_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_wPort_3_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_wPort_3_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_wPort_3_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_wPort_3_data_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_wPort_3_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_wPort_2_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_wPort_2_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_wPort_2_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_wPort_2_data_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_wPort_2_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_wPort_1_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_wPort_1_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_wPort_1_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_wPort_1_data_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_wPort_1_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_wPort_0_banks_1; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [2:0] x384_lb2_0_io_wPort_0_banks_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [8:0] x384_lb2_0_io_wPort_0_ofs_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire [31:0] x384_lb2_0_io_wPort_0_data_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x384_lb2_0_io_wPort_0_en_0; // @[m_x384_lb2_0.scala 39:17:@60017.4]
  wire  x389_1_clock; // @[Math.scala 366:24:@60152.4]
  wire [31:0] x389_1_io_a; // @[Math.scala 366:24:@60152.4]
  wire  x389_1_io_flow; // @[Math.scala 366:24:@60152.4]
  wire [31:0] x389_1_io_result; // @[Math.scala 366:24:@60152.4]
  wire  x729_sum_1_clock; // @[Math.scala 150:24:@60189.4]
  wire  x729_sum_1_reset; // @[Math.scala 150:24:@60189.4]
  wire [31:0] x729_sum_1_io_a; // @[Math.scala 150:24:@60189.4]
  wire [31:0] x729_sum_1_io_b; // @[Math.scala 150:24:@60189.4]
  wire  x729_sum_1_io_flow; // @[Math.scala 150:24:@60189.4]
  wire [31:0] x729_sum_1_io_result; // @[Math.scala 150:24:@60189.4]
  wire  x392_div_1_clock; // @[Math.scala 327:24:@60201.4]
  wire [31:0] x392_div_1_io_a; // @[Math.scala 327:24:@60201.4]
  wire  x392_div_1_io_flow; // @[Math.scala 327:24:@60201.4]
  wire [31:0] x392_div_1_io_result; // @[Math.scala 327:24:@60201.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@60211.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@60211.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@60211.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@60211.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@60211.4]
  wire  x393_sum_1_clock; // @[Math.scala 150:24:@60220.4]
  wire  x393_sum_1_reset; // @[Math.scala 150:24:@60220.4]
  wire [31:0] x393_sum_1_io_a; // @[Math.scala 150:24:@60220.4]
  wire [31:0] x393_sum_1_io_b; // @[Math.scala 150:24:@60220.4]
  wire  x393_sum_1_io_flow; // @[Math.scala 150:24:@60220.4]
  wire [31:0] x393_sum_1_io_result; // @[Math.scala 150:24:@60220.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@60230.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@60230.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@60230.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@60230.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@60230.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@60239.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@60239.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@60239.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@60239.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@60239.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@60248.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@60248.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@60248.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@60248.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@60248.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@60257.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@60257.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@60257.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@60257.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@60257.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@60266.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@60266.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@60266.4]
  wire [31:0] RetimeWrapper_6_io_in; // @[package.scala 93:22:@60266.4]
  wire [31:0] RetimeWrapper_6_io_out; // @[package.scala 93:22:@60266.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@60275.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@60275.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@60275.4]
  wire [31:0] RetimeWrapper_7_io_in; // @[package.scala 93:22:@60275.4]
  wire [31:0] RetimeWrapper_7_io_out; // @[package.scala 93:22:@60275.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@60286.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@60286.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@60286.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@60286.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@60286.4]
  wire  x395_rdcol_1_clock; // @[Math.scala 150:24:@60309.4]
  wire  x395_rdcol_1_reset; // @[Math.scala 150:24:@60309.4]
  wire [31:0] x395_rdcol_1_io_a; // @[Math.scala 150:24:@60309.4]
  wire [31:0] x395_rdcol_1_io_b; // @[Math.scala 150:24:@60309.4]
  wire  x395_rdcol_1_io_flow; // @[Math.scala 150:24:@60309.4]
  wire [31:0] x395_rdcol_1_io_result; // @[Math.scala 150:24:@60309.4]
  wire  x397_1_clock; // @[Math.scala 366:24:@60323.4]
  wire [31:0] x397_1_io_a; // @[Math.scala 366:24:@60323.4]
  wire  x397_1_io_flow; // @[Math.scala 366:24:@60323.4]
  wire [31:0] x397_1_io_result; // @[Math.scala 366:24:@60323.4]
  wire  x398_div_1_clock; // @[Math.scala 327:24:@60335.4]
  wire [31:0] x398_div_1_io_a; // @[Math.scala 327:24:@60335.4]
  wire  x398_div_1_io_flow; // @[Math.scala 327:24:@60335.4]
  wire [31:0] x398_div_1_io_result; // @[Math.scala 327:24:@60335.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@60345.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@60345.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@60345.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@60345.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@60345.4]
  wire  x399_sum_1_clock; // @[Math.scala 150:24:@60354.4]
  wire  x399_sum_1_reset; // @[Math.scala 150:24:@60354.4]
  wire [31:0] x399_sum_1_io_a; // @[Math.scala 150:24:@60354.4]
  wire [31:0] x399_sum_1_io_b; // @[Math.scala 150:24:@60354.4]
  wire  x399_sum_1_io_flow; // @[Math.scala 150:24:@60354.4]
  wire [31:0] x399_sum_1_io_result; // @[Math.scala 150:24:@60354.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@60364.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@60364.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@60364.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@60364.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@60364.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@60373.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@60373.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@60373.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@60373.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@60373.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@60382.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@60382.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@60382.4]
  wire [31:0] RetimeWrapper_12_io_in; // @[package.scala 93:22:@60382.4]
  wire [31:0] RetimeWrapper_12_io_out; // @[package.scala 93:22:@60382.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@60393.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@60393.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@60393.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@60393.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@60393.4]
  wire  x401_rdcol_1_clock; // @[Math.scala 150:24:@60416.4]
  wire  x401_rdcol_1_reset; // @[Math.scala 150:24:@60416.4]
  wire [31:0] x401_rdcol_1_io_a; // @[Math.scala 150:24:@60416.4]
  wire [31:0] x401_rdcol_1_io_b; // @[Math.scala 150:24:@60416.4]
  wire  x401_rdcol_1_io_flow; // @[Math.scala 150:24:@60416.4]
  wire [31:0] x401_rdcol_1_io_result; // @[Math.scala 150:24:@60416.4]
  wire  x403_1_clock; // @[Math.scala 366:24:@60430.4]
  wire [31:0] x403_1_io_a; // @[Math.scala 366:24:@60430.4]
  wire  x403_1_io_flow; // @[Math.scala 366:24:@60430.4]
  wire [31:0] x403_1_io_result; // @[Math.scala 366:24:@60430.4]
  wire  x404_div_1_clock; // @[Math.scala 327:24:@60442.4]
  wire [31:0] x404_div_1_io_a; // @[Math.scala 327:24:@60442.4]
  wire  x404_div_1_io_flow; // @[Math.scala 327:24:@60442.4]
  wire [31:0] x404_div_1_io_result; // @[Math.scala 327:24:@60442.4]
  wire  x405_sum_1_clock; // @[Math.scala 150:24:@60452.4]
  wire  x405_sum_1_reset; // @[Math.scala 150:24:@60452.4]
  wire [31:0] x405_sum_1_io_a; // @[Math.scala 150:24:@60452.4]
  wire [31:0] x405_sum_1_io_b; // @[Math.scala 150:24:@60452.4]
  wire  x405_sum_1_io_flow; // @[Math.scala 150:24:@60452.4]
  wire [31:0] x405_sum_1_io_result; // @[Math.scala 150:24:@60452.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@60462.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@60462.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@60462.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@60462.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@60462.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@60471.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@60471.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@60471.4]
  wire [31:0] RetimeWrapper_15_io_in; // @[package.scala 93:22:@60471.4]
  wire [31:0] RetimeWrapper_15_io_out; // @[package.scala 93:22:@60471.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@60480.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@60480.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@60480.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@60480.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@60480.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@60491.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@60491.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@60491.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@60491.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@60491.4]
  wire  x407_rdcol_1_clock; // @[Math.scala 150:24:@60514.4]
  wire  x407_rdcol_1_reset; // @[Math.scala 150:24:@60514.4]
  wire [31:0] x407_rdcol_1_io_a; // @[Math.scala 150:24:@60514.4]
  wire [31:0] x407_rdcol_1_io_b; // @[Math.scala 150:24:@60514.4]
  wire  x407_rdcol_1_io_flow; // @[Math.scala 150:24:@60514.4]
  wire [31:0] x407_rdcol_1_io_result; // @[Math.scala 150:24:@60514.4]
  wire  x409_1_clock; // @[Math.scala 366:24:@60528.4]
  wire [31:0] x409_1_io_a; // @[Math.scala 366:24:@60528.4]
  wire  x409_1_io_flow; // @[Math.scala 366:24:@60528.4]
  wire [31:0] x409_1_io_result; // @[Math.scala 366:24:@60528.4]
  wire  x410_div_1_clock; // @[Math.scala 327:24:@60540.4]
  wire [31:0] x410_div_1_io_a; // @[Math.scala 327:24:@60540.4]
  wire  x410_div_1_io_flow; // @[Math.scala 327:24:@60540.4]
  wire [31:0] x410_div_1_io_result; // @[Math.scala 327:24:@60540.4]
  wire  x411_sum_1_clock; // @[Math.scala 150:24:@60550.4]
  wire  x411_sum_1_reset; // @[Math.scala 150:24:@60550.4]
  wire [31:0] x411_sum_1_io_a; // @[Math.scala 150:24:@60550.4]
  wire [31:0] x411_sum_1_io_b; // @[Math.scala 150:24:@60550.4]
  wire  x411_sum_1_io_flow; // @[Math.scala 150:24:@60550.4]
  wire [31:0] x411_sum_1_io_result; // @[Math.scala 150:24:@60550.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@60560.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@60560.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@60560.4]
  wire [31:0] RetimeWrapper_18_io_in; // @[package.scala 93:22:@60560.4]
  wire [31:0] RetimeWrapper_18_io_out; // @[package.scala 93:22:@60560.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@60569.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@60569.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@60569.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@60569.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@60569.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@60578.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@60578.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@60578.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@60578.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@60578.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@60589.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@60589.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@60589.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@60589.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@60589.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@60610.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@60610.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@60610.4]
  wire [31:0] RetimeWrapper_22_io_in; // @[package.scala 93:22:@60610.4]
  wire [31:0] RetimeWrapper_22_io_out; // @[package.scala 93:22:@60610.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@60626.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@60626.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@60626.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@60626.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@60626.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@60635.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@60635.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@60635.4]
  wire [31:0] RetimeWrapper_24_io_in; // @[package.scala 93:22:@60635.4]
  wire [31:0] RetimeWrapper_24_io_out; // @[package.scala 93:22:@60635.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@60649.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@60649.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@60649.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@60649.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@60649.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@60658.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@60658.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@60658.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@60658.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@60658.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@60673.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@60673.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@60673.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@60673.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@60673.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@60682.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@60682.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@60682.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@60682.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@60682.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@60691.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@60691.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@60691.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@60691.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@60691.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@60700.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@60700.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@60700.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@60700.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@60700.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@60709.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@60709.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@60709.4]
  wire [31:0] RetimeWrapper_31_io_in; // @[package.scala 93:22:@60709.4]
  wire [31:0] RetimeWrapper_31_io_out; // @[package.scala 93:22:@60709.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@60718.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@60718.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@60718.4]
  wire [31:0] RetimeWrapper_32_io_in; // @[package.scala 93:22:@60718.4]
  wire [31:0] RetimeWrapper_32_io_out; // @[package.scala 93:22:@60718.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@60730.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@60730.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@60730.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@60730.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@60730.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@60751.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@60751.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@60751.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@60751.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@60751.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@60765.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@60765.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@60765.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@60765.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@60765.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@60780.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@60780.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@60780.4]
  wire [31:0] RetimeWrapper_36_io_in; // @[package.scala 93:22:@60780.4]
  wire [31:0] RetimeWrapper_36_io_out; // @[package.scala 93:22:@60780.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@60789.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@60789.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@60789.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@60789.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@60789.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@60798.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@60798.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@60798.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@60798.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@60798.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@60810.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@60810.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@60810.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@60810.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@60810.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@60831.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@60831.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@60831.4]
  wire [31:0] RetimeWrapper_40_io_in; // @[package.scala 93:22:@60831.4]
  wire [31:0] RetimeWrapper_40_io_out; // @[package.scala 93:22:@60831.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@60845.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@60845.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@60845.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@60845.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@60845.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@60860.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@60860.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@60860.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@60860.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@60860.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@60869.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@60869.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@60869.4]
  wire [31:0] RetimeWrapper_43_io_in; // @[package.scala 93:22:@60869.4]
  wire [31:0] RetimeWrapper_43_io_out; // @[package.scala 93:22:@60869.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@60878.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@60878.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@60878.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@60878.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@60878.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@60890.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@60890.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@60890.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@60890.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@60890.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@60911.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@60911.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@60911.4]
  wire [31:0] RetimeWrapper_46_io_in; // @[package.scala 93:22:@60911.4]
  wire [31:0] RetimeWrapper_46_io_out; // @[package.scala 93:22:@60911.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@60925.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@60925.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@60925.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@60925.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@60925.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@60940.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@60940.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@60940.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@60940.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@60940.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@60949.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@60949.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@60949.4]
  wire [31:0] RetimeWrapper_49_io_in; // @[package.scala 93:22:@60949.4]
  wire [31:0] RetimeWrapper_49_io_out; // @[package.scala 93:22:@60949.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@60958.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@60970.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@60970.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@60970.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@60970.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@60970.4]
  wire  x435_rdcol_1_clock; // @[Math.scala 150:24:@60993.4]
  wire  x435_rdcol_1_reset; // @[Math.scala 150:24:@60993.4]
  wire [31:0] x435_rdcol_1_io_a; // @[Math.scala 150:24:@60993.4]
  wire [31:0] x435_rdcol_1_io_b; // @[Math.scala 150:24:@60993.4]
  wire  x435_rdcol_1_io_flow; // @[Math.scala 150:24:@60993.4]
  wire [31:0] x435_rdcol_1_io_result; // @[Math.scala 150:24:@60993.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@61008.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@61008.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@61008.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@61008.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@61008.4]
  wire  x439_1_clock; // @[Math.scala 366:24:@61027.4]
  wire [31:0] x439_1_io_a; // @[Math.scala 366:24:@61027.4]
  wire  x439_1_io_flow; // @[Math.scala 366:24:@61027.4]
  wire [31:0] x439_1_io_result; // @[Math.scala 366:24:@61027.4]
  wire  x440_div_1_clock; // @[Math.scala 327:24:@61039.4]
  wire [31:0] x440_div_1_io_a; // @[Math.scala 327:24:@61039.4]
  wire  x440_div_1_io_flow; // @[Math.scala 327:24:@61039.4]
  wire [31:0] x440_div_1_io_result; // @[Math.scala 327:24:@61039.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@61049.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@61049.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@61049.4]
  wire [31:0] RetimeWrapper_53_io_in; // @[package.scala 93:22:@61049.4]
  wire [31:0] RetimeWrapper_53_io_out; // @[package.scala 93:22:@61049.4]
  wire  x441_sum_1_clock; // @[Math.scala 150:24:@61058.4]
  wire  x441_sum_1_reset; // @[Math.scala 150:24:@61058.4]
  wire [31:0] x441_sum_1_io_a; // @[Math.scala 150:24:@61058.4]
  wire [31:0] x441_sum_1_io_b; // @[Math.scala 150:24:@61058.4]
  wire  x441_sum_1_io_flow; // @[Math.scala 150:24:@61058.4]
  wire [31:0] x441_sum_1_io_result; // @[Math.scala 150:24:@61058.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@61068.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@61068.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@61068.4]
  wire [31:0] RetimeWrapper_54_io_in; // @[package.scala 93:22:@61068.4]
  wire [31:0] RetimeWrapper_54_io_out; // @[package.scala 93:22:@61068.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@61077.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@61077.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@61077.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@61077.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@61077.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@61089.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@61089.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@61089.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@61089.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@61089.4]
  wire  x444_rdcol_1_clock; // @[Math.scala 150:24:@61112.4]
  wire  x444_rdcol_1_reset; // @[Math.scala 150:24:@61112.4]
  wire [31:0] x444_rdcol_1_io_a; // @[Math.scala 150:24:@61112.4]
  wire [31:0] x444_rdcol_1_io_b; // @[Math.scala 150:24:@61112.4]
  wire  x444_rdcol_1_io_flow; // @[Math.scala 150:24:@61112.4]
  wire [31:0] x444_rdcol_1_io_result; // @[Math.scala 150:24:@61112.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@61127.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@61127.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@61127.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@61127.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@61127.4]
  wire  x448_1_clock; // @[Math.scala 366:24:@61144.4]
  wire [31:0] x448_1_io_a; // @[Math.scala 366:24:@61144.4]
  wire  x448_1_io_flow; // @[Math.scala 366:24:@61144.4]
  wire [31:0] x448_1_io_result; // @[Math.scala 366:24:@61144.4]
  wire  x449_div_1_clock; // @[Math.scala 327:24:@61156.4]
  wire [31:0] x449_div_1_io_a; // @[Math.scala 327:24:@61156.4]
  wire  x449_div_1_io_flow; // @[Math.scala 327:24:@61156.4]
  wire [31:0] x449_div_1_io_result; // @[Math.scala 327:24:@61156.4]
  wire  x450_sum_1_clock; // @[Math.scala 150:24:@61166.4]
  wire  x450_sum_1_reset; // @[Math.scala 150:24:@61166.4]
  wire [31:0] x450_sum_1_io_a; // @[Math.scala 150:24:@61166.4]
  wire [31:0] x450_sum_1_io_b; // @[Math.scala 150:24:@61166.4]
  wire  x450_sum_1_io_flow; // @[Math.scala 150:24:@61166.4]
  wire [31:0] x450_sum_1_io_result; // @[Math.scala 150:24:@61166.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@61176.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@61176.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@61176.4]
  wire [31:0] RetimeWrapper_58_io_in; // @[package.scala 93:22:@61176.4]
  wire [31:0] RetimeWrapper_58_io_out; // @[package.scala 93:22:@61176.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@61185.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@61185.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@61185.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@61185.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@61185.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@61197.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@61197.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@61197.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@61197.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@61197.4]
  wire  x453_rdrow_1_clock; // @[Math.scala 191:24:@61220.4]
  wire  x453_rdrow_1_reset; // @[Math.scala 191:24:@61220.4]
  wire [31:0] x453_rdrow_1_io_a; // @[Math.scala 191:24:@61220.4]
  wire [31:0] x453_rdrow_1_io_b; // @[Math.scala 191:24:@61220.4]
  wire  x453_rdrow_1_io_flow; // @[Math.scala 191:24:@61220.4]
  wire [31:0] x453_rdrow_1_io_result; // @[Math.scala 191:24:@61220.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@61246.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@61246.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@61246.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@61246.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@61246.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@61268.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@61268.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@61268.4]
  wire [31:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@61268.4]
  wire [31:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@61268.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@61294.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@61294.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@61294.4]
  wire [31:0] RetimeWrapper_63_io_in; // @[package.scala 93:22:@61294.4]
  wire [31:0] RetimeWrapper_63_io_out; // @[package.scala 93:22:@61294.4]
  wire  x734_sum_1_clock; // @[Math.scala 150:24:@61315.4]
  wire  x734_sum_1_reset; // @[Math.scala 150:24:@61315.4]
  wire [31:0] x734_sum_1_io_a; // @[Math.scala 150:24:@61315.4]
  wire [31:0] x734_sum_1_io_b; // @[Math.scala 150:24:@61315.4]
  wire  x734_sum_1_io_flow; // @[Math.scala 150:24:@61315.4]
  wire [31:0] x734_sum_1_io_result; // @[Math.scala 150:24:@61315.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@61325.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@61325.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@61325.4]
  wire [31:0] RetimeWrapper_64_io_in; // @[package.scala 93:22:@61325.4]
  wire [31:0] RetimeWrapper_64_io_out; // @[package.scala 93:22:@61325.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@61334.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@61334.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@61334.4]
  wire [31:0] RetimeWrapper_65_io_in; // @[package.scala 93:22:@61334.4]
  wire [31:0] RetimeWrapper_65_io_out; // @[package.scala 93:22:@61334.4]
  wire  x461_sum_1_clock; // @[Math.scala 150:24:@61343.4]
  wire  x461_sum_1_reset; // @[Math.scala 150:24:@61343.4]
  wire [31:0] x461_sum_1_io_a; // @[Math.scala 150:24:@61343.4]
  wire [31:0] x461_sum_1_io_b; // @[Math.scala 150:24:@61343.4]
  wire  x461_sum_1_io_flow; // @[Math.scala 150:24:@61343.4]
  wire [31:0] x461_sum_1_io_result; // @[Math.scala 150:24:@61343.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@61353.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@61353.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@61353.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@61353.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@61353.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@61362.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@61362.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@61362.4]
  wire [31:0] RetimeWrapper_67_io_in; // @[package.scala 93:22:@61362.4]
  wire [31:0] RetimeWrapper_67_io_out; // @[package.scala 93:22:@61362.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@61374.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@61374.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@61374.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@61374.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@61374.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@61401.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@61401.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@61401.4]
  wire [31:0] RetimeWrapper_69_io_in; // @[package.scala 93:22:@61401.4]
  wire [31:0] RetimeWrapper_69_io_out; // @[package.scala 93:22:@61401.4]
  wire  x466_sum_1_clock; // @[Math.scala 150:24:@61410.4]
  wire  x466_sum_1_reset; // @[Math.scala 150:24:@61410.4]
  wire [31:0] x466_sum_1_io_a; // @[Math.scala 150:24:@61410.4]
  wire [31:0] x466_sum_1_io_b; // @[Math.scala 150:24:@61410.4]
  wire  x466_sum_1_io_flow; // @[Math.scala 150:24:@61410.4]
  wire [31:0] x466_sum_1_io_result; // @[Math.scala 150:24:@61410.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@61420.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@61420.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@61420.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@61420.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@61420.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@61432.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@61432.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@61432.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@61432.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@61432.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@61459.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@61459.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@61459.4]
  wire [31:0] RetimeWrapper_72_io_in; // @[package.scala 93:22:@61459.4]
  wire [31:0] RetimeWrapper_72_io_out; // @[package.scala 93:22:@61459.4]
  wire  x471_sum_1_clock; // @[Math.scala 150:24:@61468.4]
  wire  x471_sum_1_reset; // @[Math.scala 150:24:@61468.4]
  wire [31:0] x471_sum_1_io_a; // @[Math.scala 150:24:@61468.4]
  wire [31:0] x471_sum_1_io_b; // @[Math.scala 150:24:@61468.4]
  wire  x471_sum_1_io_flow; // @[Math.scala 150:24:@61468.4]
  wire [31:0] x471_sum_1_io_result; // @[Math.scala 150:24:@61468.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@61478.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@61478.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@61478.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@61478.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@61478.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@61490.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@61490.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@61490.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@61490.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@61490.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@61511.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@61511.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@61511.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@61511.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@61511.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@61526.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@61526.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@61526.4]
  wire [31:0] RetimeWrapper_76_io_in; // @[package.scala 93:22:@61526.4]
  wire [31:0] RetimeWrapper_76_io_out; // @[package.scala 93:22:@61526.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@61535.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@61535.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@61535.4]
  wire [31:0] RetimeWrapper_77_io_in; // @[package.scala 93:22:@61535.4]
  wire [31:0] RetimeWrapper_77_io_out; // @[package.scala 93:22:@61535.4]
  wire  x476_sum_1_clock; // @[Math.scala 150:24:@61546.4]
  wire  x476_sum_1_reset; // @[Math.scala 150:24:@61546.4]
  wire [31:0] x476_sum_1_io_a; // @[Math.scala 150:24:@61546.4]
  wire [31:0] x476_sum_1_io_b; // @[Math.scala 150:24:@61546.4]
  wire  x476_sum_1_io_flow; // @[Math.scala 150:24:@61546.4]
  wire [31:0] x476_sum_1_io_result; // @[Math.scala 150:24:@61546.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@61556.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@61556.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@61556.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@61556.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@61556.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@61565.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@61565.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@61565.4]
  wire [31:0] RetimeWrapper_79_io_in; // @[package.scala 93:22:@61565.4]
  wire [31:0] RetimeWrapper_79_io_out; // @[package.scala 93:22:@61565.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@61577.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@61577.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@61577.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@61577.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@61577.4]
  wire  x481_sum_1_clock; // @[Math.scala 150:24:@61604.4]
  wire  x481_sum_1_reset; // @[Math.scala 150:24:@61604.4]
  wire [31:0] x481_sum_1_io_a; // @[Math.scala 150:24:@61604.4]
  wire [31:0] x481_sum_1_io_b; // @[Math.scala 150:24:@61604.4]
  wire  x481_sum_1_io_flow; // @[Math.scala 150:24:@61604.4]
  wire [31:0] x481_sum_1_io_result; // @[Math.scala 150:24:@61604.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@61614.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@61614.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@61614.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@61614.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@61614.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@61626.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@61626.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@61626.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@61626.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@61626.4]
  wire  x486_sum_1_clock; // @[Math.scala 150:24:@61653.4]
  wire  x486_sum_1_reset; // @[Math.scala 150:24:@61653.4]
  wire [31:0] x486_sum_1_io_a; // @[Math.scala 150:24:@61653.4]
  wire [31:0] x486_sum_1_io_b; // @[Math.scala 150:24:@61653.4]
  wire  x486_sum_1_io_flow; // @[Math.scala 150:24:@61653.4]
  wire [31:0] x486_sum_1_io_result; // @[Math.scala 150:24:@61653.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@61663.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@61663.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@61663.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@61663.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@61663.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@61675.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@61675.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@61675.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@61675.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@61675.4]
  wire  x489_rdrow_1_clock; // @[Math.scala 191:24:@61698.4]
  wire  x489_rdrow_1_reset; // @[Math.scala 191:24:@61698.4]
  wire [31:0] x489_rdrow_1_io_a; // @[Math.scala 191:24:@61698.4]
  wire [31:0] x489_rdrow_1_io_b; // @[Math.scala 191:24:@61698.4]
  wire  x489_rdrow_1_io_flow; // @[Math.scala 191:24:@61698.4]
  wire [31:0] x489_rdrow_1_io_result; // @[Math.scala 191:24:@61698.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@61724.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@61724.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@61724.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@61724.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@61724.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@61746.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@61746.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@61746.4]
  wire [31:0] RetimeWrapper_86_io_in; // @[package.scala 93:22:@61746.4]
  wire [31:0] RetimeWrapper_86_io_out; // @[package.scala 93:22:@61746.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@61772.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@61772.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@61772.4]
  wire [31:0] RetimeWrapper_87_io_in; // @[package.scala 93:22:@61772.4]
  wire [31:0] RetimeWrapper_87_io_out; // @[package.scala 93:22:@61772.4]
  wire  x739_sum_1_clock; // @[Math.scala 150:24:@61793.4]
  wire  x739_sum_1_reset; // @[Math.scala 150:24:@61793.4]
  wire [31:0] x739_sum_1_io_a; // @[Math.scala 150:24:@61793.4]
  wire [31:0] x739_sum_1_io_b; // @[Math.scala 150:24:@61793.4]
  wire  x739_sum_1_io_flow; // @[Math.scala 150:24:@61793.4]
  wire [31:0] x739_sum_1_io_result; // @[Math.scala 150:24:@61793.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@61803.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@61803.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@61803.4]
  wire [31:0] RetimeWrapper_88_io_in; // @[package.scala 93:22:@61803.4]
  wire [31:0] RetimeWrapper_88_io_out; // @[package.scala 93:22:@61803.4]
  wire  x497_sum_1_clock; // @[Math.scala 150:24:@61812.4]
  wire  x497_sum_1_reset; // @[Math.scala 150:24:@61812.4]
  wire [31:0] x497_sum_1_io_a; // @[Math.scala 150:24:@61812.4]
  wire [31:0] x497_sum_1_io_b; // @[Math.scala 150:24:@61812.4]
  wire  x497_sum_1_io_flow; // @[Math.scala 150:24:@61812.4]
  wire [31:0] x497_sum_1_io_result; // @[Math.scala 150:24:@61812.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@61822.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@61822.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@61822.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@61822.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@61822.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@61831.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@61831.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@61831.4]
  wire [31:0] RetimeWrapper_90_io_in; // @[package.scala 93:22:@61831.4]
  wire [31:0] RetimeWrapper_90_io_out; // @[package.scala 93:22:@61831.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@61843.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@61843.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@61843.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@61843.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@61843.4]
  wire  x502_sum_1_clock; // @[Math.scala 150:24:@61870.4]
  wire  x502_sum_1_reset; // @[Math.scala 150:24:@61870.4]
  wire [31:0] x502_sum_1_io_a; // @[Math.scala 150:24:@61870.4]
  wire [31:0] x502_sum_1_io_b; // @[Math.scala 150:24:@61870.4]
  wire  x502_sum_1_io_flow; // @[Math.scala 150:24:@61870.4]
  wire [31:0] x502_sum_1_io_result; // @[Math.scala 150:24:@61870.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@61880.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@61880.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@61880.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@61880.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@61880.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@61892.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@61892.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@61892.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@61892.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@61892.4]
  wire  x507_sum_1_clock; // @[Math.scala 150:24:@61919.4]
  wire  x507_sum_1_reset; // @[Math.scala 150:24:@61919.4]
  wire [31:0] x507_sum_1_io_a; // @[Math.scala 150:24:@61919.4]
  wire [31:0] x507_sum_1_io_b; // @[Math.scala 150:24:@61919.4]
  wire  x507_sum_1_io_flow; // @[Math.scala 150:24:@61919.4]
  wire [31:0] x507_sum_1_io_result; // @[Math.scala 150:24:@61919.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@61929.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@61929.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@61929.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@61929.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@61929.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@61941.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@61941.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@61941.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@61941.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@61941.4]
  wire  RetimeWrapper_96_clock; // @[package.scala 93:22:@61968.4]
  wire  RetimeWrapper_96_reset; // @[package.scala 93:22:@61968.4]
  wire  RetimeWrapper_96_io_flow; // @[package.scala 93:22:@61968.4]
  wire [31:0] RetimeWrapper_96_io_in; // @[package.scala 93:22:@61968.4]
  wire [31:0] RetimeWrapper_96_io_out; // @[package.scala 93:22:@61968.4]
  wire  x512_sum_1_clock; // @[Math.scala 150:24:@61979.4]
  wire  x512_sum_1_reset; // @[Math.scala 150:24:@61979.4]
  wire [31:0] x512_sum_1_io_a; // @[Math.scala 150:24:@61979.4]
  wire [31:0] x512_sum_1_io_b; // @[Math.scala 150:24:@61979.4]
  wire  x512_sum_1_io_flow; // @[Math.scala 150:24:@61979.4]
  wire [31:0] x512_sum_1_io_result; // @[Math.scala 150:24:@61979.4]
  wire  RetimeWrapper_97_clock; // @[package.scala 93:22:@61989.4]
  wire  RetimeWrapper_97_reset; // @[package.scala 93:22:@61989.4]
  wire  RetimeWrapper_97_io_flow; // @[package.scala 93:22:@61989.4]
  wire  RetimeWrapper_97_io_in; // @[package.scala 93:22:@61989.4]
  wire  RetimeWrapper_97_io_out; // @[package.scala 93:22:@61989.4]
  wire  RetimeWrapper_98_clock; // @[package.scala 93:22:@61998.4]
  wire  RetimeWrapper_98_reset; // @[package.scala 93:22:@61998.4]
  wire  RetimeWrapper_98_io_flow; // @[package.scala 93:22:@61998.4]
  wire [31:0] RetimeWrapper_98_io_in; // @[package.scala 93:22:@61998.4]
  wire [31:0] RetimeWrapper_98_io_out; // @[package.scala 93:22:@61998.4]
  wire  RetimeWrapper_99_clock; // @[package.scala 93:22:@62010.4]
  wire  RetimeWrapper_99_reset; // @[package.scala 93:22:@62010.4]
  wire  RetimeWrapper_99_io_flow; // @[package.scala 93:22:@62010.4]
  wire  RetimeWrapper_99_io_in; // @[package.scala 93:22:@62010.4]
  wire  RetimeWrapper_99_io_out; // @[package.scala 93:22:@62010.4]
  wire  x517_sum_1_clock; // @[Math.scala 150:24:@62037.4]
  wire  x517_sum_1_reset; // @[Math.scala 150:24:@62037.4]
  wire [31:0] x517_sum_1_io_a; // @[Math.scala 150:24:@62037.4]
  wire [31:0] x517_sum_1_io_b; // @[Math.scala 150:24:@62037.4]
  wire  x517_sum_1_io_flow; // @[Math.scala 150:24:@62037.4]
  wire [31:0] x517_sum_1_io_result; // @[Math.scala 150:24:@62037.4]
  wire  RetimeWrapper_100_clock; // @[package.scala 93:22:@62047.4]
  wire  RetimeWrapper_100_reset; // @[package.scala 93:22:@62047.4]
  wire  RetimeWrapper_100_io_flow; // @[package.scala 93:22:@62047.4]
  wire  RetimeWrapper_100_io_in; // @[package.scala 93:22:@62047.4]
  wire  RetimeWrapper_100_io_out; // @[package.scala 93:22:@62047.4]
  wire  RetimeWrapper_101_clock; // @[package.scala 93:22:@62059.4]
  wire  RetimeWrapper_101_reset; // @[package.scala 93:22:@62059.4]
  wire  RetimeWrapper_101_io_flow; // @[package.scala 93:22:@62059.4]
  wire  RetimeWrapper_101_io_in; // @[package.scala 93:22:@62059.4]
  wire  RetimeWrapper_101_io_out; // @[package.scala 93:22:@62059.4]
  wire  x522_sum_1_clock; // @[Math.scala 150:24:@62086.4]
  wire  x522_sum_1_reset; // @[Math.scala 150:24:@62086.4]
  wire [31:0] x522_sum_1_io_a; // @[Math.scala 150:24:@62086.4]
  wire [31:0] x522_sum_1_io_b; // @[Math.scala 150:24:@62086.4]
  wire  x522_sum_1_io_flow; // @[Math.scala 150:24:@62086.4]
  wire [31:0] x522_sum_1_io_result; // @[Math.scala 150:24:@62086.4]
  wire  RetimeWrapper_102_clock; // @[package.scala 93:22:@62096.4]
  wire  RetimeWrapper_102_reset; // @[package.scala 93:22:@62096.4]
  wire  RetimeWrapper_102_io_flow; // @[package.scala 93:22:@62096.4]
  wire  RetimeWrapper_102_io_in; // @[package.scala 93:22:@62096.4]
  wire  RetimeWrapper_102_io_out; // @[package.scala 93:22:@62096.4]
  wire  RetimeWrapper_103_clock; // @[package.scala 93:22:@62108.4]
  wire  RetimeWrapper_103_reset; // @[package.scala 93:22:@62108.4]
  wire  RetimeWrapper_103_io_flow; // @[package.scala 93:22:@62108.4]
  wire  RetimeWrapper_103_io_in; // @[package.scala 93:22:@62108.4]
  wire  RetimeWrapper_103_io_out; // @[package.scala 93:22:@62108.4]
  wire  x525_1_clock; // @[Math.scala 262:24:@62131.4]
  wire [31:0] x525_1_io_a; // @[Math.scala 262:24:@62131.4]
  wire [31:0] x525_1_io_b; // @[Math.scala 262:24:@62131.4]
  wire  x525_1_io_flow; // @[Math.scala 262:24:@62131.4]
  wire [31:0] x525_1_io_result; // @[Math.scala 262:24:@62131.4]
  wire  x526_1_clock; // @[Math.scala 262:24:@62143.4]
  wire [31:0] x526_1_io_a; // @[Math.scala 262:24:@62143.4]
  wire [31:0] x526_1_io_b; // @[Math.scala 262:24:@62143.4]
  wire  x526_1_io_flow; // @[Math.scala 262:24:@62143.4]
  wire [31:0] x526_1_io_result; // @[Math.scala 262:24:@62143.4]
  wire  x527_1_clock; // @[Math.scala 262:24:@62155.4]
  wire [31:0] x527_1_io_a; // @[Math.scala 262:24:@62155.4]
  wire [31:0] x527_1_io_b; // @[Math.scala 262:24:@62155.4]
  wire  x527_1_io_flow; // @[Math.scala 262:24:@62155.4]
  wire [31:0] x527_1_io_result; // @[Math.scala 262:24:@62155.4]
  wire  x528_1_clock; // @[Math.scala 262:24:@62167.4]
  wire [31:0] x528_1_io_a; // @[Math.scala 262:24:@62167.4]
  wire [31:0] x528_1_io_b; // @[Math.scala 262:24:@62167.4]
  wire  x528_1_io_flow; // @[Math.scala 262:24:@62167.4]
  wire [31:0] x528_1_io_result; // @[Math.scala 262:24:@62167.4]
  wire  x529_1_clock; // @[Math.scala 262:24:@62179.4]
  wire [31:0] x529_1_io_a; // @[Math.scala 262:24:@62179.4]
  wire [31:0] x529_1_io_b; // @[Math.scala 262:24:@62179.4]
  wire  x529_1_io_flow; // @[Math.scala 262:24:@62179.4]
  wire [31:0] x529_1_io_result; // @[Math.scala 262:24:@62179.4]
  wire  x530_1_clock; // @[Math.scala 262:24:@62191.4]
  wire [31:0] x530_1_io_a; // @[Math.scala 262:24:@62191.4]
  wire [31:0] x530_1_io_b; // @[Math.scala 262:24:@62191.4]
  wire  x530_1_io_flow; // @[Math.scala 262:24:@62191.4]
  wire [31:0] x530_1_io_result; // @[Math.scala 262:24:@62191.4]
  wire  x531_1_clock; // @[Math.scala 262:24:@62203.4]
  wire [31:0] x531_1_io_a; // @[Math.scala 262:24:@62203.4]
  wire [31:0] x531_1_io_b; // @[Math.scala 262:24:@62203.4]
  wire  x531_1_io_flow; // @[Math.scala 262:24:@62203.4]
  wire [31:0] x531_1_io_result; // @[Math.scala 262:24:@62203.4]
  wire  x532_1_clock; // @[Math.scala 262:24:@62215.4]
  wire [31:0] x532_1_io_a; // @[Math.scala 262:24:@62215.4]
  wire [31:0] x532_1_io_b; // @[Math.scala 262:24:@62215.4]
  wire  x532_1_io_flow; // @[Math.scala 262:24:@62215.4]
  wire [31:0] x532_1_io_result; // @[Math.scala 262:24:@62215.4]
  wire  x533_1_clock; // @[Math.scala 262:24:@62227.4]
  wire [31:0] x533_1_io_a; // @[Math.scala 262:24:@62227.4]
  wire [31:0] x533_1_io_b; // @[Math.scala 262:24:@62227.4]
  wire  x533_1_io_flow; // @[Math.scala 262:24:@62227.4]
  wire [31:0] x533_1_io_result; // @[Math.scala 262:24:@62227.4]
  wire  x534_x7_1_clock; // @[Math.scala 150:24:@62237.4]
  wire  x534_x7_1_reset; // @[Math.scala 150:24:@62237.4]
  wire [31:0] x534_x7_1_io_a; // @[Math.scala 150:24:@62237.4]
  wire [31:0] x534_x7_1_io_b; // @[Math.scala 150:24:@62237.4]
  wire  x534_x7_1_io_flow; // @[Math.scala 150:24:@62237.4]
  wire [31:0] x534_x7_1_io_result; // @[Math.scala 150:24:@62237.4]
  wire  x535_x8_1_clock; // @[Math.scala 150:24:@62247.4]
  wire  x535_x8_1_reset; // @[Math.scala 150:24:@62247.4]
  wire [31:0] x535_x8_1_io_a; // @[Math.scala 150:24:@62247.4]
  wire [31:0] x535_x8_1_io_b; // @[Math.scala 150:24:@62247.4]
  wire  x535_x8_1_io_flow; // @[Math.scala 150:24:@62247.4]
  wire [31:0] x535_x8_1_io_result; // @[Math.scala 150:24:@62247.4]
  wire  x536_x7_1_clock; // @[Math.scala 150:24:@62257.4]
  wire  x536_x7_1_reset; // @[Math.scala 150:24:@62257.4]
  wire [31:0] x536_x7_1_io_a; // @[Math.scala 150:24:@62257.4]
  wire [31:0] x536_x7_1_io_b; // @[Math.scala 150:24:@62257.4]
  wire  x536_x7_1_io_flow; // @[Math.scala 150:24:@62257.4]
  wire [31:0] x536_x7_1_io_result; // @[Math.scala 150:24:@62257.4]
  wire  x537_x8_1_clock; // @[Math.scala 150:24:@62267.4]
  wire  x537_x8_1_reset; // @[Math.scala 150:24:@62267.4]
  wire [31:0] x537_x8_1_io_a; // @[Math.scala 150:24:@62267.4]
  wire [31:0] x537_x8_1_io_b; // @[Math.scala 150:24:@62267.4]
  wire  x537_x8_1_io_flow; // @[Math.scala 150:24:@62267.4]
  wire [31:0] x537_x8_1_io_result; // @[Math.scala 150:24:@62267.4]
  wire  x538_x7_1_clock; // @[Math.scala 150:24:@62277.4]
  wire  x538_x7_1_reset; // @[Math.scala 150:24:@62277.4]
  wire [31:0] x538_x7_1_io_a; // @[Math.scala 150:24:@62277.4]
  wire [31:0] x538_x7_1_io_b; // @[Math.scala 150:24:@62277.4]
  wire  x538_x7_1_io_flow; // @[Math.scala 150:24:@62277.4]
  wire [31:0] x538_x7_1_io_result; // @[Math.scala 150:24:@62277.4]
  wire  x539_x8_1_clock; // @[Math.scala 150:24:@62287.4]
  wire  x539_x8_1_reset; // @[Math.scala 150:24:@62287.4]
  wire [31:0] x539_x8_1_io_a; // @[Math.scala 150:24:@62287.4]
  wire [31:0] x539_x8_1_io_b; // @[Math.scala 150:24:@62287.4]
  wire  x539_x8_1_io_flow; // @[Math.scala 150:24:@62287.4]
  wire [31:0] x539_x8_1_io_result; // @[Math.scala 150:24:@62287.4]
  wire  x540_x7_1_clock; // @[Math.scala 150:24:@62297.4]
  wire  x540_x7_1_reset; // @[Math.scala 150:24:@62297.4]
  wire [31:0] x540_x7_1_io_a; // @[Math.scala 150:24:@62297.4]
  wire [31:0] x540_x7_1_io_b; // @[Math.scala 150:24:@62297.4]
  wire  x540_x7_1_io_flow; // @[Math.scala 150:24:@62297.4]
  wire [31:0] x540_x7_1_io_result; // @[Math.scala 150:24:@62297.4]
  wire  RetimeWrapper_104_clock; // @[package.scala 93:22:@62307.4]
  wire  RetimeWrapper_104_reset; // @[package.scala 93:22:@62307.4]
  wire  RetimeWrapper_104_io_flow; // @[package.scala 93:22:@62307.4]
  wire [31:0] RetimeWrapper_104_io_in; // @[package.scala 93:22:@62307.4]
  wire [31:0] RetimeWrapper_104_io_out; // @[package.scala 93:22:@62307.4]
  wire  x541_sum_1_clock; // @[Math.scala 150:24:@62316.4]
  wire  x541_sum_1_reset; // @[Math.scala 150:24:@62316.4]
  wire [31:0] x541_sum_1_io_a; // @[Math.scala 150:24:@62316.4]
  wire [31:0] x541_sum_1_io_b; // @[Math.scala 150:24:@62316.4]
  wire  x541_sum_1_io_flow; // @[Math.scala 150:24:@62316.4]
  wire [31:0] x541_sum_1_io_result; // @[Math.scala 150:24:@62316.4]
  wire [31:0] x542_1_io_b; // @[Math.scala 720:24:@62326.4]
  wire [31:0] x542_1_io_result; // @[Math.scala 720:24:@62326.4]
  wire  x543_mul_1_clock; // @[Math.scala 262:24:@62337.4]
  wire [31:0] x543_mul_1_io_a; // @[Math.scala 262:24:@62337.4]
  wire [31:0] x543_mul_1_io_b; // @[Math.scala 262:24:@62337.4]
  wire  x543_mul_1_io_flow; // @[Math.scala 262:24:@62337.4]
  wire [31:0] x543_mul_1_io_result; // @[Math.scala 262:24:@62337.4]
  wire [31:0] x544_1_io_b; // @[Math.scala 720:24:@62347.4]
  wire [31:0] x544_1_io_result; // @[Math.scala 720:24:@62347.4]
  wire  x545_1_clock; // @[Math.scala 262:24:@62358.4]
  wire [31:0] x545_1_io_a; // @[Math.scala 262:24:@62358.4]
  wire [31:0] x545_1_io_b; // @[Math.scala 262:24:@62358.4]
  wire  x545_1_io_flow; // @[Math.scala 262:24:@62358.4]
  wire [31:0] x545_1_io_result; // @[Math.scala 262:24:@62358.4]
  wire  x546_1_clock; // @[Math.scala 262:24:@62370.4]
  wire [31:0] x546_1_io_a; // @[Math.scala 262:24:@62370.4]
  wire [31:0] x546_1_io_b; // @[Math.scala 262:24:@62370.4]
  wire  x546_1_io_flow; // @[Math.scala 262:24:@62370.4]
  wire [31:0] x546_1_io_result; // @[Math.scala 262:24:@62370.4]
  wire  x547_1_clock; // @[Math.scala 262:24:@62382.4]
  wire [31:0] x547_1_io_a; // @[Math.scala 262:24:@62382.4]
  wire [31:0] x547_1_io_b; // @[Math.scala 262:24:@62382.4]
  wire  x547_1_io_flow; // @[Math.scala 262:24:@62382.4]
  wire [31:0] x547_1_io_result; // @[Math.scala 262:24:@62382.4]
  wire  x548_1_clock; // @[Math.scala 262:24:@62394.4]
  wire [31:0] x548_1_io_a; // @[Math.scala 262:24:@62394.4]
  wire [31:0] x548_1_io_b; // @[Math.scala 262:24:@62394.4]
  wire  x548_1_io_flow; // @[Math.scala 262:24:@62394.4]
  wire [31:0] x548_1_io_result; // @[Math.scala 262:24:@62394.4]
  wire  x549_1_clock; // @[Math.scala 262:24:@62406.4]
  wire [31:0] x549_1_io_a; // @[Math.scala 262:24:@62406.4]
  wire [31:0] x549_1_io_b; // @[Math.scala 262:24:@62406.4]
  wire  x549_1_io_flow; // @[Math.scala 262:24:@62406.4]
  wire [31:0] x549_1_io_result; // @[Math.scala 262:24:@62406.4]
  wire  x550_1_clock; // @[Math.scala 262:24:@62420.4]
  wire [31:0] x550_1_io_a; // @[Math.scala 262:24:@62420.4]
  wire [31:0] x550_1_io_b; // @[Math.scala 262:24:@62420.4]
  wire  x550_1_io_flow; // @[Math.scala 262:24:@62420.4]
  wire [31:0] x550_1_io_result; // @[Math.scala 262:24:@62420.4]
  wire  x551_1_clock; // @[Math.scala 262:24:@62432.4]
  wire [31:0] x551_1_io_a; // @[Math.scala 262:24:@62432.4]
  wire [31:0] x551_1_io_b; // @[Math.scala 262:24:@62432.4]
  wire  x551_1_io_flow; // @[Math.scala 262:24:@62432.4]
  wire [31:0] x551_1_io_result; // @[Math.scala 262:24:@62432.4]
  wire  x552_1_clock; // @[Math.scala 262:24:@62444.4]
  wire [31:0] x552_1_io_a; // @[Math.scala 262:24:@62444.4]
  wire [31:0] x552_1_io_b; // @[Math.scala 262:24:@62444.4]
  wire  x552_1_io_flow; // @[Math.scala 262:24:@62444.4]
  wire [31:0] x552_1_io_result; // @[Math.scala 262:24:@62444.4]
  wire  x553_1_clock; // @[Math.scala 262:24:@62456.4]
  wire [31:0] x553_1_io_a; // @[Math.scala 262:24:@62456.4]
  wire [31:0] x553_1_io_b; // @[Math.scala 262:24:@62456.4]
  wire  x553_1_io_flow; // @[Math.scala 262:24:@62456.4]
  wire [31:0] x553_1_io_result; // @[Math.scala 262:24:@62456.4]
  wire  x554_x7_1_clock; // @[Math.scala 150:24:@62466.4]
  wire  x554_x7_1_reset; // @[Math.scala 150:24:@62466.4]
  wire [31:0] x554_x7_1_io_a; // @[Math.scala 150:24:@62466.4]
  wire [31:0] x554_x7_1_io_b; // @[Math.scala 150:24:@62466.4]
  wire  x554_x7_1_io_flow; // @[Math.scala 150:24:@62466.4]
  wire [31:0] x554_x7_1_io_result; // @[Math.scala 150:24:@62466.4]
  wire  x555_x8_1_clock; // @[Math.scala 150:24:@62476.4]
  wire  x555_x8_1_reset; // @[Math.scala 150:24:@62476.4]
  wire [31:0] x555_x8_1_io_a; // @[Math.scala 150:24:@62476.4]
  wire [31:0] x555_x8_1_io_b; // @[Math.scala 150:24:@62476.4]
  wire  x555_x8_1_io_flow; // @[Math.scala 150:24:@62476.4]
  wire [31:0] x555_x8_1_io_result; // @[Math.scala 150:24:@62476.4]
  wire  x556_x7_1_clock; // @[Math.scala 150:24:@62486.4]
  wire  x556_x7_1_reset; // @[Math.scala 150:24:@62486.4]
  wire [31:0] x556_x7_1_io_a; // @[Math.scala 150:24:@62486.4]
  wire [31:0] x556_x7_1_io_b; // @[Math.scala 150:24:@62486.4]
  wire  x556_x7_1_io_flow; // @[Math.scala 150:24:@62486.4]
  wire [31:0] x556_x7_1_io_result; // @[Math.scala 150:24:@62486.4]
  wire  x557_x8_1_clock; // @[Math.scala 150:24:@62496.4]
  wire  x557_x8_1_reset; // @[Math.scala 150:24:@62496.4]
  wire [31:0] x557_x8_1_io_a; // @[Math.scala 150:24:@62496.4]
  wire [31:0] x557_x8_1_io_b; // @[Math.scala 150:24:@62496.4]
  wire  x557_x8_1_io_flow; // @[Math.scala 150:24:@62496.4]
  wire [31:0] x557_x8_1_io_result; // @[Math.scala 150:24:@62496.4]
  wire  x558_x7_1_clock; // @[Math.scala 150:24:@62506.4]
  wire  x558_x7_1_reset; // @[Math.scala 150:24:@62506.4]
  wire [31:0] x558_x7_1_io_a; // @[Math.scala 150:24:@62506.4]
  wire [31:0] x558_x7_1_io_b; // @[Math.scala 150:24:@62506.4]
  wire  x558_x7_1_io_flow; // @[Math.scala 150:24:@62506.4]
  wire [31:0] x558_x7_1_io_result; // @[Math.scala 150:24:@62506.4]
  wire  x559_x8_1_clock; // @[Math.scala 150:24:@62516.4]
  wire  x559_x8_1_reset; // @[Math.scala 150:24:@62516.4]
  wire [31:0] x559_x8_1_io_a; // @[Math.scala 150:24:@62516.4]
  wire [31:0] x559_x8_1_io_b; // @[Math.scala 150:24:@62516.4]
  wire  x559_x8_1_io_flow; // @[Math.scala 150:24:@62516.4]
  wire [31:0] x559_x8_1_io_result; // @[Math.scala 150:24:@62516.4]
  wire  x560_x7_1_clock; // @[Math.scala 150:24:@62526.4]
  wire  x560_x7_1_reset; // @[Math.scala 150:24:@62526.4]
  wire [31:0] x560_x7_1_io_a; // @[Math.scala 150:24:@62526.4]
  wire [31:0] x560_x7_1_io_b; // @[Math.scala 150:24:@62526.4]
  wire  x560_x7_1_io_flow; // @[Math.scala 150:24:@62526.4]
  wire [31:0] x560_x7_1_io_result; // @[Math.scala 150:24:@62526.4]
  wire  RetimeWrapper_105_clock; // @[package.scala 93:22:@62536.4]
  wire  RetimeWrapper_105_reset; // @[package.scala 93:22:@62536.4]
  wire  RetimeWrapper_105_io_flow; // @[package.scala 93:22:@62536.4]
  wire [31:0] RetimeWrapper_105_io_in; // @[package.scala 93:22:@62536.4]
  wire [31:0] RetimeWrapper_105_io_out; // @[package.scala 93:22:@62536.4]
  wire  x561_sum_1_clock; // @[Math.scala 150:24:@62545.4]
  wire  x561_sum_1_reset; // @[Math.scala 150:24:@62545.4]
  wire [31:0] x561_sum_1_io_a; // @[Math.scala 150:24:@62545.4]
  wire [31:0] x561_sum_1_io_b; // @[Math.scala 150:24:@62545.4]
  wire  x561_sum_1_io_flow; // @[Math.scala 150:24:@62545.4]
  wire [31:0] x561_sum_1_io_result; // @[Math.scala 150:24:@62545.4]
  wire [31:0] x562_1_io_b; // @[Math.scala 720:24:@62555.4]
  wire [31:0] x562_1_io_result; // @[Math.scala 720:24:@62555.4]
  wire  x563_mul_1_clock; // @[Math.scala 262:24:@62566.4]
  wire [31:0] x563_mul_1_io_a; // @[Math.scala 262:24:@62566.4]
  wire [31:0] x563_mul_1_io_b; // @[Math.scala 262:24:@62566.4]
  wire  x563_mul_1_io_flow; // @[Math.scala 262:24:@62566.4]
  wire [31:0] x563_mul_1_io_result; // @[Math.scala 262:24:@62566.4]
  wire [31:0] x564_1_io_b; // @[Math.scala 720:24:@62576.4]
  wire [31:0] x564_1_io_result; // @[Math.scala 720:24:@62576.4]
  wire  x565_1_clock; // @[Math.scala 262:24:@62587.4]
  wire [31:0] x565_1_io_a; // @[Math.scala 262:24:@62587.4]
  wire [31:0] x565_1_io_b; // @[Math.scala 262:24:@62587.4]
  wire  x565_1_io_flow; // @[Math.scala 262:24:@62587.4]
  wire [31:0] x565_1_io_result; // @[Math.scala 262:24:@62587.4]
  wire  x566_1_clock; // @[Math.scala 262:24:@62599.4]
  wire [31:0] x566_1_io_a; // @[Math.scala 262:24:@62599.4]
  wire [31:0] x566_1_io_b; // @[Math.scala 262:24:@62599.4]
  wire  x566_1_io_flow; // @[Math.scala 262:24:@62599.4]
  wire [31:0] x566_1_io_result; // @[Math.scala 262:24:@62599.4]
  wire  x567_1_clock; // @[Math.scala 262:24:@62611.4]
  wire [31:0] x567_1_io_a; // @[Math.scala 262:24:@62611.4]
  wire [31:0] x567_1_io_b; // @[Math.scala 262:24:@62611.4]
  wire  x567_1_io_flow; // @[Math.scala 262:24:@62611.4]
  wire [31:0] x567_1_io_result; // @[Math.scala 262:24:@62611.4]
  wire  x568_1_clock; // @[Math.scala 262:24:@62623.4]
  wire [31:0] x568_1_io_a; // @[Math.scala 262:24:@62623.4]
  wire [31:0] x568_1_io_b; // @[Math.scala 262:24:@62623.4]
  wire  x568_1_io_flow; // @[Math.scala 262:24:@62623.4]
  wire [31:0] x568_1_io_result; // @[Math.scala 262:24:@62623.4]
  wire  x569_1_clock; // @[Math.scala 262:24:@62635.4]
  wire [31:0] x569_1_io_a; // @[Math.scala 262:24:@62635.4]
  wire [31:0] x569_1_io_b; // @[Math.scala 262:24:@62635.4]
  wire  x569_1_io_flow; // @[Math.scala 262:24:@62635.4]
  wire [31:0] x569_1_io_result; // @[Math.scala 262:24:@62635.4]
  wire  x570_1_clock; // @[Math.scala 262:24:@62647.4]
  wire [31:0] x570_1_io_a; // @[Math.scala 262:24:@62647.4]
  wire [31:0] x570_1_io_b; // @[Math.scala 262:24:@62647.4]
  wire  x570_1_io_flow; // @[Math.scala 262:24:@62647.4]
  wire [31:0] x570_1_io_result; // @[Math.scala 262:24:@62647.4]
  wire  x571_x7_1_clock; // @[Math.scala 150:24:@62657.4]
  wire  x571_x7_1_reset; // @[Math.scala 150:24:@62657.4]
  wire [31:0] x571_x7_1_io_a; // @[Math.scala 150:24:@62657.4]
  wire [31:0] x571_x7_1_io_b; // @[Math.scala 150:24:@62657.4]
  wire  x571_x7_1_io_flow; // @[Math.scala 150:24:@62657.4]
  wire [31:0] x571_x7_1_io_result; // @[Math.scala 150:24:@62657.4]
  wire  x572_x8_1_clock; // @[Math.scala 150:24:@62667.4]
  wire  x572_x8_1_reset; // @[Math.scala 150:24:@62667.4]
  wire [31:0] x572_x8_1_io_a; // @[Math.scala 150:24:@62667.4]
  wire [31:0] x572_x8_1_io_b; // @[Math.scala 150:24:@62667.4]
  wire  x572_x8_1_io_flow; // @[Math.scala 150:24:@62667.4]
  wire [31:0] x572_x8_1_io_result; // @[Math.scala 150:24:@62667.4]
  wire  x573_x7_1_clock; // @[Math.scala 150:24:@62677.4]
  wire  x573_x7_1_reset; // @[Math.scala 150:24:@62677.4]
  wire [31:0] x573_x7_1_io_a; // @[Math.scala 150:24:@62677.4]
  wire [31:0] x573_x7_1_io_b; // @[Math.scala 150:24:@62677.4]
  wire  x573_x7_1_io_flow; // @[Math.scala 150:24:@62677.4]
  wire [31:0] x573_x7_1_io_result; // @[Math.scala 150:24:@62677.4]
  wire  x574_x8_1_clock; // @[Math.scala 150:24:@62687.4]
  wire  x574_x8_1_reset; // @[Math.scala 150:24:@62687.4]
  wire [31:0] x574_x8_1_io_a; // @[Math.scala 150:24:@62687.4]
  wire [31:0] x574_x8_1_io_b; // @[Math.scala 150:24:@62687.4]
  wire  x574_x8_1_io_flow; // @[Math.scala 150:24:@62687.4]
  wire [31:0] x574_x8_1_io_result; // @[Math.scala 150:24:@62687.4]
  wire  x575_x7_1_clock; // @[Math.scala 150:24:@62697.4]
  wire  x575_x7_1_reset; // @[Math.scala 150:24:@62697.4]
  wire [31:0] x575_x7_1_io_a; // @[Math.scala 150:24:@62697.4]
  wire [31:0] x575_x7_1_io_b; // @[Math.scala 150:24:@62697.4]
  wire  x575_x7_1_io_flow; // @[Math.scala 150:24:@62697.4]
  wire [31:0] x575_x7_1_io_result; // @[Math.scala 150:24:@62697.4]
  wire  x576_x8_1_clock; // @[Math.scala 150:24:@62707.4]
  wire  x576_x8_1_reset; // @[Math.scala 150:24:@62707.4]
  wire [31:0] x576_x8_1_io_a; // @[Math.scala 150:24:@62707.4]
  wire [31:0] x576_x8_1_io_b; // @[Math.scala 150:24:@62707.4]
  wire  x576_x8_1_io_flow; // @[Math.scala 150:24:@62707.4]
  wire [31:0] x576_x8_1_io_result; // @[Math.scala 150:24:@62707.4]
  wire  x577_x7_1_clock; // @[Math.scala 150:24:@62717.4]
  wire  x577_x7_1_reset; // @[Math.scala 150:24:@62717.4]
  wire [31:0] x577_x7_1_io_a; // @[Math.scala 150:24:@62717.4]
  wire [31:0] x577_x7_1_io_b; // @[Math.scala 150:24:@62717.4]
  wire  x577_x7_1_io_flow; // @[Math.scala 150:24:@62717.4]
  wire [31:0] x577_x7_1_io_result; // @[Math.scala 150:24:@62717.4]
  wire  RetimeWrapper_106_clock; // @[package.scala 93:22:@62727.4]
  wire  RetimeWrapper_106_reset; // @[package.scala 93:22:@62727.4]
  wire  RetimeWrapper_106_io_flow; // @[package.scala 93:22:@62727.4]
  wire [31:0] RetimeWrapper_106_io_in; // @[package.scala 93:22:@62727.4]
  wire [31:0] RetimeWrapper_106_io_out; // @[package.scala 93:22:@62727.4]
  wire  x578_sum_1_clock; // @[Math.scala 150:24:@62736.4]
  wire  x578_sum_1_reset; // @[Math.scala 150:24:@62736.4]
  wire [31:0] x578_sum_1_io_a; // @[Math.scala 150:24:@62736.4]
  wire [31:0] x578_sum_1_io_b; // @[Math.scala 150:24:@62736.4]
  wire  x578_sum_1_io_flow; // @[Math.scala 150:24:@62736.4]
  wire [31:0] x578_sum_1_io_result; // @[Math.scala 150:24:@62736.4]
  wire [31:0] x579_1_io_b; // @[Math.scala 720:24:@62746.4]
  wire [31:0] x579_1_io_result; // @[Math.scala 720:24:@62746.4]
  wire  x580_mul_1_clock; // @[Math.scala 262:24:@62757.4]
  wire [31:0] x580_mul_1_io_a; // @[Math.scala 262:24:@62757.4]
  wire [31:0] x580_mul_1_io_b; // @[Math.scala 262:24:@62757.4]
  wire  x580_mul_1_io_flow; // @[Math.scala 262:24:@62757.4]
  wire [31:0] x580_mul_1_io_result; // @[Math.scala 262:24:@62757.4]
  wire [31:0] x581_1_io_b; // @[Math.scala 720:24:@62767.4]
  wire [31:0] x581_1_io_result; // @[Math.scala 720:24:@62767.4]
  wire  x582_1_clock; // @[Math.scala 262:24:@62778.4]
  wire [31:0] x582_1_io_a; // @[Math.scala 262:24:@62778.4]
  wire [31:0] x582_1_io_b; // @[Math.scala 262:24:@62778.4]
  wire  x582_1_io_flow; // @[Math.scala 262:24:@62778.4]
  wire [31:0] x582_1_io_result; // @[Math.scala 262:24:@62778.4]
  wire  x583_1_clock; // @[Math.scala 262:24:@62790.4]
  wire [31:0] x583_1_io_a; // @[Math.scala 262:24:@62790.4]
  wire [31:0] x583_1_io_b; // @[Math.scala 262:24:@62790.4]
  wire  x583_1_io_flow; // @[Math.scala 262:24:@62790.4]
  wire [31:0] x583_1_io_result; // @[Math.scala 262:24:@62790.4]
  wire  x584_1_clock; // @[Math.scala 262:24:@62802.4]
  wire [31:0] x584_1_io_a; // @[Math.scala 262:24:@62802.4]
  wire [31:0] x584_1_io_b; // @[Math.scala 262:24:@62802.4]
  wire  x584_1_io_flow; // @[Math.scala 262:24:@62802.4]
  wire [31:0] x584_1_io_result; // @[Math.scala 262:24:@62802.4]
  wire  x585_1_clock; // @[Math.scala 262:24:@62814.4]
  wire [31:0] x585_1_io_a; // @[Math.scala 262:24:@62814.4]
  wire [31:0] x585_1_io_b; // @[Math.scala 262:24:@62814.4]
  wire  x585_1_io_flow; // @[Math.scala 262:24:@62814.4]
  wire [31:0] x585_1_io_result; // @[Math.scala 262:24:@62814.4]
  wire  x586_1_clock; // @[Math.scala 262:24:@62826.4]
  wire [31:0] x586_1_io_a; // @[Math.scala 262:24:@62826.4]
  wire [31:0] x586_1_io_b; // @[Math.scala 262:24:@62826.4]
  wire  x586_1_io_flow; // @[Math.scala 262:24:@62826.4]
  wire [31:0] x586_1_io_result; // @[Math.scala 262:24:@62826.4]
  wire  x587_1_clock; // @[Math.scala 262:24:@62838.4]
  wire [31:0] x587_1_io_a; // @[Math.scala 262:24:@62838.4]
  wire [31:0] x587_1_io_b; // @[Math.scala 262:24:@62838.4]
  wire  x587_1_io_flow; // @[Math.scala 262:24:@62838.4]
  wire [31:0] x587_1_io_result; // @[Math.scala 262:24:@62838.4]
  wire  x588_x7_1_clock; // @[Math.scala 150:24:@62848.4]
  wire  x588_x7_1_reset; // @[Math.scala 150:24:@62848.4]
  wire [31:0] x588_x7_1_io_a; // @[Math.scala 150:24:@62848.4]
  wire [31:0] x588_x7_1_io_b; // @[Math.scala 150:24:@62848.4]
  wire  x588_x7_1_io_flow; // @[Math.scala 150:24:@62848.4]
  wire [31:0] x588_x7_1_io_result; // @[Math.scala 150:24:@62848.4]
  wire  x589_x8_1_clock; // @[Math.scala 150:24:@62858.4]
  wire  x589_x8_1_reset; // @[Math.scala 150:24:@62858.4]
  wire [31:0] x589_x8_1_io_a; // @[Math.scala 150:24:@62858.4]
  wire [31:0] x589_x8_1_io_b; // @[Math.scala 150:24:@62858.4]
  wire  x589_x8_1_io_flow; // @[Math.scala 150:24:@62858.4]
  wire [31:0] x589_x8_1_io_result; // @[Math.scala 150:24:@62858.4]
  wire  x590_x7_1_clock; // @[Math.scala 150:24:@62868.4]
  wire  x590_x7_1_reset; // @[Math.scala 150:24:@62868.4]
  wire [31:0] x590_x7_1_io_a; // @[Math.scala 150:24:@62868.4]
  wire [31:0] x590_x7_1_io_b; // @[Math.scala 150:24:@62868.4]
  wire  x590_x7_1_io_flow; // @[Math.scala 150:24:@62868.4]
  wire [31:0] x590_x7_1_io_result; // @[Math.scala 150:24:@62868.4]
  wire  x591_x8_1_clock; // @[Math.scala 150:24:@62878.4]
  wire  x591_x8_1_reset; // @[Math.scala 150:24:@62878.4]
  wire [31:0] x591_x8_1_io_a; // @[Math.scala 150:24:@62878.4]
  wire [31:0] x591_x8_1_io_b; // @[Math.scala 150:24:@62878.4]
  wire  x591_x8_1_io_flow; // @[Math.scala 150:24:@62878.4]
  wire [31:0] x591_x8_1_io_result; // @[Math.scala 150:24:@62878.4]
  wire  x592_x7_1_clock; // @[Math.scala 150:24:@62888.4]
  wire  x592_x7_1_reset; // @[Math.scala 150:24:@62888.4]
  wire [31:0] x592_x7_1_io_a; // @[Math.scala 150:24:@62888.4]
  wire [31:0] x592_x7_1_io_b; // @[Math.scala 150:24:@62888.4]
  wire  x592_x7_1_io_flow; // @[Math.scala 150:24:@62888.4]
  wire [31:0] x592_x7_1_io_result; // @[Math.scala 150:24:@62888.4]
  wire  x593_x8_1_clock; // @[Math.scala 150:24:@62898.4]
  wire  x593_x8_1_reset; // @[Math.scala 150:24:@62898.4]
  wire [31:0] x593_x8_1_io_a; // @[Math.scala 150:24:@62898.4]
  wire [31:0] x593_x8_1_io_b; // @[Math.scala 150:24:@62898.4]
  wire  x593_x8_1_io_flow; // @[Math.scala 150:24:@62898.4]
  wire [31:0] x593_x8_1_io_result; // @[Math.scala 150:24:@62898.4]
  wire  x594_x7_1_clock; // @[Math.scala 150:24:@62908.4]
  wire  x594_x7_1_reset; // @[Math.scala 150:24:@62908.4]
  wire [31:0] x594_x7_1_io_a; // @[Math.scala 150:24:@62908.4]
  wire [31:0] x594_x7_1_io_b; // @[Math.scala 150:24:@62908.4]
  wire  x594_x7_1_io_flow; // @[Math.scala 150:24:@62908.4]
  wire [31:0] x594_x7_1_io_result; // @[Math.scala 150:24:@62908.4]
  wire  RetimeWrapper_107_clock; // @[package.scala 93:22:@62918.4]
  wire  RetimeWrapper_107_reset; // @[package.scala 93:22:@62918.4]
  wire  RetimeWrapper_107_io_flow; // @[package.scala 93:22:@62918.4]
  wire [31:0] RetimeWrapper_107_io_in; // @[package.scala 93:22:@62918.4]
  wire [31:0] RetimeWrapper_107_io_out; // @[package.scala 93:22:@62918.4]
  wire  x595_sum_1_clock; // @[Math.scala 150:24:@62927.4]
  wire  x595_sum_1_reset; // @[Math.scala 150:24:@62927.4]
  wire [31:0] x595_sum_1_io_a; // @[Math.scala 150:24:@62927.4]
  wire [31:0] x595_sum_1_io_b; // @[Math.scala 150:24:@62927.4]
  wire  x595_sum_1_io_flow; // @[Math.scala 150:24:@62927.4]
  wire [31:0] x595_sum_1_io_result; // @[Math.scala 150:24:@62927.4]
  wire [31:0] x596_1_io_b; // @[Math.scala 720:24:@62939.4]
  wire [31:0] x596_1_io_result; // @[Math.scala 720:24:@62939.4]
  wire  x597_mul_1_clock; // @[Math.scala 262:24:@62950.4]
  wire [31:0] x597_mul_1_io_a; // @[Math.scala 262:24:@62950.4]
  wire [31:0] x597_mul_1_io_b; // @[Math.scala 262:24:@62950.4]
  wire  x597_mul_1_io_flow; // @[Math.scala 262:24:@62950.4]
  wire [31:0] x597_mul_1_io_result; // @[Math.scala 262:24:@62950.4]
  wire [31:0] x598_1_io_b; // @[Math.scala 720:24:@62960.4]
  wire [31:0] x598_1_io_result; // @[Math.scala 720:24:@62960.4]
  wire  RetimeWrapper_108_clock; // @[package.scala 93:22:@62969.4]
  wire  RetimeWrapper_108_reset; // @[package.scala 93:22:@62969.4]
  wire  RetimeWrapper_108_io_flow; // @[package.scala 93:22:@62969.4]
  wire  RetimeWrapper_108_io_in; // @[package.scala 93:22:@62969.4]
  wire  RetimeWrapper_108_io_out; // @[package.scala 93:22:@62969.4]
  wire  RetimeWrapper_109_clock; // @[package.scala 93:22:@62978.4]
  wire  RetimeWrapper_109_reset; // @[package.scala 93:22:@62978.4]
  wire  RetimeWrapper_109_io_flow; // @[package.scala 93:22:@62978.4]
  wire [31:0] RetimeWrapper_109_io_in; // @[package.scala 93:22:@62978.4]
  wire [31:0] RetimeWrapper_109_io_out; // @[package.scala 93:22:@62978.4]
  wire  RetimeWrapper_110_clock; // @[package.scala 93:22:@62987.4]
  wire  RetimeWrapper_110_reset; // @[package.scala 93:22:@62987.4]
  wire  RetimeWrapper_110_io_flow; // @[package.scala 93:22:@62987.4]
  wire  RetimeWrapper_110_io_in; // @[package.scala 93:22:@62987.4]
  wire  RetimeWrapper_110_io_out; // @[package.scala 93:22:@62987.4]
  wire  RetimeWrapper_111_clock; // @[package.scala 93:22:@62996.4]
  wire  RetimeWrapper_111_reset; // @[package.scala 93:22:@62996.4]
  wire  RetimeWrapper_111_io_flow; // @[package.scala 93:22:@62996.4]
  wire [31:0] RetimeWrapper_111_io_in; // @[package.scala 93:22:@62996.4]
  wire [31:0] RetimeWrapper_111_io_out; // @[package.scala 93:22:@62996.4]
  wire  RetimeWrapper_112_clock; // @[package.scala 93:22:@63005.4]
  wire  RetimeWrapper_112_reset; // @[package.scala 93:22:@63005.4]
  wire  RetimeWrapper_112_io_flow; // @[package.scala 93:22:@63005.4]
  wire [31:0] RetimeWrapper_112_io_in; // @[package.scala 93:22:@63005.4]
  wire [31:0] RetimeWrapper_112_io_out; // @[package.scala 93:22:@63005.4]
  wire  RetimeWrapper_113_clock; // @[package.scala 93:22:@63014.4]
  wire  RetimeWrapper_113_reset; // @[package.scala 93:22:@63014.4]
  wire  RetimeWrapper_113_io_flow; // @[package.scala 93:22:@63014.4]
  wire [31:0] RetimeWrapper_113_io_in; // @[package.scala 93:22:@63014.4]
  wire [31:0] RetimeWrapper_113_io_out; // @[package.scala 93:22:@63014.4]
  wire  RetimeWrapper_114_clock; // @[package.scala 93:22:@63025.4]
  wire  RetimeWrapper_114_reset; // @[package.scala 93:22:@63025.4]
  wire  RetimeWrapper_114_io_flow; // @[package.scala 93:22:@63025.4]
  wire  RetimeWrapper_114_io_in; // @[package.scala 93:22:@63025.4]
  wire  RetimeWrapper_114_io_out; // @[package.scala 93:22:@63025.4]
  wire  RetimeWrapper_115_clock; // @[package.scala 93:22:@63046.4]
  wire  RetimeWrapper_115_reset; // @[package.scala 93:22:@63046.4]
  wire  RetimeWrapper_115_io_flow; // @[package.scala 93:22:@63046.4]
  wire [31:0] RetimeWrapper_115_io_in; // @[package.scala 93:22:@63046.4]
  wire [31:0] RetimeWrapper_115_io_out; // @[package.scala 93:22:@63046.4]
  wire  RetimeWrapper_116_clock; // @[package.scala 93:22:@63055.4]
  wire  RetimeWrapper_116_reset; // @[package.scala 93:22:@63055.4]
  wire  RetimeWrapper_116_io_flow; // @[package.scala 93:22:@63055.4]
  wire [31:0] RetimeWrapper_116_io_in; // @[package.scala 93:22:@63055.4]
  wire [31:0] RetimeWrapper_116_io_out; // @[package.scala 93:22:@63055.4]
  wire  RetimeWrapper_117_clock; // @[package.scala 93:22:@63064.4]
  wire  RetimeWrapper_117_reset; // @[package.scala 93:22:@63064.4]
  wire  RetimeWrapper_117_io_flow; // @[package.scala 93:22:@63064.4]
  wire [31:0] RetimeWrapper_117_io_in; // @[package.scala 93:22:@63064.4]
  wire [31:0] RetimeWrapper_117_io_out; // @[package.scala 93:22:@63064.4]
  wire  RetimeWrapper_118_clock; // @[package.scala 93:22:@63075.4]
  wire  RetimeWrapper_118_reset; // @[package.scala 93:22:@63075.4]
  wire  RetimeWrapper_118_io_flow; // @[package.scala 93:22:@63075.4]
  wire  RetimeWrapper_118_io_in; // @[package.scala 93:22:@63075.4]
  wire  RetimeWrapper_118_io_out; // @[package.scala 93:22:@63075.4]
  wire  RetimeWrapper_119_clock; // @[package.scala 93:22:@63096.4]
  wire  RetimeWrapper_119_reset; // @[package.scala 93:22:@63096.4]
  wire  RetimeWrapper_119_io_flow; // @[package.scala 93:22:@63096.4]
  wire [31:0] RetimeWrapper_119_io_in; // @[package.scala 93:22:@63096.4]
  wire [31:0] RetimeWrapper_119_io_out; // @[package.scala 93:22:@63096.4]
  wire  RetimeWrapper_120_clock; // @[package.scala 93:22:@63105.4]
  wire  RetimeWrapper_120_reset; // @[package.scala 93:22:@63105.4]
  wire  RetimeWrapper_120_io_flow; // @[package.scala 93:22:@63105.4]
  wire [31:0] RetimeWrapper_120_io_in; // @[package.scala 93:22:@63105.4]
  wire [31:0] RetimeWrapper_120_io_out; // @[package.scala 93:22:@63105.4]
  wire  RetimeWrapper_121_clock; // @[package.scala 93:22:@63114.4]
  wire  RetimeWrapper_121_reset; // @[package.scala 93:22:@63114.4]
  wire  RetimeWrapper_121_io_flow; // @[package.scala 93:22:@63114.4]
  wire [31:0] RetimeWrapper_121_io_in; // @[package.scala 93:22:@63114.4]
  wire [31:0] RetimeWrapper_121_io_out; // @[package.scala 93:22:@63114.4]
  wire  RetimeWrapper_122_clock; // @[package.scala 93:22:@63125.4]
  wire  RetimeWrapper_122_reset; // @[package.scala 93:22:@63125.4]
  wire  RetimeWrapper_122_io_flow; // @[package.scala 93:22:@63125.4]
  wire  RetimeWrapper_122_io_in; // @[package.scala 93:22:@63125.4]
  wire  RetimeWrapper_122_io_out; // @[package.scala 93:22:@63125.4]
  wire  RetimeWrapper_123_clock; // @[package.scala 93:22:@63146.4]
  wire  RetimeWrapper_123_reset; // @[package.scala 93:22:@63146.4]
  wire  RetimeWrapper_123_io_flow; // @[package.scala 93:22:@63146.4]
  wire [31:0] RetimeWrapper_123_io_in; // @[package.scala 93:22:@63146.4]
  wire [31:0] RetimeWrapper_123_io_out; // @[package.scala 93:22:@63146.4]
  wire  RetimeWrapper_124_clock; // @[package.scala 93:22:@63155.4]
  wire  RetimeWrapper_124_reset; // @[package.scala 93:22:@63155.4]
  wire  RetimeWrapper_124_io_flow; // @[package.scala 93:22:@63155.4]
  wire [31:0] RetimeWrapper_124_io_in; // @[package.scala 93:22:@63155.4]
  wire [31:0] RetimeWrapper_124_io_out; // @[package.scala 93:22:@63155.4]
  wire  RetimeWrapper_125_clock; // @[package.scala 93:22:@63164.4]
  wire  RetimeWrapper_125_reset; // @[package.scala 93:22:@63164.4]
  wire  RetimeWrapper_125_io_flow; // @[package.scala 93:22:@63164.4]
  wire [31:0] RetimeWrapper_125_io_in; // @[package.scala 93:22:@63164.4]
  wire [31:0] RetimeWrapper_125_io_out; // @[package.scala 93:22:@63164.4]
  wire  RetimeWrapper_126_clock; // @[package.scala 93:22:@63175.4]
  wire  RetimeWrapper_126_reset; // @[package.scala 93:22:@63175.4]
  wire  RetimeWrapper_126_io_flow; // @[package.scala 93:22:@63175.4]
  wire  RetimeWrapper_126_io_in; // @[package.scala 93:22:@63175.4]
  wire  RetimeWrapper_126_io_out; // @[package.scala 93:22:@63175.4]
  wire  RetimeWrapper_127_clock; // @[package.scala 93:22:@63196.4]
  wire  RetimeWrapper_127_reset; // @[package.scala 93:22:@63196.4]
  wire  RetimeWrapper_127_io_flow; // @[package.scala 93:22:@63196.4]
  wire  RetimeWrapper_127_io_in; // @[package.scala 93:22:@63196.4]
  wire  RetimeWrapper_127_io_out; // @[package.scala 93:22:@63196.4]
  wire  RetimeWrapper_128_clock; // @[package.scala 93:22:@63205.4]
  wire  RetimeWrapper_128_reset; // @[package.scala 93:22:@63205.4]
  wire  RetimeWrapper_128_io_flow; // @[package.scala 93:22:@63205.4]
  wire  RetimeWrapper_128_io_in; // @[package.scala 93:22:@63205.4]
  wire  RetimeWrapper_128_io_out; // @[package.scala 93:22:@63205.4]
  wire  RetimeWrapper_129_clock; // @[package.scala 93:22:@63214.4]
  wire  RetimeWrapper_129_reset; // @[package.scala 93:22:@63214.4]
  wire  RetimeWrapper_129_io_flow; // @[package.scala 93:22:@63214.4]
  wire [31:0] RetimeWrapper_129_io_in; // @[package.scala 93:22:@63214.4]
  wire [31:0] RetimeWrapper_129_io_out; // @[package.scala 93:22:@63214.4]
  wire  RetimeWrapper_130_clock; // @[package.scala 93:22:@63223.4]
  wire  RetimeWrapper_130_reset; // @[package.scala 93:22:@63223.4]
  wire  RetimeWrapper_130_io_flow; // @[package.scala 93:22:@63223.4]
  wire  RetimeWrapper_130_io_in; // @[package.scala 93:22:@63223.4]
  wire  RetimeWrapper_130_io_out; // @[package.scala 93:22:@63223.4]
  wire  RetimeWrapper_131_clock; // @[package.scala 93:22:@63232.4]
  wire  RetimeWrapper_131_reset; // @[package.scala 93:22:@63232.4]
  wire  RetimeWrapper_131_io_flow; // @[package.scala 93:22:@63232.4]
  wire [31:0] RetimeWrapper_131_io_in; // @[package.scala 93:22:@63232.4]
  wire [31:0] RetimeWrapper_131_io_out; // @[package.scala 93:22:@63232.4]
  wire  RetimeWrapper_132_clock; // @[package.scala 93:22:@63241.4]
  wire  RetimeWrapper_132_reset; // @[package.scala 93:22:@63241.4]
  wire  RetimeWrapper_132_io_flow; // @[package.scala 93:22:@63241.4]
  wire [31:0] RetimeWrapper_132_io_in; // @[package.scala 93:22:@63241.4]
  wire [31:0] RetimeWrapper_132_io_out; // @[package.scala 93:22:@63241.4]
  wire  RetimeWrapper_133_clock; // @[package.scala 93:22:@63253.4]
  wire  RetimeWrapper_133_reset; // @[package.scala 93:22:@63253.4]
  wire  RetimeWrapper_133_io_flow; // @[package.scala 93:22:@63253.4]
  wire  RetimeWrapper_133_io_in; // @[package.scala 93:22:@63253.4]
  wire  RetimeWrapper_133_io_out; // @[package.scala 93:22:@63253.4]
  wire  RetimeWrapper_134_clock; // @[package.scala 93:22:@63274.4]
  wire  RetimeWrapper_134_reset; // @[package.scala 93:22:@63274.4]
  wire  RetimeWrapper_134_io_flow; // @[package.scala 93:22:@63274.4]
  wire [31:0] RetimeWrapper_134_io_in; // @[package.scala 93:22:@63274.4]
  wire [31:0] RetimeWrapper_134_io_out; // @[package.scala 93:22:@63274.4]
  wire  RetimeWrapper_135_clock; // @[package.scala 93:22:@63283.4]
  wire  RetimeWrapper_135_reset; // @[package.scala 93:22:@63283.4]
  wire  RetimeWrapper_135_io_flow; // @[package.scala 93:22:@63283.4]
  wire [31:0] RetimeWrapper_135_io_in; // @[package.scala 93:22:@63283.4]
  wire [31:0] RetimeWrapper_135_io_out; // @[package.scala 93:22:@63283.4]
  wire  RetimeWrapper_136_clock; // @[package.scala 93:22:@63292.4]
  wire  RetimeWrapper_136_reset; // @[package.scala 93:22:@63292.4]
  wire  RetimeWrapper_136_io_flow; // @[package.scala 93:22:@63292.4]
  wire  RetimeWrapper_136_io_in; // @[package.scala 93:22:@63292.4]
  wire  RetimeWrapper_136_io_out; // @[package.scala 93:22:@63292.4]
  wire  RetimeWrapper_137_clock; // @[package.scala 93:22:@63304.4]
  wire  RetimeWrapper_137_reset; // @[package.scala 93:22:@63304.4]
  wire  RetimeWrapper_137_io_flow; // @[package.scala 93:22:@63304.4]
  wire  RetimeWrapper_137_io_in; // @[package.scala 93:22:@63304.4]
  wire  RetimeWrapper_137_io_out; // @[package.scala 93:22:@63304.4]
  wire  RetimeWrapper_138_clock; // @[package.scala 93:22:@63325.4]
  wire  RetimeWrapper_138_reset; // @[package.scala 93:22:@63325.4]
  wire  RetimeWrapper_138_io_flow; // @[package.scala 93:22:@63325.4]
  wire [31:0] RetimeWrapper_138_io_in; // @[package.scala 93:22:@63325.4]
  wire [31:0] RetimeWrapper_138_io_out; // @[package.scala 93:22:@63325.4]
  wire  RetimeWrapper_139_clock; // @[package.scala 93:22:@63334.4]
  wire  RetimeWrapper_139_reset; // @[package.scala 93:22:@63334.4]
  wire  RetimeWrapper_139_io_flow; // @[package.scala 93:22:@63334.4]
  wire [31:0] RetimeWrapper_139_io_in; // @[package.scala 93:22:@63334.4]
  wire [31:0] RetimeWrapper_139_io_out; // @[package.scala 93:22:@63334.4]
  wire  RetimeWrapper_140_clock; // @[package.scala 93:22:@63343.4]
  wire  RetimeWrapper_140_reset; // @[package.scala 93:22:@63343.4]
  wire  RetimeWrapper_140_io_flow; // @[package.scala 93:22:@63343.4]
  wire  RetimeWrapper_140_io_in; // @[package.scala 93:22:@63343.4]
  wire  RetimeWrapper_140_io_out; // @[package.scala 93:22:@63343.4]
  wire  RetimeWrapper_141_clock; // @[package.scala 93:22:@63355.4]
  wire  RetimeWrapper_141_reset; // @[package.scala 93:22:@63355.4]
  wire  RetimeWrapper_141_io_flow; // @[package.scala 93:22:@63355.4]
  wire  RetimeWrapper_141_io_in; // @[package.scala 93:22:@63355.4]
  wire  RetimeWrapper_141_io_out; // @[package.scala 93:22:@63355.4]
  wire  RetimeWrapper_142_clock; // @[package.scala 93:22:@63376.4]
  wire  RetimeWrapper_142_reset; // @[package.scala 93:22:@63376.4]
  wire  RetimeWrapper_142_io_flow; // @[package.scala 93:22:@63376.4]
  wire [31:0] RetimeWrapper_142_io_in; // @[package.scala 93:22:@63376.4]
  wire [31:0] RetimeWrapper_142_io_out; // @[package.scala 93:22:@63376.4]
  wire  RetimeWrapper_143_clock; // @[package.scala 93:22:@63385.4]
  wire  RetimeWrapper_143_reset; // @[package.scala 93:22:@63385.4]
  wire  RetimeWrapper_143_io_flow; // @[package.scala 93:22:@63385.4]
  wire [31:0] RetimeWrapper_143_io_in; // @[package.scala 93:22:@63385.4]
  wire [31:0] RetimeWrapper_143_io_out; // @[package.scala 93:22:@63385.4]
  wire  RetimeWrapper_144_clock; // @[package.scala 93:22:@63394.4]
  wire  RetimeWrapper_144_reset; // @[package.scala 93:22:@63394.4]
  wire  RetimeWrapper_144_io_flow; // @[package.scala 93:22:@63394.4]
  wire  RetimeWrapper_144_io_in; // @[package.scala 93:22:@63394.4]
  wire  RetimeWrapper_144_io_out; // @[package.scala 93:22:@63394.4]
  wire  RetimeWrapper_145_clock; // @[package.scala 93:22:@63406.4]
  wire  RetimeWrapper_145_reset; // @[package.scala 93:22:@63406.4]
  wire  RetimeWrapper_145_io_flow; // @[package.scala 93:22:@63406.4]
  wire  RetimeWrapper_145_io_in; // @[package.scala 93:22:@63406.4]
  wire  RetimeWrapper_145_io_out; // @[package.scala 93:22:@63406.4]
  wire  RetimeWrapper_146_clock; // @[package.scala 93:22:@63427.4]
  wire  RetimeWrapper_146_reset; // @[package.scala 93:22:@63427.4]
  wire  RetimeWrapper_146_io_flow; // @[package.scala 93:22:@63427.4]
  wire [31:0] RetimeWrapper_146_io_in; // @[package.scala 93:22:@63427.4]
  wire [31:0] RetimeWrapper_146_io_out; // @[package.scala 93:22:@63427.4]
  wire  RetimeWrapper_147_clock; // @[package.scala 93:22:@63436.4]
  wire  RetimeWrapper_147_reset; // @[package.scala 93:22:@63436.4]
  wire  RetimeWrapper_147_io_flow; // @[package.scala 93:22:@63436.4]
  wire  RetimeWrapper_147_io_in; // @[package.scala 93:22:@63436.4]
  wire  RetimeWrapper_147_io_out; // @[package.scala 93:22:@63436.4]
  wire  RetimeWrapper_148_clock; // @[package.scala 93:22:@63445.4]
  wire  RetimeWrapper_148_reset; // @[package.scala 93:22:@63445.4]
  wire  RetimeWrapper_148_io_flow; // @[package.scala 93:22:@63445.4]
  wire [31:0] RetimeWrapper_148_io_in; // @[package.scala 93:22:@63445.4]
  wire [31:0] RetimeWrapper_148_io_out; // @[package.scala 93:22:@63445.4]
  wire  RetimeWrapper_149_clock; // @[package.scala 93:22:@63457.4]
  wire  RetimeWrapper_149_reset; // @[package.scala 93:22:@63457.4]
  wire  RetimeWrapper_149_io_flow; // @[package.scala 93:22:@63457.4]
  wire  RetimeWrapper_149_io_in; // @[package.scala 93:22:@63457.4]
  wire  RetimeWrapper_149_io_out; // @[package.scala 93:22:@63457.4]
  wire  RetimeWrapper_150_clock; // @[package.scala 93:22:@63478.4]
  wire  RetimeWrapper_150_reset; // @[package.scala 93:22:@63478.4]
  wire  RetimeWrapper_150_io_flow; // @[package.scala 93:22:@63478.4]
  wire [31:0] RetimeWrapper_150_io_in; // @[package.scala 93:22:@63478.4]
  wire [31:0] RetimeWrapper_150_io_out; // @[package.scala 93:22:@63478.4]
  wire  RetimeWrapper_151_clock; // @[package.scala 93:22:@63487.4]
  wire  RetimeWrapper_151_reset; // @[package.scala 93:22:@63487.4]
  wire  RetimeWrapper_151_io_flow; // @[package.scala 93:22:@63487.4]
  wire  RetimeWrapper_151_io_in; // @[package.scala 93:22:@63487.4]
  wire  RetimeWrapper_151_io_out; // @[package.scala 93:22:@63487.4]
  wire  RetimeWrapper_152_clock; // @[package.scala 93:22:@63496.4]
  wire  RetimeWrapper_152_reset; // @[package.scala 93:22:@63496.4]
  wire  RetimeWrapper_152_io_flow; // @[package.scala 93:22:@63496.4]
  wire [31:0] RetimeWrapper_152_io_in; // @[package.scala 93:22:@63496.4]
  wire [31:0] RetimeWrapper_152_io_out; // @[package.scala 93:22:@63496.4]
  wire  RetimeWrapper_153_clock; // @[package.scala 93:22:@63508.4]
  wire  RetimeWrapper_153_reset; // @[package.scala 93:22:@63508.4]
  wire  RetimeWrapper_153_io_flow; // @[package.scala 93:22:@63508.4]
  wire  RetimeWrapper_153_io_in; // @[package.scala 93:22:@63508.4]
  wire  RetimeWrapper_153_io_out; // @[package.scala 93:22:@63508.4]
  wire  RetimeWrapper_154_clock; // @[package.scala 93:22:@63529.4]
  wire  RetimeWrapper_154_reset; // @[package.scala 93:22:@63529.4]
  wire  RetimeWrapper_154_io_flow; // @[package.scala 93:22:@63529.4]
  wire [31:0] RetimeWrapper_154_io_in; // @[package.scala 93:22:@63529.4]
  wire [31:0] RetimeWrapper_154_io_out; // @[package.scala 93:22:@63529.4]
  wire  RetimeWrapper_155_clock; // @[package.scala 93:22:@63538.4]
  wire  RetimeWrapper_155_reset; // @[package.scala 93:22:@63538.4]
  wire  RetimeWrapper_155_io_flow; // @[package.scala 93:22:@63538.4]
  wire  RetimeWrapper_155_io_in; // @[package.scala 93:22:@63538.4]
  wire  RetimeWrapper_155_io_out; // @[package.scala 93:22:@63538.4]
  wire  RetimeWrapper_156_clock; // @[package.scala 93:22:@63550.4]
  wire  RetimeWrapper_156_reset; // @[package.scala 93:22:@63550.4]
  wire  RetimeWrapper_156_io_flow; // @[package.scala 93:22:@63550.4]
  wire  RetimeWrapper_156_io_in; // @[package.scala 93:22:@63550.4]
  wire  RetimeWrapper_156_io_out; // @[package.scala 93:22:@63550.4]
  wire  RetimeWrapper_157_clock; // @[package.scala 93:22:@63571.4]
  wire  RetimeWrapper_157_reset; // @[package.scala 93:22:@63571.4]
  wire  RetimeWrapper_157_io_flow; // @[package.scala 93:22:@63571.4]
  wire [31:0] RetimeWrapper_157_io_in; // @[package.scala 93:22:@63571.4]
  wire [31:0] RetimeWrapper_157_io_out; // @[package.scala 93:22:@63571.4]
  wire  RetimeWrapper_158_clock; // @[package.scala 93:22:@63580.4]
  wire  RetimeWrapper_158_reset; // @[package.scala 93:22:@63580.4]
  wire  RetimeWrapper_158_io_flow; // @[package.scala 93:22:@63580.4]
  wire  RetimeWrapper_158_io_in; // @[package.scala 93:22:@63580.4]
  wire  RetimeWrapper_158_io_out; // @[package.scala 93:22:@63580.4]
  wire  RetimeWrapper_159_clock; // @[package.scala 93:22:@63592.4]
  wire  RetimeWrapper_159_reset; // @[package.scala 93:22:@63592.4]
  wire  RetimeWrapper_159_io_flow; // @[package.scala 93:22:@63592.4]
  wire  RetimeWrapper_159_io_in; // @[package.scala 93:22:@63592.4]
  wire  RetimeWrapper_159_io_out; // @[package.scala 93:22:@63592.4]
  wire  RetimeWrapper_160_clock; // @[package.scala 93:22:@63613.4]
  wire  RetimeWrapper_160_reset; // @[package.scala 93:22:@63613.4]
  wire  RetimeWrapper_160_io_flow; // @[package.scala 93:22:@63613.4]
  wire  RetimeWrapper_160_io_in; // @[package.scala 93:22:@63613.4]
  wire  RetimeWrapper_160_io_out; // @[package.scala 93:22:@63613.4]
  wire  RetimeWrapper_161_clock; // @[package.scala 93:22:@63622.4]
  wire  RetimeWrapper_161_reset; // @[package.scala 93:22:@63622.4]
  wire  RetimeWrapper_161_io_flow; // @[package.scala 93:22:@63622.4]
  wire [31:0] RetimeWrapper_161_io_in; // @[package.scala 93:22:@63622.4]
  wire [31:0] RetimeWrapper_161_io_out; // @[package.scala 93:22:@63622.4]
  wire  RetimeWrapper_162_clock; // @[package.scala 93:22:@63634.4]
  wire  RetimeWrapper_162_reset; // @[package.scala 93:22:@63634.4]
  wire  RetimeWrapper_162_io_flow; // @[package.scala 93:22:@63634.4]
  wire  RetimeWrapper_162_io_in; // @[package.scala 93:22:@63634.4]
  wire  RetimeWrapper_162_io_out; // @[package.scala 93:22:@63634.4]
  wire  RetimeWrapper_163_clock; // @[package.scala 93:22:@63655.4]
  wire  RetimeWrapper_163_reset; // @[package.scala 93:22:@63655.4]
  wire  RetimeWrapper_163_io_flow; // @[package.scala 93:22:@63655.4]
  wire [31:0] RetimeWrapper_163_io_in; // @[package.scala 93:22:@63655.4]
  wire [31:0] RetimeWrapper_163_io_out; // @[package.scala 93:22:@63655.4]
  wire  RetimeWrapper_164_clock; // @[package.scala 93:22:@63664.4]
  wire  RetimeWrapper_164_reset; // @[package.scala 93:22:@63664.4]
  wire  RetimeWrapper_164_io_flow; // @[package.scala 93:22:@63664.4]
  wire  RetimeWrapper_164_io_in; // @[package.scala 93:22:@63664.4]
  wire  RetimeWrapper_164_io_out; // @[package.scala 93:22:@63664.4]
  wire  RetimeWrapper_165_clock; // @[package.scala 93:22:@63676.4]
  wire  RetimeWrapper_165_reset; // @[package.scala 93:22:@63676.4]
  wire  RetimeWrapper_165_io_flow; // @[package.scala 93:22:@63676.4]
  wire  RetimeWrapper_165_io_in; // @[package.scala 93:22:@63676.4]
  wire  RetimeWrapper_165_io_out; // @[package.scala 93:22:@63676.4]
  wire  x625_1_clock; // @[Math.scala 262:24:@63701.4]
  wire [31:0] x625_1_io_a; // @[Math.scala 262:24:@63701.4]
  wire [31:0] x625_1_io_b; // @[Math.scala 262:24:@63701.4]
  wire  x625_1_io_flow; // @[Math.scala 262:24:@63701.4]
  wire [31:0] x625_1_io_result; // @[Math.scala 262:24:@63701.4]
  wire  x626_1_clock; // @[Math.scala 262:24:@63713.4]
  wire [31:0] x626_1_io_a; // @[Math.scala 262:24:@63713.4]
  wire [31:0] x626_1_io_b; // @[Math.scala 262:24:@63713.4]
  wire  x626_1_io_flow; // @[Math.scala 262:24:@63713.4]
  wire [31:0] x626_1_io_result; // @[Math.scala 262:24:@63713.4]
  wire  x627_1_clock; // @[Math.scala 262:24:@63725.4]
  wire [31:0] x627_1_io_a; // @[Math.scala 262:24:@63725.4]
  wire [31:0] x627_1_io_b; // @[Math.scala 262:24:@63725.4]
  wire  x627_1_io_flow; // @[Math.scala 262:24:@63725.4]
  wire [31:0] x627_1_io_result; // @[Math.scala 262:24:@63725.4]
  wire  x628_1_clock; // @[Math.scala 262:24:@63737.4]
  wire [31:0] x628_1_io_a; // @[Math.scala 262:24:@63737.4]
  wire [31:0] x628_1_io_b; // @[Math.scala 262:24:@63737.4]
  wire  x628_1_io_flow; // @[Math.scala 262:24:@63737.4]
  wire [31:0] x628_1_io_result; // @[Math.scala 262:24:@63737.4]
  wire  x629_x9_1_clock; // @[Math.scala 150:24:@63747.4]
  wire  x629_x9_1_reset; // @[Math.scala 150:24:@63747.4]
  wire [31:0] x629_x9_1_io_a; // @[Math.scala 150:24:@63747.4]
  wire [31:0] x629_x9_1_io_b; // @[Math.scala 150:24:@63747.4]
  wire  x629_x9_1_io_flow; // @[Math.scala 150:24:@63747.4]
  wire [31:0] x629_x9_1_io_result; // @[Math.scala 150:24:@63747.4]
  wire  x630_x10_1_clock; // @[Math.scala 150:24:@63757.4]
  wire  x630_x10_1_reset; // @[Math.scala 150:24:@63757.4]
  wire [31:0] x630_x10_1_io_a; // @[Math.scala 150:24:@63757.4]
  wire [31:0] x630_x10_1_io_b; // @[Math.scala 150:24:@63757.4]
  wire  x630_x10_1_io_flow; // @[Math.scala 150:24:@63757.4]
  wire [31:0] x630_x10_1_io_result; // @[Math.scala 150:24:@63757.4]
  wire  x631_sum_1_clock; // @[Math.scala 150:24:@63767.4]
  wire  x631_sum_1_reset; // @[Math.scala 150:24:@63767.4]
  wire [31:0] x631_sum_1_io_a; // @[Math.scala 150:24:@63767.4]
  wire [31:0] x631_sum_1_io_b; // @[Math.scala 150:24:@63767.4]
  wire  x631_sum_1_io_flow; // @[Math.scala 150:24:@63767.4]
  wire [31:0] x631_sum_1_io_result; // @[Math.scala 150:24:@63767.4]
  wire [31:0] x632_1_io_b; // @[Math.scala 720:24:@63777.4]
  wire [31:0] x632_1_io_result; // @[Math.scala 720:24:@63777.4]
  wire  x633_mul_1_clock; // @[Math.scala 262:24:@63788.4]
  wire [31:0] x633_mul_1_io_a; // @[Math.scala 262:24:@63788.4]
  wire [31:0] x633_mul_1_io_b; // @[Math.scala 262:24:@63788.4]
  wire  x633_mul_1_io_flow; // @[Math.scala 262:24:@63788.4]
  wire [31:0] x633_mul_1_io_result; // @[Math.scala 262:24:@63788.4]
  wire [31:0] x634_1_io_b; // @[Math.scala 720:24:@63798.4]
  wire [31:0] x634_1_io_result; // @[Math.scala 720:24:@63798.4]
  wire  x635_1_clock; // @[Math.scala 262:24:@63809.4]
  wire [31:0] x635_1_io_a; // @[Math.scala 262:24:@63809.4]
  wire [31:0] x635_1_io_b; // @[Math.scala 262:24:@63809.4]
  wire  x635_1_io_flow; // @[Math.scala 262:24:@63809.4]
  wire [31:0] x635_1_io_result; // @[Math.scala 262:24:@63809.4]
  wire  x636_1_clock; // @[Math.scala 262:24:@63821.4]
  wire [31:0] x636_1_io_a; // @[Math.scala 262:24:@63821.4]
  wire [31:0] x636_1_io_b; // @[Math.scala 262:24:@63821.4]
  wire  x636_1_io_flow; // @[Math.scala 262:24:@63821.4]
  wire [31:0] x636_1_io_result; // @[Math.scala 262:24:@63821.4]
  wire  x637_1_clock; // @[Math.scala 262:24:@63833.4]
  wire [31:0] x637_1_io_a; // @[Math.scala 262:24:@63833.4]
  wire [31:0] x637_1_io_b; // @[Math.scala 262:24:@63833.4]
  wire  x637_1_io_flow; // @[Math.scala 262:24:@63833.4]
  wire [31:0] x637_1_io_result; // @[Math.scala 262:24:@63833.4]
  wire  x638_1_clock; // @[Math.scala 262:24:@63845.4]
  wire [31:0] x638_1_io_a; // @[Math.scala 262:24:@63845.4]
  wire [31:0] x638_1_io_b; // @[Math.scala 262:24:@63845.4]
  wire  x638_1_io_flow; // @[Math.scala 262:24:@63845.4]
  wire [31:0] x638_1_io_result; // @[Math.scala 262:24:@63845.4]
  wire  x639_x9_1_clock; // @[Math.scala 150:24:@63855.4]
  wire  x639_x9_1_reset; // @[Math.scala 150:24:@63855.4]
  wire [31:0] x639_x9_1_io_a; // @[Math.scala 150:24:@63855.4]
  wire [31:0] x639_x9_1_io_b; // @[Math.scala 150:24:@63855.4]
  wire  x639_x9_1_io_flow; // @[Math.scala 150:24:@63855.4]
  wire [31:0] x639_x9_1_io_result; // @[Math.scala 150:24:@63855.4]
  wire  x640_x10_1_clock; // @[Math.scala 150:24:@63865.4]
  wire  x640_x10_1_reset; // @[Math.scala 150:24:@63865.4]
  wire [31:0] x640_x10_1_io_a; // @[Math.scala 150:24:@63865.4]
  wire [31:0] x640_x10_1_io_b; // @[Math.scala 150:24:@63865.4]
  wire  x640_x10_1_io_flow; // @[Math.scala 150:24:@63865.4]
  wire [31:0] x640_x10_1_io_result; // @[Math.scala 150:24:@63865.4]
  wire  x641_sum_1_clock; // @[Math.scala 150:24:@63875.4]
  wire  x641_sum_1_reset; // @[Math.scala 150:24:@63875.4]
  wire [31:0] x641_sum_1_io_a; // @[Math.scala 150:24:@63875.4]
  wire [31:0] x641_sum_1_io_b; // @[Math.scala 150:24:@63875.4]
  wire  x641_sum_1_io_flow; // @[Math.scala 150:24:@63875.4]
  wire [31:0] x641_sum_1_io_result; // @[Math.scala 150:24:@63875.4]
  wire [31:0] x642_1_io_b; // @[Math.scala 720:24:@63885.4]
  wire [31:0] x642_1_io_result; // @[Math.scala 720:24:@63885.4]
  wire  x643_mul_1_clock; // @[Math.scala 262:24:@63896.4]
  wire [31:0] x643_mul_1_io_a; // @[Math.scala 262:24:@63896.4]
  wire [31:0] x643_mul_1_io_b; // @[Math.scala 262:24:@63896.4]
  wire  x643_mul_1_io_flow; // @[Math.scala 262:24:@63896.4]
  wire [31:0] x643_mul_1_io_result; // @[Math.scala 262:24:@63896.4]
  wire [31:0] x644_1_io_b; // @[Math.scala 720:24:@63906.4]
  wire [31:0] x644_1_io_result; // @[Math.scala 720:24:@63906.4]
  wire  x645_1_clock; // @[Math.scala 262:24:@63917.4]
  wire [31:0] x645_1_io_a; // @[Math.scala 262:24:@63917.4]
  wire [31:0] x645_1_io_b; // @[Math.scala 262:24:@63917.4]
  wire  x645_1_io_flow; // @[Math.scala 262:24:@63917.4]
  wire [31:0] x645_1_io_result; // @[Math.scala 262:24:@63917.4]
  wire  x646_1_clock; // @[Math.scala 262:24:@63929.4]
  wire [31:0] x646_1_io_a; // @[Math.scala 262:24:@63929.4]
  wire [31:0] x646_1_io_b; // @[Math.scala 262:24:@63929.4]
  wire  x646_1_io_flow; // @[Math.scala 262:24:@63929.4]
  wire [31:0] x646_1_io_result; // @[Math.scala 262:24:@63929.4]
  wire  x647_1_clock; // @[Math.scala 262:24:@63941.4]
  wire [31:0] x647_1_io_a; // @[Math.scala 262:24:@63941.4]
  wire [31:0] x647_1_io_b; // @[Math.scala 262:24:@63941.4]
  wire  x647_1_io_flow; // @[Math.scala 262:24:@63941.4]
  wire [31:0] x647_1_io_result; // @[Math.scala 262:24:@63941.4]
  wire  x648_1_clock; // @[Math.scala 262:24:@63953.4]
  wire [31:0] x648_1_io_a; // @[Math.scala 262:24:@63953.4]
  wire [31:0] x648_1_io_b; // @[Math.scala 262:24:@63953.4]
  wire  x648_1_io_flow; // @[Math.scala 262:24:@63953.4]
  wire [31:0] x648_1_io_result; // @[Math.scala 262:24:@63953.4]
  wire  x649_x9_1_clock; // @[Math.scala 150:24:@63963.4]
  wire  x649_x9_1_reset; // @[Math.scala 150:24:@63963.4]
  wire [31:0] x649_x9_1_io_a; // @[Math.scala 150:24:@63963.4]
  wire [31:0] x649_x9_1_io_b; // @[Math.scala 150:24:@63963.4]
  wire  x649_x9_1_io_flow; // @[Math.scala 150:24:@63963.4]
  wire [31:0] x649_x9_1_io_result; // @[Math.scala 150:24:@63963.4]
  wire  x650_x10_1_clock; // @[Math.scala 150:24:@63975.4]
  wire  x650_x10_1_reset; // @[Math.scala 150:24:@63975.4]
  wire [31:0] x650_x10_1_io_a; // @[Math.scala 150:24:@63975.4]
  wire [31:0] x650_x10_1_io_b; // @[Math.scala 150:24:@63975.4]
  wire  x650_x10_1_io_flow; // @[Math.scala 150:24:@63975.4]
  wire [31:0] x650_x10_1_io_result; // @[Math.scala 150:24:@63975.4]
  wire  x651_sum_1_clock; // @[Math.scala 150:24:@63985.4]
  wire  x651_sum_1_reset; // @[Math.scala 150:24:@63985.4]
  wire [31:0] x651_sum_1_io_a; // @[Math.scala 150:24:@63985.4]
  wire [31:0] x651_sum_1_io_b; // @[Math.scala 150:24:@63985.4]
  wire  x651_sum_1_io_flow; // @[Math.scala 150:24:@63985.4]
  wire [31:0] x651_sum_1_io_result; // @[Math.scala 150:24:@63985.4]
  wire [31:0] x652_1_io_b; // @[Math.scala 720:24:@63995.4]
  wire [31:0] x652_1_io_result; // @[Math.scala 720:24:@63995.4]
  wire  x653_mul_1_clock; // @[Math.scala 262:24:@64006.4]
  wire [31:0] x653_mul_1_io_a; // @[Math.scala 262:24:@64006.4]
  wire [31:0] x653_mul_1_io_b; // @[Math.scala 262:24:@64006.4]
  wire  x653_mul_1_io_flow; // @[Math.scala 262:24:@64006.4]
  wire [31:0] x653_mul_1_io_result; // @[Math.scala 262:24:@64006.4]
  wire [31:0] x654_1_io_b; // @[Math.scala 720:24:@64016.4]
  wire [31:0] x654_1_io_result; // @[Math.scala 720:24:@64016.4]
  wire  x655_1_clock; // @[Math.scala 262:24:@64027.4]
  wire [31:0] x655_1_io_a; // @[Math.scala 262:24:@64027.4]
  wire [31:0] x655_1_io_b; // @[Math.scala 262:24:@64027.4]
  wire  x655_1_io_flow; // @[Math.scala 262:24:@64027.4]
  wire [31:0] x655_1_io_result; // @[Math.scala 262:24:@64027.4]
  wire  x656_1_clock; // @[Math.scala 262:24:@64039.4]
  wire [31:0] x656_1_io_a; // @[Math.scala 262:24:@64039.4]
  wire [31:0] x656_1_io_b; // @[Math.scala 262:24:@64039.4]
  wire  x656_1_io_flow; // @[Math.scala 262:24:@64039.4]
  wire [31:0] x656_1_io_result; // @[Math.scala 262:24:@64039.4]
  wire  x657_1_clock; // @[Math.scala 262:24:@64051.4]
  wire [31:0] x657_1_io_a; // @[Math.scala 262:24:@64051.4]
  wire [31:0] x657_1_io_b; // @[Math.scala 262:24:@64051.4]
  wire  x657_1_io_flow; // @[Math.scala 262:24:@64051.4]
  wire [31:0] x657_1_io_result; // @[Math.scala 262:24:@64051.4]
  wire  x658_1_clock; // @[Math.scala 262:24:@64063.4]
  wire [31:0] x658_1_io_a; // @[Math.scala 262:24:@64063.4]
  wire [31:0] x658_1_io_b; // @[Math.scala 262:24:@64063.4]
  wire  x658_1_io_flow; // @[Math.scala 262:24:@64063.4]
  wire [31:0] x658_1_io_result; // @[Math.scala 262:24:@64063.4]
  wire  x659_x9_1_clock; // @[Math.scala 150:24:@64073.4]
  wire  x659_x9_1_reset; // @[Math.scala 150:24:@64073.4]
  wire [31:0] x659_x9_1_io_a; // @[Math.scala 150:24:@64073.4]
  wire [31:0] x659_x9_1_io_b; // @[Math.scala 150:24:@64073.4]
  wire  x659_x9_1_io_flow; // @[Math.scala 150:24:@64073.4]
  wire [31:0] x659_x9_1_io_result; // @[Math.scala 150:24:@64073.4]
  wire  x660_x10_1_clock; // @[Math.scala 150:24:@64083.4]
  wire  x660_x10_1_reset; // @[Math.scala 150:24:@64083.4]
  wire [31:0] x660_x10_1_io_a; // @[Math.scala 150:24:@64083.4]
  wire [31:0] x660_x10_1_io_b; // @[Math.scala 150:24:@64083.4]
  wire  x660_x10_1_io_flow; // @[Math.scala 150:24:@64083.4]
  wire [31:0] x660_x10_1_io_result; // @[Math.scala 150:24:@64083.4]
  wire  x661_sum_1_clock; // @[Math.scala 150:24:@64093.4]
  wire  x661_sum_1_reset; // @[Math.scala 150:24:@64093.4]
  wire [31:0] x661_sum_1_io_a; // @[Math.scala 150:24:@64093.4]
  wire [31:0] x661_sum_1_io_b; // @[Math.scala 150:24:@64093.4]
  wire  x661_sum_1_io_flow; // @[Math.scala 150:24:@64093.4]
  wire [31:0] x661_sum_1_io_result; // @[Math.scala 150:24:@64093.4]
  wire [31:0] x662_1_io_b; // @[Math.scala 720:24:@64103.4]
  wire [31:0] x662_1_io_result; // @[Math.scala 720:24:@64103.4]
  wire  x663_mul_1_clock; // @[Math.scala 262:24:@64114.4]
  wire [31:0] x663_mul_1_io_a; // @[Math.scala 262:24:@64114.4]
  wire [31:0] x663_mul_1_io_b; // @[Math.scala 262:24:@64114.4]
  wire  x663_mul_1_io_flow; // @[Math.scala 262:24:@64114.4]
  wire [31:0] x663_mul_1_io_result; // @[Math.scala 262:24:@64114.4]
  wire [31:0] x664_1_io_b; // @[Math.scala 720:24:@64124.4]
  wire [31:0] x664_1_io_result; // @[Math.scala 720:24:@64124.4]
  wire  RetimeWrapper_166_clock; // @[package.scala 93:22:@64143.4]
  wire  RetimeWrapper_166_reset; // @[package.scala 93:22:@64143.4]
  wire  RetimeWrapper_166_io_flow; // @[package.scala 93:22:@64143.4]
  wire [127:0] RetimeWrapper_166_io_in; // @[package.scala 93:22:@64143.4]
  wire [127:0] RetimeWrapper_166_io_out; // @[package.scala 93:22:@64143.4]
  wire  RetimeWrapper_167_clock; // @[package.scala 93:22:@64152.4]
  wire  RetimeWrapper_167_reset; // @[package.scala 93:22:@64152.4]
  wire  RetimeWrapper_167_io_flow; // @[package.scala 93:22:@64152.4]
  wire  RetimeWrapper_167_io_in; // @[package.scala 93:22:@64152.4]
  wire  RetimeWrapper_167_io_out; // @[package.scala 93:22:@64152.4]
  wire  RetimeWrapper_168_clock; // @[package.scala 93:22:@64161.4]
  wire  RetimeWrapper_168_reset; // @[package.scala 93:22:@64161.4]
  wire  RetimeWrapper_168_io_flow; // @[package.scala 93:22:@64161.4]
  wire  RetimeWrapper_168_io_in; // @[package.scala 93:22:@64161.4]
  wire  RetimeWrapper_168_io_out; // @[package.scala 93:22:@64161.4]
  wire  RetimeWrapper_169_clock; // @[package.scala 93:22:@64170.4]
  wire  RetimeWrapper_169_reset; // @[package.scala 93:22:@64170.4]
  wire  RetimeWrapper_169_io_flow; // @[package.scala 93:22:@64170.4]
  wire  RetimeWrapper_169_io_in; // @[package.scala 93:22:@64170.4]
  wire  RetimeWrapper_169_io_out; // @[package.scala 93:22:@64170.4]
  wire  b379; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 62:18:@59847.4]
  wire  b380; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 63:18:@59848.4]
  wire  _T_205; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 67:30:@59850.4]
  wire  _T_206; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 67:37:@59851.4]
  wire  _T_210; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 69:76:@59856.4]
  wire  _T_211; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 69:62:@59857.4]
  wire  _T_213; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 69:101:@59858.4]
  wire [127:0] x745_x381_D1_0_number; // @[package.scala 96:25:@59867.4 package.scala 96:25:@59868.4]
  wire [31:0] b377_number; // @[Math.scala 723:22:@59832.4 Math.scala 724:14:@59833.4]
  wire [31:0] _T_248; // @[Math.scala 406:49:@60129.4]
  wire [31:0] _T_250; // @[Math.scala 406:56:@60131.4]
  wire [31:0] _T_251; // @[Math.scala 406:56:@60132.4]
  wire [31:0] x725_number; // @[implicits.scala 133:21:@60133.4]
  wire [31:0] _T_261; // @[Math.scala 406:49:@60142.4]
  wire [31:0] _T_263; // @[Math.scala 406:56:@60144.4]
  wire [31:0] _T_264; // @[Math.scala 406:56:@60145.4]
  wire  _T_275; // @[FixedPoint.scala 50:25:@60163.4]
  wire [1:0] _T_279; // @[Bitwise.scala 72:12:@60165.4]
  wire [29:0] _T_280; // @[FixedPoint.scala 18:52:@60166.4]
  wire  _T_286; // @[Math.scala 451:55:@60168.4]
  wire [1:0] _T_287; // @[FixedPoint.scala 18:52:@60169.4]
  wire  _T_293; // @[Math.scala 451:110:@60171.4]
  wire  _T_294; // @[Math.scala 451:94:@60172.4]
  wire [31:0] _T_296; // @[Cat.scala 30:58:@60174.4]
  wire [31:0] x390_1_number; // @[Math.scala 454:20:@60175.4]
  wire [39:0] _GEN_0; // @[Math.scala 461:32:@60180.4]
  wire [39:0] _T_301; // @[Math.scala 461:32:@60180.4]
  wire [37:0] _GEN_1; // @[Math.scala 461:32:@60185.4]
  wire [37:0] _T_304; // @[Math.scala 461:32:@60185.4]
  wire  _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:101:@60283.4]
  wire  _T_344; // @[package.scala 96:25:@60291.4 package.scala 96:25:@60292.4]
  wire  _T_346; // @[implicits.scala 55:10:@60293.4]
  wire  _T_347; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:118:@60294.4]
  wire  _T_349; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:207:@60296.4]
  wire  _T_350; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:226:@60297.4]
  wire  x747_b379_D24; // @[package.scala 96:25:@60235.4 package.scala 96:25:@60236.4]
  wire  _T_351; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:252:@60298.4]
  wire  x749_b380_D24; // @[package.scala 96:25:@60253.4 package.scala 96:25:@60254.4]
  wire  _T_395; // @[package.scala 96:25:@60398.4 package.scala 96:25:@60399.4]
  wire  _T_397; // @[implicits.scala 55:10:@60400.4]
  wire  _T_398; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 141:118:@60401.4]
  wire  _T_400; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 141:207:@60403.4]
  wire  _T_401; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 141:226:@60404.4]
  wire  _T_402; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 141:252:@60405.4]
  wire  _T_443; // @[package.scala 96:25:@60496.4 package.scala 96:25:@60497.4]
  wire  _T_445; // @[implicits.scala 55:10:@60498.4]
  wire  _T_446; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 162:118:@60499.4]
  wire  _T_448; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 162:207:@60501.4]
  wire  _T_449; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 162:226:@60502.4]
  wire  _T_450; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 162:252:@60503.4]
  wire  _T_491; // @[package.scala 96:25:@60594.4 package.scala 96:25:@60595.4]
  wire  _T_493; // @[implicits.scala 55:10:@60596.4]
  wire  _T_494; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 189:166:@60597.4]
  wire  _T_496; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 189:255:@60599.4]
  wire  _T_497; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 189:274:@60600.4]
  wire  _T_498; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 189:300:@60601.4]
  wire [31:0] x763_b377_D26_number; // @[package.scala 96:25:@60615.4 package.scala 96:25:@60616.4]
  wire [31:0] _T_510; // @[Math.scala 476:37:@60623.4]
  wire [31:0] x764_x407_rdcol_D26_number; // @[package.scala 96:25:@60640.4 package.scala 96:25:@60641.4]
  wire [31:0] _T_523; // @[Math.scala 476:37:@60646.4]
  wire  x765_x414_D1; // @[package.scala 96:25:@60663.4 package.scala 96:25:@60664.4]
  wire  x415; // @[package.scala 96:25:@60654.4 package.scala 96:25:@60655.4]
  wire  x416; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 204:24:@60667.4]
  wire  _T_564; // @[package.scala 96:25:@60735.4 package.scala 96:25:@60736.4]
  wire  _T_566; // @[implicits.scala 55:10:@60737.4]
  wire  _T_567; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 223:194:@60738.4]
  wire  x767_x417_D20; // @[package.scala 96:25:@60687.4 package.scala 96:25:@60688.4]
  wire  _T_568; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 223:283:@60739.4]
  wire  x766_b379_D48; // @[package.scala 96:25:@60678.4 package.scala 96:25:@60679.4]
  wire  _T_569; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 223:291:@60740.4]
  wire  x769_b380_D48; // @[package.scala 96:25:@60705.4 package.scala 96:25:@60706.4]
  wire [31:0] x772_x401_rdcol_D26_number; // @[package.scala 96:25:@60756.4 package.scala 96:25:@60757.4]
  wire [31:0] _T_580; // @[Math.scala 476:37:@60762.4]
  wire  x420; // @[package.scala 96:25:@60770.4 package.scala 96:25:@60771.4]
  wire  x421; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 231:24:@60774.4]
  wire  _T_609; // @[package.scala 96:25:@60815.4 package.scala 96:25:@60816.4]
  wire  _T_611; // @[implicits.scala 55:10:@60817.4]
  wire  _T_612; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 244:194:@60818.4]
  wire  x775_x422_D20; // @[package.scala 96:25:@60803.4 package.scala 96:25:@60804.4]
  wire  _T_613; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 244:283:@60819.4]
  wire  _T_614; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 244:291:@60820.4]
  wire [31:0] x776_x395_rdcol_D26_number; // @[package.scala 96:25:@60836.4 package.scala 96:25:@60837.4]
  wire [31:0] _T_625; // @[Math.scala 476:37:@60842.4]
  wire  x425; // @[package.scala 96:25:@60850.4 package.scala 96:25:@60851.4]
  wire  x426; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 252:24:@60854.4]
  wire  _T_654; // @[package.scala 96:25:@60895.4 package.scala 96:25:@60896.4]
  wire  _T_656; // @[implicits.scala 55:10:@60897.4]
  wire  _T_657; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 265:194:@60898.4]
  wire  x779_x427_D20; // @[package.scala 96:25:@60883.4 package.scala 96:25:@60884.4]
  wire  _T_658; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 265:283:@60899.4]
  wire  _T_659; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 265:291:@60900.4]
  wire [31:0] x780_b378_D26_number; // @[package.scala 96:25:@60916.4 package.scala 96:25:@60917.4]
  wire [31:0] _T_670; // @[Math.scala 476:37:@60922.4]
  wire  x414; // @[package.scala 96:25:@60631.4 package.scala 96:25:@60632.4]
  wire  x430; // @[package.scala 96:25:@60930.4 package.scala 96:25:@60931.4]
  wire  x431; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 273:24:@60934.4]
  wire  _T_699; // @[package.scala 96:25:@60975.4 package.scala 96:25:@60976.4]
  wire  _T_701; // @[implicits.scala 55:10:@60977.4]
  wire  _T_702; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 286:194:@60978.4]
  wire  x783_x432_D21; // @[package.scala 96:25:@60963.4 package.scala 96:25:@60964.4]
  wire  _T_703; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 286:283:@60979.4]
  wire  _T_704; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 286:291:@60980.4]
  wire [31:0] x435_rdcol_number; // @[Math.scala 154:22:@60999.4 Math.scala 155:14:@61000.4]
  wire [31:0] _T_719; // @[Math.scala 476:37:@61005.4]
  wire  x436; // @[package.scala 96:25:@61013.4 package.scala 96:25:@61014.4]
  wire  x437; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 294:24:@61017.4]
  wire  _T_767; // @[package.scala 96:25:@61094.4 package.scala 96:25:@61095.4]
  wire  _T_769; // @[implicits.scala 55:10:@61096.4]
  wire  _T_770; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 321:194:@61097.4]
  wire  x786_x438_D20; // @[package.scala 96:25:@61082.4 package.scala 96:25:@61083.4]
  wire  _T_771; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 321:283:@61098.4]
  wire  _T_772; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 321:291:@61099.4]
  wire [31:0] x444_rdcol_number; // @[Math.scala 154:22:@61118.4 Math.scala 155:14:@61119.4]
  wire [31:0] _T_787; // @[Math.scala 476:37:@61124.4]
  wire  x445; // @[package.scala 96:25:@61132.4 package.scala 96:25:@61133.4]
  wire  x446; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 329:59:@61136.4]
  wire  _T_830; // @[package.scala 96:25:@61202.4 package.scala 96:25:@61203.4]
  wire  _T_832; // @[implicits.scala 55:10:@61204.4]
  wire  _T_833; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 346:194:@61205.4]
  wire  x788_x447_D20; // @[package.scala 96:25:@61190.4 package.scala 96:25:@61191.4]
  wire  _T_834; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 346:283:@61206.4]
  wire  _T_835; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 346:291:@61207.4]
  wire [31:0] x453_rdrow_number; // @[Math.scala 195:22:@61226.4 Math.scala 196:14:@61227.4]
  wire [31:0] _T_852; // @[Math.scala 406:49:@61233.4]
  wire [31:0] _T_854; // @[Math.scala 406:56:@61235.4]
  wire [31:0] _T_855; // @[Math.scala 406:56:@61236.4]
  wire [31:0] x730_number; // @[implicits.scala 133:21:@61237.4]
  wire  x455; // @[package.scala 96:25:@61251.4 package.scala 96:25:@61252.4]
  wire  x456; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 356:24:@61255.4]
  wire [31:0] _T_878; // @[Math.scala 406:49:@61264.4]
  wire [31:0] _T_880; // @[Math.scala 406:56:@61266.4]
  wire [31:0] _T_881; // @[Math.scala 406:56:@61267.4]
  wire [31:0] _T_885; // @[package.scala 96:25:@61275.4]
  wire  _T_889; // @[FixedPoint.scala 50:25:@61282.4]
  wire [1:0] _T_893; // @[Bitwise.scala 72:12:@61284.4]
  wire [29:0] _T_894; // @[FixedPoint.scala 18:52:@61285.4]
  wire  _T_900; // @[Math.scala 451:55:@61287.4]
  wire [1:0] _T_901; // @[FixedPoint.scala 18:52:@61288.4]
  wire  _T_907; // @[Math.scala 451:110:@61290.4]
  wire  _T_908; // @[Math.scala 451:94:@61291.4]
  wire [31:0] _T_912; // @[package.scala 96:25:@61299.4 package.scala 96:25:@61300.4]
  wire [31:0] x459_1_number; // @[Math.scala 454:20:@61301.4]
  wire [39:0] _GEN_2; // @[Math.scala 461:32:@61306.4]
  wire [39:0] _T_917; // @[Math.scala 461:32:@61306.4]
  wire [37:0] _GEN_3; // @[Math.scala 461:32:@61311.4]
  wire [37:0] _T_920; // @[Math.scala 461:32:@61311.4]
  wire  _T_950; // @[package.scala 96:25:@61379.4 package.scala 96:25:@61380.4]
  wire  _T_952; // @[implicits.scala 55:10:@61381.4]
  wire  _T_953; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 383:194:@61382.4]
  wire  x791_x457_D20; // @[package.scala 96:25:@61358.4 package.scala 96:25:@61359.4]
  wire  _T_954; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 383:283:@61383.4]
  wire  _T_955; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 383:291:@61384.4]
  wire  x464; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 387:24:@61395.4]
  wire  _T_982; // @[package.scala 96:25:@61437.4 package.scala 96:25:@61438.4]
  wire  _T_984; // @[implicits.scala 55:10:@61439.4]
  wire  _T_985; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 400:194:@61440.4]
  wire  x794_x465_D20; // @[package.scala 96:25:@61425.4 package.scala 96:25:@61426.4]
  wire  _T_986; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 400:283:@61441.4]
  wire  _T_987; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 400:291:@61442.4]
  wire  x469; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 404:24:@61453.4]
  wire  _T_1014; // @[package.scala 96:25:@61495.4 package.scala 96:25:@61496.4]
  wire  _T_1016; // @[implicits.scala 55:10:@61497.4]
  wire  _T_1017; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 423:194:@61498.4]
  wire  x796_x470_D20; // @[package.scala 96:25:@61483.4 package.scala 96:25:@61484.4]
  wire  _T_1018; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 423:283:@61499.4]
  wire  _T_1019; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 423:326:@61500.4]
  wire  x797_x430_D1; // @[package.scala 96:25:@61516.4 package.scala 96:25:@61517.4]
  wire  x474; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 429:59:@61520.4]
  wire  _T_1057; // @[package.scala 96:25:@61582.4 package.scala 96:25:@61583.4]
  wire  _T_1059; // @[implicits.scala 55:10:@61584.4]
  wire  _T_1060; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 448:194:@61585.4]
  wire  x800_x475_D20; // @[package.scala 96:25:@61561.4 package.scala 96:25:@61562.4]
  wire  _T_1061; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 448:283:@61586.4]
  wire  _T_1062; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 448:291:@61587.4]
  wire  x479; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 452:59:@61598.4]
  wire  _T_1086; // @[package.scala 96:25:@61631.4 package.scala 96:25:@61632.4]
  wire  _T_1088; // @[implicits.scala 55:10:@61633.4]
  wire  _T_1089; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 463:194:@61634.4]
  wire  x802_x480_D20; // @[package.scala 96:25:@61619.4 package.scala 96:25:@61620.4]
  wire  _T_1090; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 463:283:@61635.4]
  wire  _T_1091; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 463:291:@61636.4]
  wire  x484; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 467:59:@61647.4]
  wire  _T_1115; // @[package.scala 96:25:@61680.4 package.scala 96:25:@61681.4]
  wire  _T_1117; // @[implicits.scala 55:10:@61682.4]
  wire  _T_1118; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 478:194:@61683.4]
  wire  x803_x485_D20; // @[package.scala 96:25:@61668.4 package.scala 96:25:@61669.4]
  wire  _T_1119; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 478:283:@61684.4]
  wire  _T_1120; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 478:291:@61685.4]
  wire [31:0] x489_rdrow_number; // @[Math.scala 195:22:@61704.4 Math.scala 196:14:@61705.4]
  wire [31:0] _T_1137; // @[Math.scala 406:49:@61711.4]
  wire [31:0] _T_1139; // @[Math.scala 406:56:@61713.4]
  wire [31:0] _T_1140; // @[Math.scala 406:56:@61714.4]
  wire [31:0] x735_number; // @[implicits.scala 133:21:@61715.4]
  wire  x491; // @[package.scala 96:25:@61729.4 package.scala 96:25:@61730.4]
  wire  x492; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 488:24:@61733.4]
  wire [31:0] _T_1163; // @[Math.scala 406:49:@61742.4]
  wire [31:0] _T_1165; // @[Math.scala 406:56:@61744.4]
  wire [31:0] _T_1166; // @[Math.scala 406:56:@61745.4]
  wire [31:0] _T_1170; // @[package.scala 96:25:@61753.4]
  wire  _T_1174; // @[FixedPoint.scala 50:25:@61760.4]
  wire [1:0] _T_1178; // @[Bitwise.scala 72:12:@61762.4]
  wire [29:0] _T_1179; // @[FixedPoint.scala 18:52:@61763.4]
  wire  _T_1185; // @[Math.scala 451:55:@61765.4]
  wire [1:0] _T_1186; // @[FixedPoint.scala 18:52:@61766.4]
  wire  _T_1192; // @[Math.scala 451:110:@61768.4]
  wire  _T_1193; // @[Math.scala 451:94:@61769.4]
  wire [31:0] _T_1197; // @[package.scala 96:25:@61777.4 package.scala 96:25:@61778.4]
  wire [31:0] x495_1_number; // @[Math.scala 454:20:@61779.4]
  wire [39:0] _GEN_4; // @[Math.scala 461:32:@61784.4]
  wire [39:0] _T_1202; // @[Math.scala 461:32:@61784.4]
  wire [37:0] _GEN_5; // @[Math.scala 461:32:@61789.4]
  wire [37:0] _T_1205; // @[Math.scala 461:32:@61789.4]
  wire  _T_1232; // @[package.scala 96:25:@61848.4 package.scala 96:25:@61849.4]
  wire  _T_1234; // @[implicits.scala 55:10:@61850.4]
  wire  _T_1235; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 513:194:@61851.4]
  wire  x805_x493_D20; // @[package.scala 96:25:@61827.4 package.scala 96:25:@61828.4]
  wire  _T_1236; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 513:283:@61852.4]
  wire  _T_1237; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 513:291:@61853.4]
  wire  x500; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 517:24:@61864.4]
  wire  _T_1261; // @[package.scala 96:25:@61897.4 package.scala 96:25:@61898.4]
  wire  _T_1263; // @[implicits.scala 55:10:@61899.4]
  wire  _T_1264; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 528:194:@61900.4]
  wire  x807_x501_D20; // @[package.scala 96:25:@61885.4 package.scala 96:25:@61886.4]
  wire  _T_1265; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 528:283:@61901.4]
  wire  _T_1266; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 528:291:@61902.4]
  wire  x505; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 532:24:@61913.4]
  wire  _T_1290; // @[package.scala 96:25:@61946.4 package.scala 96:25:@61947.4]
  wire  _T_1292; // @[implicits.scala 55:10:@61948.4]
  wire  _T_1293; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 549:194:@61949.4]
  wire  x808_x506_D20; // @[package.scala 96:25:@61934.4 package.scala 96:25:@61935.4]
  wire  _T_1294; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 549:283:@61950.4]
  wire  _T_1295; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 549:291:@61951.4]
  wire  x510; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 553:59:@61962.4]
  wire  _T_1327; // @[package.scala 96:25:@62015.4 package.scala 96:25:@62016.4]
  wire  _T_1329; // @[implicits.scala 55:10:@62017.4]
  wire  _T_1330; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 570:194:@62018.4]
  wire  x810_x511_D20; // @[package.scala 96:25:@61994.4 package.scala 96:25:@61995.4]
  wire  _T_1331; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 570:283:@62019.4]
  wire  _T_1332; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 570:291:@62020.4]
  wire  x515; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 574:59:@62031.4]
  wire  _T_1356; // @[package.scala 96:25:@62064.4 package.scala 96:25:@62065.4]
  wire  _T_1358; // @[implicits.scala 55:10:@62066.4]
  wire  _T_1359; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 585:194:@62067.4]
  wire  x812_x516_D20; // @[package.scala 96:25:@62052.4 package.scala 96:25:@62053.4]
  wire  _T_1360; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 585:283:@62068.4]
  wire  _T_1361; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 585:291:@62069.4]
  wire  x520; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 589:59:@62080.4]
  wire  _T_1385; // @[package.scala 96:25:@62113.4 package.scala 96:25:@62114.4]
  wire  _T_1387; // @[implicits.scala 55:10:@62115.4]
  wire  _T_1388; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 600:194:@62116.4]
  wire  x813_x521_D20; // @[package.scala 96:25:@62101.4 package.scala 96:25:@62102.4]
  wire  _T_1389; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 600:283:@62117.4]
  wire  _T_1390; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 600:291:@62118.4]
  wire  _T_1790; // @[package.scala 96:25:@63030.4 package.scala 96:25:@63031.4]
  wire  _T_1792; // @[implicits.scala 55:10:@63032.4]
  wire  _T_1793; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 792:167:@63033.4]
  wire  _T_1795; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 792:256:@63035.4]
  wire  _T_1796; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 792:275:@63036.4]
  wire  x818_b379_D67; // @[package.scala 96:25:@62974.4 package.scala 96:25:@62975.4]
  wire  _T_1797; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 792:301:@63037.4]
  wire  x820_b380_D67; // @[package.scala 96:25:@62992.4 package.scala 96:25:@62993.4]
  wire  _T_1813; // @[package.scala 96:25:@63080.4 package.scala 96:25:@63081.4]
  wire  _T_1815; // @[implicits.scala 55:10:@63082.4]
  wire  _T_1816; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 803:167:@63083.4]
  wire  _T_1818; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 803:256:@63085.4]
  wire  _T_1819; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 803:275:@63086.4]
  wire  _T_1820; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 803:301:@63087.4]
  wire  _T_1836; // @[package.scala 96:25:@63130.4 package.scala 96:25:@63131.4]
  wire  _T_1838; // @[implicits.scala 55:10:@63132.4]
  wire  _T_1839; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 814:167:@63133.4]
  wire  _T_1841; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 814:256:@63135.4]
  wire  _T_1842; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 814:275:@63136.4]
  wire  _T_1843; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 814:301:@63137.4]
  wire  _T_1859; // @[package.scala 96:25:@63180.4 package.scala 96:25:@63181.4]
  wire  _T_1861; // @[implicits.scala 55:10:@63182.4]
  wire  _T_1862; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 825:167:@63183.4]
  wire  _T_1864; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 825:256:@63185.4]
  wire  _T_1865; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 825:275:@63186.4]
  wire  _T_1866; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 825:301:@63187.4]
  wire  _T_1897; // @[package.scala 96:25:@63258.4 package.scala 96:25:@63259.4]
  wire  _T_1899; // @[implicits.scala 55:10:@63260.4]
  wire  _T_1900; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 843:195:@63261.4]
  wire  x834_x417_D40; // @[package.scala 96:25:@63210.4 package.scala 96:25:@63211.4]
  wire  _T_1901; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 843:284:@63262.4]
  wire  x833_b379_D68; // @[package.scala 96:25:@63201.4 package.scala 96:25:@63202.4]
  wire  _T_1902; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 843:292:@63263.4]
  wire  x836_b380_D68; // @[package.scala 96:25:@63228.4 package.scala 96:25:@63229.4]
  wire  _T_1925; // @[package.scala 96:25:@63309.4 package.scala 96:25:@63310.4]
  wire  _T_1927; // @[implicits.scala 55:10:@63311.4]
  wire  _T_1928; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 856:195:@63312.4]
  wire  x841_x422_D40; // @[package.scala 96:25:@63297.4 package.scala 96:25:@63298.4]
  wire  _T_1929; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 856:284:@63313.4]
  wire  _T_1930; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 856:292:@63314.4]
  wire  _T_1953; // @[package.scala 96:25:@63360.4 package.scala 96:25:@63361.4]
  wire  _T_1955; // @[implicits.scala 55:10:@63362.4]
  wire  _T_1956; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 869:195:@63363.4]
  wire  x844_x427_D40; // @[package.scala 96:25:@63348.4 package.scala 96:25:@63349.4]
  wire  _T_1957; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 869:284:@63364.4]
  wire  _T_1958; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 869:292:@63365.4]
  wire  _T_1981; // @[package.scala 96:25:@63411.4 package.scala 96:25:@63412.4]
  wire  _T_1983; // @[implicits.scala 55:10:@63413.4]
  wire  _T_1984; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 882:195:@63414.4]
  wire  x847_x432_D41; // @[package.scala 96:25:@63399.4 package.scala 96:25:@63400.4]
  wire  _T_1985; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 882:284:@63415.4]
  wire  _T_1986; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 882:292:@63416.4]
  wire  _T_2009; // @[package.scala 96:25:@63462.4 package.scala 96:25:@63463.4]
  wire  _T_2011; // @[implicits.scala 55:10:@63464.4]
  wire  _T_2012; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 901:195:@63465.4]
  wire  x849_x438_D40; // @[package.scala 96:25:@63441.4 package.scala 96:25:@63442.4]
  wire  _T_2013; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 901:284:@63466.4]
  wire  _T_2014; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 901:327:@63467.4]
  wire  _T_2037; // @[package.scala 96:25:@63513.4 package.scala 96:25:@63514.4]
  wire  _T_2039; // @[implicits.scala 55:10:@63515.4]
  wire  _T_2040; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 914:195:@63516.4]
  wire  x852_x457_D40; // @[package.scala 96:25:@63492.4 package.scala 96:25:@63493.4]
  wire  _T_2041; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 914:284:@63517.4]
  wire  _T_2042; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 914:292:@63518.4]
  wire  _T_2062; // @[package.scala 96:25:@63555.4 package.scala 96:25:@63556.4]
  wire  _T_2064; // @[implicits.scala 55:10:@63557.4]
  wire  _T_2065; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 925:195:@63558.4]
  wire  x855_x465_D40; // @[package.scala 96:25:@63543.4 package.scala 96:25:@63544.4]
  wire  _T_2066; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 925:284:@63559.4]
  wire  _T_2067; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 925:292:@63560.4]
  wire  _T_2087; // @[package.scala 96:25:@63597.4 package.scala 96:25:@63598.4]
  wire  _T_2089; // @[implicits.scala 55:10:@63599.4]
  wire  _T_2090; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 936:195:@63600.4]
  wire  x857_x470_D40; // @[package.scala 96:25:@63585.4 package.scala 96:25:@63586.4]
  wire  _T_2091; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 936:284:@63601.4]
  wire  _T_2092; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 936:292:@63602.4]
  wire  _T_2112; // @[package.scala 96:25:@63639.4 package.scala 96:25:@63640.4]
  wire  _T_2114; // @[implicits.scala 55:10:@63641.4]
  wire  _T_2115; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 947:195:@63642.4]
  wire  x858_x475_D40; // @[package.scala 96:25:@63618.4 package.scala 96:25:@63619.4]
  wire  _T_2116; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 947:284:@63643.4]
  wire  _T_2117; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 947:292:@63644.4]
  wire  _T_2137; // @[package.scala 96:25:@63681.4 package.scala 96:25:@63682.4]
  wire  _T_2139; // @[implicits.scala 55:10:@63683.4]
  wire  _T_2140; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 958:195:@63684.4]
  wire  x861_x480_D40; // @[package.scala 96:25:@63669.4 package.scala 96:25:@63670.4]
  wire  _T_2141; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 958:284:@63685.4]
  wire  _T_2142; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 958:292:@63686.4]
  wire [31:0] x654_number; // @[Math.scala 723:22:@64021.4 Math.scala 724:14:@64022.4]
  wire [31:0] x664_number; // @[Math.scala 723:22:@64129.4 Math.scala 724:14:@64130.4]
  wire [63:0] _T_2360; // @[Cat.scala 30:58:@64138.4]
  wire [31:0] x634_number; // @[Math.scala 723:22:@63803.4 Math.scala 724:14:@63804.4]
  wire [31:0] x644_number; // @[Math.scala 723:22:@63911.4 Math.scala 724:14:@63912.4]
  wire [63:0] _T_2361; // @[Cat.scala 30:58:@64139.4]
  wire  _T_2374; // @[package.scala 96:25:@64175.4 package.scala 96:25:@64176.4]
  wire  _T_2376; // @[implicits.scala 55:10:@64177.4]
  wire  x863_b379_D87; // @[package.scala 96:25:@64166.4 package.scala 96:25:@64167.4]
  wire  _T_2377; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1060:117:@64178.4]
  wire  x862_b380_D87; // @[package.scala 96:25:@64157.4 package.scala 96:25:@64158.4]
  wire  _T_2378; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1060:123:@64179.4]
  wire [31:0] x748_x389_D8_number; // @[package.scala 96:25:@60244.4 package.scala 96:25:@60245.4]
  wire [31:0] x750_x393_sum_D3_number; // @[package.scala 96:25:@60262.4 package.scala 96:25:@60263.4]
  wire [31:0] x752_x726_D24_number; // @[package.scala 96:25:@60280.4 package.scala 96:25:@60281.4]
  wire [31:0] x754_x397_D7_number; // @[package.scala 96:25:@60369.4 package.scala 96:25:@60370.4]
  wire [31:0] x756_x399_sum_D2_number; // @[package.scala 96:25:@60387.4 package.scala 96:25:@60388.4]
  wire [31:0] x757_x403_D7_number; // @[package.scala 96:25:@60467.4 package.scala 96:25:@60468.4]
  wire [31:0] x759_x405_sum_D2_number; // @[package.scala 96:25:@60485.4 package.scala 96:25:@60486.4]
  wire [31:0] x761_x411_sum_D2_number; // @[package.scala 96:25:@60574.4 package.scala 96:25:@60575.4]
  wire [31:0] x762_x409_D7_number; // @[package.scala 96:25:@60583.4 package.scala 96:25:@60584.4]
  wire [31:0] x768_x411_sum_D26_number; // @[package.scala 96:25:@60696.4 package.scala 96:25:@60697.4]
  wire [31:0] x770_x726_D48_number; // @[package.scala 96:25:@60714.4 package.scala 96:25:@60715.4]
  wire [31:0] x771_x409_D31_number; // @[package.scala 96:25:@60723.4 package.scala 96:25:@60724.4]
  wire [31:0] x773_x403_D31_number; // @[package.scala 96:25:@60785.4 package.scala 96:25:@60786.4]
  wire [31:0] x774_x405_sum_D26_number; // @[package.scala 96:25:@60794.4 package.scala 96:25:@60795.4]
  wire [31:0] x777_x397_D31_number; // @[package.scala 96:25:@60865.4 package.scala 96:25:@60866.4]
  wire [31:0] x778_x399_sum_D26_number; // @[package.scala 96:25:@60874.4 package.scala 96:25:@60875.4]
  wire [31:0] x781_x389_D32_number; // @[package.scala 96:25:@60945.4 package.scala 96:25:@60946.4]
  wire [31:0] x782_x393_sum_D27_number; // @[package.scala 96:25:@60954.4 package.scala 96:25:@60955.4]
  wire [31:0] x441_sum_number; // @[Math.scala 154:22:@61064.4 Math.scala 155:14:@61065.4]
  wire [31:0] x785_x439_D5_number; // @[package.scala 96:25:@61073.4 package.scala 96:25:@61074.4]
  wire [31:0] x450_sum_number; // @[Math.scala 154:22:@61172.4 Math.scala 155:14:@61173.4]
  wire [31:0] x787_x448_D5_number; // @[package.scala 96:25:@61181.4 package.scala 96:25:@61182.4]
  wire [31:0] x461_sum_number; // @[Math.scala 154:22:@61349.4 Math.scala 155:14:@61350.4]
  wire [31:0] x792_x731_D20_number; // @[package.scala 96:25:@61367.4 package.scala 96:25:@61368.4]
  wire [31:0] x466_sum_number; // @[Math.scala 154:22:@61416.4 Math.scala 155:14:@61417.4]
  wire [31:0] x471_sum_number; // @[Math.scala 154:22:@61474.4 Math.scala 155:14:@61475.4]
  wire [31:0] x801_x476_sum_D1_number; // @[package.scala 96:25:@61570.4 package.scala 96:25:@61571.4]
  wire [31:0] x481_sum_number; // @[Math.scala 154:22:@61610.4 Math.scala 155:14:@61611.4]
  wire [31:0] x486_sum_number; // @[Math.scala 154:22:@61659.4 Math.scala 155:14:@61660.4]
  wire [31:0] x497_sum_number; // @[Math.scala 154:22:@61818.4 Math.scala 155:14:@61819.4]
  wire [31:0] x806_x736_D20_number; // @[package.scala 96:25:@61836.4 package.scala 96:25:@61837.4]
  wire [31:0] x502_sum_number; // @[Math.scala 154:22:@61876.4 Math.scala 155:14:@61877.4]
  wire [31:0] x507_sum_number; // @[Math.scala 154:22:@61925.4 Math.scala 155:14:@61926.4]
  wire [31:0] x811_x512_sum_D1_number; // @[package.scala 96:25:@62003.4 package.scala 96:25:@62004.4]
  wire [31:0] x517_sum_number; // @[Math.scala 154:22:@62043.4 Math.scala 155:14:@62044.4]
  wire [31:0] x522_sum_number; // @[Math.scala 154:22:@62092.4 Math.scala 155:14:@62093.4]
  wire [31:0] x819_x389_D51_number; // @[package.scala 96:25:@62983.4 package.scala 96:25:@62984.4]
  wire [31:0] x822_x393_sum_D46_number; // @[package.scala 96:25:@63010.4 package.scala 96:25:@63011.4]
  wire [31:0] x823_x726_D67_number; // @[package.scala 96:25:@63019.4 package.scala 96:25:@63020.4]
  wire [31:0] x824_x397_D50_number; // @[package.scala 96:25:@63051.4 package.scala 96:25:@63052.4]
  wire [31:0] x825_x399_sum_D45_number; // @[package.scala 96:25:@63060.4 package.scala 96:25:@63061.4]
  wire [31:0] x827_x403_D50_number; // @[package.scala 96:25:@63101.4 package.scala 96:25:@63102.4]
  wire [31:0] x828_x405_sum_D45_number; // @[package.scala 96:25:@63110.4 package.scala 96:25:@63111.4]
  wire [31:0] x830_x411_sum_D45_number; // @[package.scala 96:25:@63151.4 package.scala 96:25:@63152.4]
  wire [31:0] x831_x409_D50_number; // @[package.scala 96:25:@63160.4 package.scala 96:25:@63161.4]
  wire [31:0] x835_x411_sum_D46_number; // @[package.scala 96:25:@63219.4 package.scala 96:25:@63220.4]
  wire [31:0] x837_x726_D68_number; // @[package.scala 96:25:@63237.4 package.scala 96:25:@63238.4]
  wire [31:0] x838_x409_D51_number; // @[package.scala 96:25:@63246.4 package.scala 96:25:@63247.4]
  wire [31:0] x839_x403_D51_number; // @[package.scala 96:25:@63279.4 package.scala 96:25:@63280.4]
  wire [31:0] x840_x405_sum_D46_number; // @[package.scala 96:25:@63288.4 package.scala 96:25:@63289.4]
  wire [31:0] x842_x397_D51_number; // @[package.scala 96:25:@63330.4 package.scala 96:25:@63331.4]
  wire [31:0] x843_x399_sum_D46_number; // @[package.scala 96:25:@63339.4 package.scala 96:25:@63340.4]
  wire [31:0] x845_x389_D52_number; // @[package.scala 96:25:@63381.4 package.scala 96:25:@63382.4]
  wire [31:0] x846_x393_sum_D47_number; // @[package.scala 96:25:@63390.4 package.scala 96:25:@63391.4]
  wire [31:0] x848_x439_D25_number; // @[package.scala 96:25:@63432.4 package.scala 96:25:@63433.4]
  wire [31:0] x850_x441_sum_D20_number; // @[package.scala 96:25:@63450.4 package.scala 96:25:@63451.4]
  wire [31:0] x851_x461_sum_D20_number; // @[package.scala 96:25:@63483.4 package.scala 96:25:@63484.4]
  wire [31:0] x853_x731_D40_number; // @[package.scala 96:25:@63501.4 package.scala 96:25:@63502.4]
  wire [31:0] x854_x466_sum_D20_number; // @[package.scala 96:25:@63534.4 package.scala 96:25:@63535.4]
  wire [31:0] x856_x471_sum_D20_number; // @[package.scala 96:25:@63576.4 package.scala 96:25:@63577.4]
  wire [31:0] x859_x476_sum_D21_number; // @[package.scala 96:25:@63627.4 package.scala 96:25:@63628.4]
  wire [31:0] x860_x481_sum_D20_number; // @[package.scala 96:25:@63660.4 package.scala 96:25:@63661.4]
  _ _ ( // @[Math.scala 720:24:@59827.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@59839.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@59862.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x383_lb_0 x383_lb_0 ( // @[m_x383_lb_0.scala 47:17:@59872.4]
    .clock(x383_lb_0_clock),
    .reset(x383_lb_0_reset),
    .io_rPort_17_banks_1(x383_lb_0_io_rPort_17_banks_1),
    .io_rPort_17_banks_0(x383_lb_0_io_rPort_17_banks_0),
    .io_rPort_17_ofs_0(x383_lb_0_io_rPort_17_ofs_0),
    .io_rPort_17_en_0(x383_lb_0_io_rPort_17_en_0),
    .io_rPort_17_backpressure(x383_lb_0_io_rPort_17_backpressure),
    .io_rPort_17_output_0(x383_lb_0_io_rPort_17_output_0),
    .io_rPort_16_banks_1(x383_lb_0_io_rPort_16_banks_1),
    .io_rPort_16_banks_0(x383_lb_0_io_rPort_16_banks_0),
    .io_rPort_16_ofs_0(x383_lb_0_io_rPort_16_ofs_0),
    .io_rPort_16_en_0(x383_lb_0_io_rPort_16_en_0),
    .io_rPort_16_backpressure(x383_lb_0_io_rPort_16_backpressure),
    .io_rPort_16_output_0(x383_lb_0_io_rPort_16_output_0),
    .io_rPort_15_banks_1(x383_lb_0_io_rPort_15_banks_1),
    .io_rPort_15_banks_0(x383_lb_0_io_rPort_15_banks_0),
    .io_rPort_15_ofs_0(x383_lb_0_io_rPort_15_ofs_0),
    .io_rPort_15_en_0(x383_lb_0_io_rPort_15_en_0),
    .io_rPort_15_backpressure(x383_lb_0_io_rPort_15_backpressure),
    .io_rPort_15_output_0(x383_lb_0_io_rPort_15_output_0),
    .io_rPort_14_banks_1(x383_lb_0_io_rPort_14_banks_1),
    .io_rPort_14_banks_0(x383_lb_0_io_rPort_14_banks_0),
    .io_rPort_14_ofs_0(x383_lb_0_io_rPort_14_ofs_0),
    .io_rPort_14_en_0(x383_lb_0_io_rPort_14_en_0),
    .io_rPort_14_backpressure(x383_lb_0_io_rPort_14_backpressure),
    .io_rPort_14_output_0(x383_lb_0_io_rPort_14_output_0),
    .io_rPort_13_banks_1(x383_lb_0_io_rPort_13_banks_1),
    .io_rPort_13_banks_0(x383_lb_0_io_rPort_13_banks_0),
    .io_rPort_13_ofs_0(x383_lb_0_io_rPort_13_ofs_0),
    .io_rPort_13_en_0(x383_lb_0_io_rPort_13_en_0),
    .io_rPort_13_backpressure(x383_lb_0_io_rPort_13_backpressure),
    .io_rPort_13_output_0(x383_lb_0_io_rPort_13_output_0),
    .io_rPort_12_banks_1(x383_lb_0_io_rPort_12_banks_1),
    .io_rPort_12_banks_0(x383_lb_0_io_rPort_12_banks_0),
    .io_rPort_12_ofs_0(x383_lb_0_io_rPort_12_ofs_0),
    .io_rPort_12_en_0(x383_lb_0_io_rPort_12_en_0),
    .io_rPort_12_backpressure(x383_lb_0_io_rPort_12_backpressure),
    .io_rPort_12_output_0(x383_lb_0_io_rPort_12_output_0),
    .io_rPort_11_banks_1(x383_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x383_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x383_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x383_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x383_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x383_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x383_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x383_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x383_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x383_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x383_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x383_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x383_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x383_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x383_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x383_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x383_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x383_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x383_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x383_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x383_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x383_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x383_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x383_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x383_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x383_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x383_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x383_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x383_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x383_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x383_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x383_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x383_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x383_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x383_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x383_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x383_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x383_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x383_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x383_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x383_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x383_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x383_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x383_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x383_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x383_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x383_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x383_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x383_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x383_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x383_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x383_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x383_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x383_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x383_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x383_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x383_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x383_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x383_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x383_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x383_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x383_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x383_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x383_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x383_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x383_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x383_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x383_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x383_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x383_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x383_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x383_lb_0_io_rPort_0_output_0),
    .io_wPort_3_banks_1(x383_lb_0_io_wPort_3_banks_1),
    .io_wPort_3_banks_0(x383_lb_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x383_lb_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x383_lb_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x383_lb_0_io_wPort_3_en_0),
    .io_wPort_2_banks_1(x383_lb_0_io_wPort_2_banks_1),
    .io_wPort_2_banks_0(x383_lb_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x383_lb_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x383_lb_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x383_lb_0_io_wPort_2_en_0),
    .io_wPort_1_banks_1(x383_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x383_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x383_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x383_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x383_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x383_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x383_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x383_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x383_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x383_lb_0_io_wPort_0_en_0)
  );
  x384_lb2_0 x384_lb2_0 ( // @[m_x384_lb2_0.scala 39:17:@60017.4]
    .clock(x384_lb2_0_clock),
    .reset(x384_lb2_0_reset),
    .io_rPort_9_banks_1(x384_lb2_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x384_lb2_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x384_lb2_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x384_lb2_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x384_lb2_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x384_lb2_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x384_lb2_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x384_lb2_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x384_lb2_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x384_lb2_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x384_lb2_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x384_lb2_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x384_lb2_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x384_lb2_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x384_lb2_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x384_lb2_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x384_lb2_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x384_lb2_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x384_lb2_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x384_lb2_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x384_lb2_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x384_lb2_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x384_lb2_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x384_lb2_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x384_lb2_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x384_lb2_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x384_lb2_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x384_lb2_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x384_lb2_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x384_lb2_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x384_lb2_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x384_lb2_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x384_lb2_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x384_lb2_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x384_lb2_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x384_lb2_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x384_lb2_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x384_lb2_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x384_lb2_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x384_lb2_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x384_lb2_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x384_lb2_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x384_lb2_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x384_lb2_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x384_lb2_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x384_lb2_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x384_lb2_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x384_lb2_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x384_lb2_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x384_lb2_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x384_lb2_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x384_lb2_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x384_lb2_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x384_lb2_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x384_lb2_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x384_lb2_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x384_lb2_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x384_lb2_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x384_lb2_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x384_lb2_0_io_rPort_0_output_0),
    .io_wPort_3_banks_1(x384_lb2_0_io_wPort_3_banks_1),
    .io_wPort_3_banks_0(x384_lb2_0_io_wPort_3_banks_0),
    .io_wPort_3_ofs_0(x384_lb2_0_io_wPort_3_ofs_0),
    .io_wPort_3_data_0(x384_lb2_0_io_wPort_3_data_0),
    .io_wPort_3_en_0(x384_lb2_0_io_wPort_3_en_0),
    .io_wPort_2_banks_1(x384_lb2_0_io_wPort_2_banks_1),
    .io_wPort_2_banks_0(x384_lb2_0_io_wPort_2_banks_0),
    .io_wPort_2_ofs_0(x384_lb2_0_io_wPort_2_ofs_0),
    .io_wPort_2_data_0(x384_lb2_0_io_wPort_2_data_0),
    .io_wPort_2_en_0(x384_lb2_0_io_wPort_2_en_0),
    .io_wPort_1_banks_1(x384_lb2_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x384_lb2_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x384_lb2_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x384_lb2_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x384_lb2_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x384_lb2_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x384_lb2_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x384_lb2_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x384_lb2_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x384_lb2_0_io_wPort_0_en_0)
  );
  x389 x389_1 ( // @[Math.scala 366:24:@60152.4]
    .clock(x389_1_clock),
    .io_a(x389_1_io_a),
    .io_flow(x389_1_io_flow),
    .io_result(x389_1_io_result)
  );
  x356_sum x729_sum_1 ( // @[Math.scala 150:24:@60189.4]
    .clock(x729_sum_1_clock),
    .reset(x729_sum_1_reset),
    .io_a(x729_sum_1_io_a),
    .io_b(x729_sum_1_io_b),
    .io_flow(x729_sum_1_io_flow),
    .io_result(x729_sum_1_io_result)
  );
  x392_div x392_div_1 ( // @[Math.scala 327:24:@60201.4]
    .clock(x392_div_1_clock),
    .io_a(x392_div_1_io_a),
    .io_flow(x392_div_1_io_flow),
    .io_result(x392_div_1_io_result)
  );
  RetimeWrapper_438 RetimeWrapper_1 ( // @[package.scala 93:22:@60211.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x356_sum x393_sum_1 ( // @[Math.scala 150:24:@60220.4]
    .clock(x393_sum_1_clock),
    .reset(x393_sum_1_reset),
    .io_a(x393_sum_1_io_a),
    .io_b(x393_sum_1_io_b),
    .io_flow(x393_sum_1_io_flow),
    .io_result(x393_sum_1_io_result)
  );
  RetimeWrapper_440 RetimeWrapper_2 ( // @[package.scala 93:22:@60230.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_441 RetimeWrapper_3 ( // @[package.scala 93:22:@60239.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_440 RetimeWrapper_4 ( // @[package.scala 93:22:@60248.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_443 RetimeWrapper_5 ( // @[package.scala 93:22:@60257.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_444 RetimeWrapper_6 ( // @[package.scala 93:22:@60266.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_445 RetimeWrapper_7 ( // @[package.scala 93:22:@60275.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_440 RetimeWrapper_8 ( // @[package.scala 93:22:@60286.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x356_sum x395_rdcol_1 ( // @[Math.scala 150:24:@60309.4]
    .clock(x395_rdcol_1_clock),
    .reset(x395_rdcol_1_reset),
    .io_a(x395_rdcol_1_io_a),
    .io_b(x395_rdcol_1_io_b),
    .io_flow(x395_rdcol_1_io_flow),
    .io_result(x395_rdcol_1_io_result)
  );
  x389 x397_1 ( // @[Math.scala 366:24:@60323.4]
    .clock(x397_1_clock),
    .io_a(x397_1_io_a),
    .io_flow(x397_1_io_flow),
    .io_result(x397_1_io_result)
  );
  x392_div x398_div_1 ( // @[Math.scala 327:24:@60335.4]
    .clock(x398_div_1_clock),
    .io_a(x398_div_1_io_a),
    .io_flow(x398_div_1_io_flow),
    .io_result(x398_div_1_io_result)
  );
  RetimeWrapper_448 RetimeWrapper_9 ( // @[package.scala 93:22:@60345.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  x356_sum x399_sum_1 ( // @[Math.scala 150:24:@60354.4]
    .clock(x399_sum_1_clock),
    .reset(x399_sum_1_reset),
    .io_a(x399_sum_1_io_a),
    .io_b(x399_sum_1_io_b),
    .io_flow(x399_sum_1_io_flow),
    .io_result(x399_sum_1_io_result)
  );
  RetimeWrapper_450 RetimeWrapper_10 ( // @[package.scala 93:22:@60364.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_444 RetimeWrapper_11 ( // @[package.scala 93:22:@60373.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_452 RetimeWrapper_12 ( // @[package.scala 93:22:@60382.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_440 RetimeWrapper_13 ( // @[package.scala 93:22:@60393.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  x356_sum x401_rdcol_1 ( // @[Math.scala 150:24:@60416.4]
    .clock(x401_rdcol_1_clock),
    .reset(x401_rdcol_1_reset),
    .io_a(x401_rdcol_1_io_a),
    .io_b(x401_rdcol_1_io_b),
    .io_flow(x401_rdcol_1_io_flow),
    .io_result(x401_rdcol_1_io_result)
  );
  x389 x403_1 ( // @[Math.scala 366:24:@60430.4]
    .clock(x403_1_clock),
    .io_a(x403_1_io_a),
    .io_flow(x403_1_io_flow),
    .io_result(x403_1_io_result)
  );
  x392_div x404_div_1 ( // @[Math.scala 327:24:@60442.4]
    .clock(x404_div_1_clock),
    .io_a(x404_div_1_io_a),
    .io_flow(x404_div_1_io_flow),
    .io_result(x404_div_1_io_result)
  );
  x356_sum x405_sum_1 ( // @[Math.scala 150:24:@60452.4]
    .clock(x405_sum_1_clock),
    .reset(x405_sum_1_reset),
    .io_a(x405_sum_1_io_a),
    .io_b(x405_sum_1_io_b),
    .io_flow(x405_sum_1_io_flow),
    .io_result(x405_sum_1_io_result)
  );
  RetimeWrapper_450 RetimeWrapper_14 ( // @[package.scala 93:22:@60462.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_444 RetimeWrapper_15 ( // @[package.scala 93:22:@60471.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_452 RetimeWrapper_16 ( // @[package.scala 93:22:@60480.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_440 RetimeWrapper_17 ( // @[package.scala 93:22:@60491.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  x356_sum x407_rdcol_1 ( // @[Math.scala 150:24:@60514.4]
    .clock(x407_rdcol_1_clock),
    .reset(x407_rdcol_1_reset),
    .io_a(x407_rdcol_1_io_a),
    .io_b(x407_rdcol_1_io_b),
    .io_flow(x407_rdcol_1_io_flow),
    .io_result(x407_rdcol_1_io_result)
  );
  x389 x409_1 ( // @[Math.scala 366:24:@60528.4]
    .clock(x409_1_clock),
    .io_a(x409_1_io_a),
    .io_flow(x409_1_io_flow),
    .io_result(x409_1_io_result)
  );
  x392_div x410_div_1 ( // @[Math.scala 327:24:@60540.4]
    .clock(x410_div_1_clock),
    .io_a(x410_div_1_io_a),
    .io_flow(x410_div_1_io_flow),
    .io_result(x410_div_1_io_result)
  );
  x356_sum x411_sum_1 ( // @[Math.scala 150:24:@60550.4]
    .clock(x411_sum_1_clock),
    .reset(x411_sum_1_reset),
    .io_a(x411_sum_1_io_a),
    .io_b(x411_sum_1_io_b),
    .io_flow(x411_sum_1_io_flow),
    .io_result(x411_sum_1_io_result)
  );
  RetimeWrapper_444 RetimeWrapper_18 ( // @[package.scala 93:22:@60560.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_452 RetimeWrapper_19 ( // @[package.scala 93:22:@60569.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_450 RetimeWrapper_20 ( // @[package.scala 93:22:@60578.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_440 RetimeWrapper_21 ( // @[package.scala 93:22:@60589.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_22 ( // @[package.scala 93:22:@60610.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper RetimeWrapper_23 ( // @[package.scala 93:22:@60626.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_24 ( // @[package.scala 93:22:@60635.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper RetimeWrapper_25 ( // @[package.scala 93:22:@60649.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper RetimeWrapper_26 ( // @[package.scala 93:22:@60658.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_27 ( // @[package.scala 93:22:@60673.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_472 RetimeWrapper_28 ( // @[package.scala 93:22:@60682.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_29 ( // @[package.scala 93:22:@60691.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_30 ( // @[package.scala 93:22:@60700.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_475 RetimeWrapper_31 ( // @[package.scala 93:22:@60709.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_476 RetimeWrapper_32 ( // @[package.scala 93:22:@60718.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_33 ( // @[package.scala 93:22:@60730.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_34 ( // @[package.scala 93:22:@60751.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper RetimeWrapper_35 ( // @[package.scala 93:22:@60765.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_476 RetimeWrapper_36 ( // @[package.scala 93:22:@60780.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_37 ( // @[package.scala 93:22:@60789.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_472 RetimeWrapper_38 ( // @[package.scala 93:22:@60798.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_39 ( // @[package.scala 93:22:@60810.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_40 ( // @[package.scala 93:22:@60831.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@60845.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_476 RetimeWrapper_42 ( // @[package.scala 93:22:@60860.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_43 ( // @[package.scala 93:22:@60869.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_472 RetimeWrapper_44 ( // @[package.scala 93:22:@60878.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_45 ( // @[package.scala 93:22:@60890.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_46 ( // @[package.scala 93:22:@60911.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper RetimeWrapper_47 ( // @[package.scala 93:22:@60925.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_492 RetimeWrapper_48 ( // @[package.scala 93:22:@60940.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_493 RetimeWrapper_49 ( // @[package.scala 93:22:@60949.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_494 RetimeWrapper_50 ( // @[package.scala 93:22:@60958.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_51 ( // @[package.scala 93:22:@60970.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  x356_sum x435_rdcol_1 ( // @[Math.scala 150:24:@60993.4]
    .clock(x435_rdcol_1_clock),
    .reset(x435_rdcol_1_reset),
    .io_a(x435_rdcol_1_io_a),
    .io_b(x435_rdcol_1_io_b),
    .io_flow(x435_rdcol_1_io_flow),
    .io_result(x435_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_52 ( // @[package.scala 93:22:@61008.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  x389 x439_1 ( // @[Math.scala 366:24:@61027.4]
    .clock(x439_1_clock),
    .io_a(x439_1_io_a),
    .io_flow(x439_1_io_flow),
    .io_result(x439_1_io_result)
  );
  x392_div x440_div_1 ( // @[Math.scala 327:24:@61039.4]
    .clock(x440_div_1_clock),
    .io_a(x440_div_1_io_a),
    .io_flow(x440_div_1_io_flow),
    .io_result(x440_div_1_io_result)
  );
  RetimeWrapper_498 RetimeWrapper_53 ( // @[package.scala 93:22:@61049.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x356_sum x441_sum_1 ( // @[Math.scala 150:24:@61058.4]
    .clock(x441_sum_1_clock),
    .reset(x441_sum_1_reset),
    .io_a(x441_sum_1_io_a),
    .io_b(x441_sum_1_io_b),
    .io_flow(x441_sum_1_io_flow),
    .io_result(x441_sum_1_io_result)
  );
  RetimeWrapper_500 RetimeWrapper_54 ( // @[package.scala 93:22:@61068.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_472 RetimeWrapper_55 ( // @[package.scala 93:22:@61077.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_56 ( // @[package.scala 93:22:@61089.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  x356_sum x444_rdcol_1 ( // @[Math.scala 150:24:@61112.4]
    .clock(x444_rdcol_1_clock),
    .reset(x444_rdcol_1_reset),
    .io_a(x444_rdcol_1_io_a),
    .io_b(x444_rdcol_1_io_b),
    .io_flow(x444_rdcol_1_io_flow),
    .io_result(x444_rdcol_1_io_result)
  );
  RetimeWrapper RetimeWrapper_57 ( // @[package.scala 93:22:@61127.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x389 x448_1 ( // @[Math.scala 366:24:@61144.4]
    .clock(x448_1_clock),
    .io_a(x448_1_io_a),
    .io_flow(x448_1_io_flow),
    .io_result(x448_1_io_result)
  );
  x392_div x449_div_1 ( // @[Math.scala 327:24:@61156.4]
    .clock(x449_div_1_clock),
    .io_a(x449_div_1_io_a),
    .io_flow(x449_div_1_io_flow),
    .io_result(x449_div_1_io_result)
  );
  x356_sum x450_sum_1 ( // @[Math.scala 150:24:@61166.4]
    .clock(x450_sum_1_clock),
    .reset(x450_sum_1_reset),
    .io_a(x450_sum_1_io_a),
    .io_b(x450_sum_1_io_b),
    .io_flow(x450_sum_1_io_flow),
    .io_result(x450_sum_1_io_result)
  );
  RetimeWrapper_500 RetimeWrapper_58 ( // @[package.scala 93:22:@61176.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_472 RetimeWrapper_59 ( // @[package.scala 93:22:@61185.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_60 ( // @[package.scala 93:22:@61197.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  x720_sub x453_rdrow_1 ( // @[Math.scala 191:24:@61220.4]
    .clock(x453_rdrow_1_clock),
    .reset(x453_rdrow_1_reset),
    .io_a(x453_rdrow_1_io_a),
    .io_b(x453_rdrow_1_io_b),
    .io_flow(x453_rdrow_1_io_flow),
    .io_result(x453_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_61 ( // @[package.scala 93:22:@61246.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_62 ( // @[package.scala 93:22:@61268.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_63 ( // @[package.scala 93:22:@61294.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  x356_sum x734_sum_1 ( // @[Math.scala 150:24:@61315.4]
    .clock(x734_sum_1_clock),
    .reset(x734_sum_1_reset),
    .io_a(x734_sum_1_io_a),
    .io_b(x734_sum_1_io_b),
    .io_flow(x734_sum_1_io_flow),
    .io_result(x734_sum_1_io_result)
  );
  RetimeWrapper_466 RetimeWrapper_64 ( // @[package.scala 93:22:@61325.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_515 RetimeWrapper_65 ( // @[package.scala 93:22:@61334.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  x356_sum x461_sum_1 ( // @[Math.scala 150:24:@61343.4]
    .clock(x461_sum_1_clock),
    .reset(x461_sum_1_reset),
    .io_a(x461_sum_1_io_a),
    .io_b(x461_sum_1_io_b),
    .io_flow(x461_sum_1_io_flow),
    .io_result(x461_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_66 ( // @[package.scala 93:22:@61353.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_67 ( // @[package.scala 93:22:@61362.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_68 ( // @[package.scala 93:22:@61374.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_69 ( // @[package.scala 93:22:@61401.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  x356_sum x466_sum_1 ( // @[Math.scala 150:24:@61410.4]
    .clock(x466_sum_1_clock),
    .reset(x466_sum_1_reset),
    .io_a(x466_sum_1_io_a),
    .io_b(x466_sum_1_io_b),
    .io_flow(x466_sum_1_io_flow),
    .io_result(x466_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_70 ( // @[package.scala 93:22:@61420.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_71 ( // @[package.scala 93:22:@61432.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_72 ( // @[package.scala 93:22:@61459.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  x356_sum x471_sum_1 ( // @[Math.scala 150:24:@61468.4]
    .clock(x471_sum_1_clock),
    .reset(x471_sum_1_reset),
    .io_a(x471_sum_1_io_a),
    .io_b(x471_sum_1_io_b),
    .io_flow(x471_sum_1_io_flow),
    .io_result(x471_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_73 ( // @[package.scala 93:22:@61478.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_74 ( // @[package.scala 93:22:@61490.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper RetimeWrapper_75 ( // @[package.scala 93:22:@61511.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_466 RetimeWrapper_76 ( // @[package.scala 93:22:@61526.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_530 RetimeWrapper_77 ( // @[package.scala 93:22:@61535.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  x356_sum x476_sum_1 ( // @[Math.scala 150:24:@61546.4]
    .clock(x476_sum_1_clock),
    .reset(x476_sum_1_reset),
    .io_a(x476_sum_1_io_a),
    .io_b(x476_sum_1_io_b),
    .io_flow(x476_sum_1_io_flow),
    .io_result(x476_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_78 ( // @[package.scala 93:22:@61556.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_79 ( // @[package.scala 93:22:@61565.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_80 ( // @[package.scala 93:22:@61577.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  x356_sum x481_sum_1 ( // @[Math.scala 150:24:@61604.4]
    .clock(x481_sum_1_clock),
    .reset(x481_sum_1_reset),
    .io_a(x481_sum_1_io_a),
    .io_b(x481_sum_1_io_b),
    .io_flow(x481_sum_1_io_flow),
    .io_result(x481_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_81 ( // @[package.scala 93:22:@61614.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_82 ( // @[package.scala 93:22:@61626.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  x356_sum x486_sum_1 ( // @[Math.scala 150:24:@61653.4]
    .clock(x486_sum_1_clock),
    .reset(x486_sum_1_reset),
    .io_a(x486_sum_1_io_a),
    .io_b(x486_sum_1_io_b),
    .io_flow(x486_sum_1_io_flow),
    .io_result(x486_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_83 ( // @[package.scala 93:22:@61663.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_84 ( // @[package.scala 93:22:@61675.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  x720_sub x489_rdrow_1 ( // @[Math.scala 191:24:@61698.4]
    .clock(x489_rdrow_1_clock),
    .reset(x489_rdrow_1_reset),
    .io_a(x489_rdrow_1_io_a),
    .io_b(x489_rdrow_1_io_b),
    .io_flow(x489_rdrow_1_io_flow),
    .io_result(x489_rdrow_1_io_result)
  );
  RetimeWrapper RetimeWrapper_85 ( // @[package.scala 93:22:@61724.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_86 ( // @[package.scala 93:22:@61746.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_87 ( // @[package.scala 93:22:@61772.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  x356_sum x739_sum_1 ( // @[Math.scala 150:24:@61793.4]
    .clock(x739_sum_1_clock),
    .reset(x739_sum_1_reset),
    .io_a(x739_sum_1_io_a),
    .io_b(x739_sum_1_io_b),
    .io_flow(x739_sum_1_io_flow),
    .io_result(x739_sum_1_io_result)
  );
  RetimeWrapper_515 RetimeWrapper_88 ( // @[package.scala 93:22:@61803.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  x356_sum x497_sum_1 ( // @[Math.scala 150:24:@61812.4]
    .clock(x497_sum_1_clock),
    .reset(x497_sum_1_reset),
    .io_a(x497_sum_1_io_a),
    .io_b(x497_sum_1_io_b),
    .io_flow(x497_sum_1_io_flow),
    .io_result(x497_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_89 ( // @[package.scala 93:22:@61822.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_90 ( // @[package.scala 93:22:@61831.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_91 ( // @[package.scala 93:22:@61843.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  x356_sum x502_sum_1 ( // @[Math.scala 150:24:@61870.4]
    .clock(x502_sum_1_clock),
    .reset(x502_sum_1_reset),
    .io_a(x502_sum_1_io_a),
    .io_b(x502_sum_1_io_b),
    .io_flow(x502_sum_1_io_flow),
    .io_result(x502_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_92 ( // @[package.scala 93:22:@61880.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_93 ( // @[package.scala 93:22:@61892.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  x356_sum x507_sum_1 ( // @[Math.scala 150:24:@61919.4]
    .clock(x507_sum_1_clock),
    .reset(x507_sum_1_reset),
    .io_a(x507_sum_1_io_a),
    .io_b(x507_sum_1_io_b),
    .io_flow(x507_sum_1_io_flow),
    .io_result(x507_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_94 ( // @[package.scala 93:22:@61929.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_95 ( // @[package.scala 93:22:@61941.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  RetimeWrapper_530 RetimeWrapper_96 ( // @[package.scala 93:22:@61968.4]
    .clock(RetimeWrapper_96_clock),
    .reset(RetimeWrapper_96_reset),
    .io_flow(RetimeWrapper_96_io_flow),
    .io_in(RetimeWrapper_96_io_in),
    .io_out(RetimeWrapper_96_io_out)
  );
  x356_sum x512_sum_1 ( // @[Math.scala 150:24:@61979.4]
    .clock(x512_sum_1_clock),
    .reset(x512_sum_1_reset),
    .io_a(x512_sum_1_io_a),
    .io_b(x512_sum_1_io_b),
    .io_flow(x512_sum_1_io_flow),
    .io_result(x512_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_97 ( // @[package.scala 93:22:@61989.4]
    .clock(RetimeWrapper_97_clock),
    .reset(RetimeWrapper_97_reset),
    .io_flow(RetimeWrapper_97_io_flow),
    .io_in(RetimeWrapper_97_io_in),
    .io_out(RetimeWrapper_97_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_98 ( // @[package.scala 93:22:@61998.4]
    .clock(RetimeWrapper_98_clock),
    .reset(RetimeWrapper_98_reset),
    .io_flow(RetimeWrapper_98_io_flow),
    .io_in(RetimeWrapper_98_io_in),
    .io_out(RetimeWrapper_98_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_99 ( // @[package.scala 93:22:@62010.4]
    .clock(RetimeWrapper_99_clock),
    .reset(RetimeWrapper_99_reset),
    .io_flow(RetimeWrapper_99_io_flow),
    .io_in(RetimeWrapper_99_io_in),
    .io_out(RetimeWrapper_99_io_out)
  );
  x356_sum x517_sum_1 ( // @[Math.scala 150:24:@62037.4]
    .clock(x517_sum_1_clock),
    .reset(x517_sum_1_reset),
    .io_a(x517_sum_1_io_a),
    .io_b(x517_sum_1_io_b),
    .io_flow(x517_sum_1_io_flow),
    .io_result(x517_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_100 ( // @[package.scala 93:22:@62047.4]
    .clock(RetimeWrapper_100_clock),
    .reset(RetimeWrapper_100_reset),
    .io_flow(RetimeWrapper_100_io_flow),
    .io_in(RetimeWrapper_100_io_in),
    .io_out(RetimeWrapper_100_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_101 ( // @[package.scala 93:22:@62059.4]
    .clock(RetimeWrapper_101_clock),
    .reset(RetimeWrapper_101_reset),
    .io_flow(RetimeWrapper_101_io_flow),
    .io_in(RetimeWrapper_101_io_in),
    .io_out(RetimeWrapper_101_io_out)
  );
  x356_sum x522_sum_1 ( // @[Math.scala 150:24:@62086.4]
    .clock(x522_sum_1_clock),
    .reset(x522_sum_1_reset),
    .io_a(x522_sum_1_io_a),
    .io_b(x522_sum_1_io_b),
    .io_flow(x522_sum_1_io_flow),
    .io_result(x522_sum_1_io_result)
  );
  RetimeWrapper_472 RetimeWrapper_102 ( // @[package.scala 93:22:@62096.4]
    .clock(RetimeWrapper_102_clock),
    .reset(RetimeWrapper_102_reset),
    .io_flow(RetimeWrapper_102_io_flow),
    .io_in(RetimeWrapper_102_io_in),
    .io_out(RetimeWrapper_102_io_out)
  );
  RetimeWrapper_471 RetimeWrapper_103 ( // @[package.scala 93:22:@62108.4]
    .clock(RetimeWrapper_103_clock),
    .reset(RetimeWrapper_103_reset),
    .io_flow(RetimeWrapper_103_io_flow),
    .io_in(RetimeWrapper_103_io_in),
    .io_out(RetimeWrapper_103_io_out)
  );
  x525 x525_1 ( // @[Math.scala 262:24:@62131.4]
    .clock(x525_1_clock),
    .io_a(x525_1_io_a),
    .io_b(x525_1_io_b),
    .io_flow(x525_1_io_flow),
    .io_result(x525_1_io_result)
  );
  x525 x526_1 ( // @[Math.scala 262:24:@62143.4]
    .clock(x526_1_clock),
    .io_a(x526_1_io_a),
    .io_b(x526_1_io_b),
    .io_flow(x526_1_io_flow),
    .io_result(x526_1_io_result)
  );
  x525 x527_1 ( // @[Math.scala 262:24:@62155.4]
    .clock(x527_1_clock),
    .io_a(x527_1_io_a),
    .io_b(x527_1_io_b),
    .io_flow(x527_1_io_flow),
    .io_result(x527_1_io_result)
  );
  x525 x528_1 ( // @[Math.scala 262:24:@62167.4]
    .clock(x528_1_clock),
    .io_a(x528_1_io_a),
    .io_b(x528_1_io_b),
    .io_flow(x528_1_io_flow),
    .io_result(x528_1_io_result)
  );
  x525 x529_1 ( // @[Math.scala 262:24:@62179.4]
    .clock(x529_1_clock),
    .io_a(x529_1_io_a),
    .io_b(x529_1_io_b),
    .io_flow(x529_1_io_flow),
    .io_result(x529_1_io_result)
  );
  x525 x530_1 ( // @[Math.scala 262:24:@62191.4]
    .clock(x530_1_clock),
    .io_a(x530_1_io_a),
    .io_b(x530_1_io_b),
    .io_flow(x530_1_io_flow),
    .io_result(x530_1_io_result)
  );
  x525 x531_1 ( // @[Math.scala 262:24:@62203.4]
    .clock(x531_1_clock),
    .io_a(x531_1_io_a),
    .io_b(x531_1_io_b),
    .io_flow(x531_1_io_flow),
    .io_result(x531_1_io_result)
  );
  x525 x532_1 ( // @[Math.scala 262:24:@62215.4]
    .clock(x532_1_clock),
    .io_a(x532_1_io_a),
    .io_b(x532_1_io_b),
    .io_flow(x532_1_io_flow),
    .io_result(x532_1_io_result)
  );
  x525 x533_1 ( // @[Math.scala 262:24:@62227.4]
    .clock(x533_1_clock),
    .io_a(x533_1_io_a),
    .io_b(x533_1_io_b),
    .io_flow(x533_1_io_flow),
    .io_result(x533_1_io_result)
  );
  x534_x7 x534_x7_1 ( // @[Math.scala 150:24:@62237.4]
    .clock(x534_x7_1_clock),
    .reset(x534_x7_1_reset),
    .io_a(x534_x7_1_io_a),
    .io_b(x534_x7_1_io_b),
    .io_flow(x534_x7_1_io_flow),
    .io_result(x534_x7_1_io_result)
  );
  x534_x7 x535_x8_1 ( // @[Math.scala 150:24:@62247.4]
    .clock(x535_x8_1_clock),
    .reset(x535_x8_1_reset),
    .io_a(x535_x8_1_io_a),
    .io_b(x535_x8_1_io_b),
    .io_flow(x535_x8_1_io_flow),
    .io_result(x535_x8_1_io_result)
  );
  x534_x7 x536_x7_1 ( // @[Math.scala 150:24:@62257.4]
    .clock(x536_x7_1_clock),
    .reset(x536_x7_1_reset),
    .io_a(x536_x7_1_io_a),
    .io_b(x536_x7_1_io_b),
    .io_flow(x536_x7_1_io_flow),
    .io_result(x536_x7_1_io_result)
  );
  x534_x7 x537_x8_1 ( // @[Math.scala 150:24:@62267.4]
    .clock(x537_x8_1_clock),
    .reset(x537_x8_1_reset),
    .io_a(x537_x8_1_io_a),
    .io_b(x537_x8_1_io_b),
    .io_flow(x537_x8_1_io_flow),
    .io_result(x537_x8_1_io_result)
  );
  x534_x7 x538_x7_1 ( // @[Math.scala 150:24:@62277.4]
    .clock(x538_x7_1_clock),
    .reset(x538_x7_1_reset),
    .io_a(x538_x7_1_io_a),
    .io_b(x538_x7_1_io_b),
    .io_flow(x538_x7_1_io_flow),
    .io_result(x538_x7_1_io_result)
  );
  x534_x7 x539_x8_1 ( // @[Math.scala 150:24:@62287.4]
    .clock(x539_x8_1_clock),
    .reset(x539_x8_1_reset),
    .io_a(x539_x8_1_io_a),
    .io_b(x539_x8_1_io_b),
    .io_flow(x539_x8_1_io_flow),
    .io_result(x539_x8_1_io_result)
  );
  x534_x7 x540_x7_1 ( // @[Math.scala 150:24:@62297.4]
    .clock(x540_x7_1_clock),
    .reset(x540_x7_1_reset),
    .io_a(x540_x7_1_io_a),
    .io_b(x540_x7_1_io_b),
    .io_flow(x540_x7_1_io_flow),
    .io_result(x540_x7_1_io_result)
  );
  RetimeWrapper_443 RetimeWrapper_104 ( // @[package.scala 93:22:@62307.4]
    .clock(RetimeWrapper_104_clock),
    .reset(RetimeWrapper_104_reset),
    .io_flow(RetimeWrapper_104_io_flow),
    .io_in(RetimeWrapper_104_io_in),
    .io_out(RetimeWrapper_104_io_out)
  );
  x534_x7 x541_sum_1 ( // @[Math.scala 150:24:@62316.4]
    .clock(x541_sum_1_clock),
    .reset(x541_sum_1_reset),
    .io_a(x541_sum_1_io_a),
    .io_b(x541_sum_1_io_b),
    .io_flow(x541_sum_1_io_flow),
    .io_result(x541_sum_1_io_result)
  );
  x542 x542_1 ( // @[Math.scala 720:24:@62326.4]
    .io_b(x542_1_io_b),
    .io_result(x542_1_io_result)
  );
  x543_mul x543_mul_1 ( // @[Math.scala 262:24:@62337.4]
    .clock(x543_mul_1_clock),
    .io_a(x543_mul_1_io_a),
    .io_b(x543_mul_1_io_b),
    .io_flow(x543_mul_1_io_flow),
    .io_result(x543_mul_1_io_result)
  );
  x544 x544_1 ( // @[Math.scala 720:24:@62347.4]
    .io_b(x544_1_io_b),
    .io_result(x544_1_io_result)
  );
  x525 x545_1 ( // @[Math.scala 262:24:@62358.4]
    .clock(x545_1_clock),
    .io_a(x545_1_io_a),
    .io_b(x545_1_io_b),
    .io_flow(x545_1_io_flow),
    .io_result(x545_1_io_result)
  );
  x525 x546_1 ( // @[Math.scala 262:24:@62370.4]
    .clock(x546_1_clock),
    .io_a(x546_1_io_a),
    .io_b(x546_1_io_b),
    .io_flow(x546_1_io_flow),
    .io_result(x546_1_io_result)
  );
  x525 x547_1 ( // @[Math.scala 262:24:@62382.4]
    .clock(x547_1_clock),
    .io_a(x547_1_io_a),
    .io_b(x547_1_io_b),
    .io_flow(x547_1_io_flow),
    .io_result(x547_1_io_result)
  );
  x525 x548_1 ( // @[Math.scala 262:24:@62394.4]
    .clock(x548_1_clock),
    .io_a(x548_1_io_a),
    .io_b(x548_1_io_b),
    .io_flow(x548_1_io_flow),
    .io_result(x548_1_io_result)
  );
  x525 x549_1 ( // @[Math.scala 262:24:@62406.4]
    .clock(x549_1_clock),
    .io_a(x549_1_io_a),
    .io_b(x549_1_io_b),
    .io_flow(x549_1_io_flow),
    .io_result(x549_1_io_result)
  );
  x525 x550_1 ( // @[Math.scala 262:24:@62420.4]
    .clock(x550_1_clock),
    .io_a(x550_1_io_a),
    .io_b(x550_1_io_b),
    .io_flow(x550_1_io_flow),
    .io_result(x550_1_io_result)
  );
  x525 x551_1 ( // @[Math.scala 262:24:@62432.4]
    .clock(x551_1_clock),
    .io_a(x551_1_io_a),
    .io_b(x551_1_io_b),
    .io_flow(x551_1_io_flow),
    .io_result(x551_1_io_result)
  );
  x525 x552_1 ( // @[Math.scala 262:24:@62444.4]
    .clock(x552_1_clock),
    .io_a(x552_1_io_a),
    .io_b(x552_1_io_b),
    .io_flow(x552_1_io_flow),
    .io_result(x552_1_io_result)
  );
  x525 x553_1 ( // @[Math.scala 262:24:@62456.4]
    .clock(x553_1_clock),
    .io_a(x553_1_io_a),
    .io_b(x553_1_io_b),
    .io_flow(x553_1_io_flow),
    .io_result(x553_1_io_result)
  );
  x534_x7 x554_x7_1 ( // @[Math.scala 150:24:@62466.4]
    .clock(x554_x7_1_clock),
    .reset(x554_x7_1_reset),
    .io_a(x554_x7_1_io_a),
    .io_b(x554_x7_1_io_b),
    .io_flow(x554_x7_1_io_flow),
    .io_result(x554_x7_1_io_result)
  );
  x534_x7 x555_x8_1 ( // @[Math.scala 150:24:@62476.4]
    .clock(x555_x8_1_clock),
    .reset(x555_x8_1_reset),
    .io_a(x555_x8_1_io_a),
    .io_b(x555_x8_1_io_b),
    .io_flow(x555_x8_1_io_flow),
    .io_result(x555_x8_1_io_result)
  );
  x534_x7 x556_x7_1 ( // @[Math.scala 150:24:@62486.4]
    .clock(x556_x7_1_clock),
    .reset(x556_x7_1_reset),
    .io_a(x556_x7_1_io_a),
    .io_b(x556_x7_1_io_b),
    .io_flow(x556_x7_1_io_flow),
    .io_result(x556_x7_1_io_result)
  );
  x534_x7 x557_x8_1 ( // @[Math.scala 150:24:@62496.4]
    .clock(x557_x8_1_clock),
    .reset(x557_x8_1_reset),
    .io_a(x557_x8_1_io_a),
    .io_b(x557_x8_1_io_b),
    .io_flow(x557_x8_1_io_flow),
    .io_result(x557_x8_1_io_result)
  );
  x534_x7 x558_x7_1 ( // @[Math.scala 150:24:@62506.4]
    .clock(x558_x7_1_clock),
    .reset(x558_x7_1_reset),
    .io_a(x558_x7_1_io_a),
    .io_b(x558_x7_1_io_b),
    .io_flow(x558_x7_1_io_flow),
    .io_result(x558_x7_1_io_result)
  );
  x534_x7 x559_x8_1 ( // @[Math.scala 150:24:@62516.4]
    .clock(x559_x8_1_clock),
    .reset(x559_x8_1_reset),
    .io_a(x559_x8_1_io_a),
    .io_b(x559_x8_1_io_b),
    .io_flow(x559_x8_1_io_flow),
    .io_result(x559_x8_1_io_result)
  );
  x534_x7 x560_x7_1 ( // @[Math.scala 150:24:@62526.4]
    .clock(x560_x7_1_clock),
    .reset(x560_x7_1_reset),
    .io_a(x560_x7_1_io_a),
    .io_b(x560_x7_1_io_b),
    .io_flow(x560_x7_1_io_flow),
    .io_result(x560_x7_1_io_result)
  );
  RetimeWrapper_443 RetimeWrapper_105 ( // @[package.scala 93:22:@62536.4]
    .clock(RetimeWrapper_105_clock),
    .reset(RetimeWrapper_105_reset),
    .io_flow(RetimeWrapper_105_io_flow),
    .io_in(RetimeWrapper_105_io_in),
    .io_out(RetimeWrapper_105_io_out)
  );
  x534_x7 x561_sum_1 ( // @[Math.scala 150:24:@62545.4]
    .clock(x561_sum_1_clock),
    .reset(x561_sum_1_reset),
    .io_a(x561_sum_1_io_a),
    .io_b(x561_sum_1_io_b),
    .io_flow(x561_sum_1_io_flow),
    .io_result(x561_sum_1_io_result)
  );
  x542 x562_1 ( // @[Math.scala 720:24:@62555.4]
    .io_b(x562_1_io_b),
    .io_result(x562_1_io_result)
  );
  x543_mul x563_mul_1 ( // @[Math.scala 262:24:@62566.4]
    .clock(x563_mul_1_clock),
    .io_a(x563_mul_1_io_a),
    .io_b(x563_mul_1_io_b),
    .io_flow(x563_mul_1_io_flow),
    .io_result(x563_mul_1_io_result)
  );
  x544 x564_1 ( // @[Math.scala 720:24:@62576.4]
    .io_b(x564_1_io_b),
    .io_result(x564_1_io_result)
  );
  x525 x565_1 ( // @[Math.scala 262:24:@62587.4]
    .clock(x565_1_clock),
    .io_a(x565_1_io_a),
    .io_b(x565_1_io_b),
    .io_flow(x565_1_io_flow),
    .io_result(x565_1_io_result)
  );
  x525 x566_1 ( // @[Math.scala 262:24:@62599.4]
    .clock(x566_1_clock),
    .io_a(x566_1_io_a),
    .io_b(x566_1_io_b),
    .io_flow(x566_1_io_flow),
    .io_result(x566_1_io_result)
  );
  x525 x567_1 ( // @[Math.scala 262:24:@62611.4]
    .clock(x567_1_clock),
    .io_a(x567_1_io_a),
    .io_b(x567_1_io_b),
    .io_flow(x567_1_io_flow),
    .io_result(x567_1_io_result)
  );
  x525 x568_1 ( // @[Math.scala 262:24:@62623.4]
    .clock(x568_1_clock),
    .io_a(x568_1_io_a),
    .io_b(x568_1_io_b),
    .io_flow(x568_1_io_flow),
    .io_result(x568_1_io_result)
  );
  x525 x569_1 ( // @[Math.scala 262:24:@62635.4]
    .clock(x569_1_clock),
    .io_a(x569_1_io_a),
    .io_b(x569_1_io_b),
    .io_flow(x569_1_io_flow),
    .io_result(x569_1_io_result)
  );
  x525 x570_1 ( // @[Math.scala 262:24:@62647.4]
    .clock(x570_1_clock),
    .io_a(x570_1_io_a),
    .io_b(x570_1_io_b),
    .io_flow(x570_1_io_flow),
    .io_result(x570_1_io_result)
  );
  x534_x7 x571_x7_1 ( // @[Math.scala 150:24:@62657.4]
    .clock(x571_x7_1_clock),
    .reset(x571_x7_1_reset),
    .io_a(x571_x7_1_io_a),
    .io_b(x571_x7_1_io_b),
    .io_flow(x571_x7_1_io_flow),
    .io_result(x571_x7_1_io_result)
  );
  x534_x7 x572_x8_1 ( // @[Math.scala 150:24:@62667.4]
    .clock(x572_x8_1_clock),
    .reset(x572_x8_1_reset),
    .io_a(x572_x8_1_io_a),
    .io_b(x572_x8_1_io_b),
    .io_flow(x572_x8_1_io_flow),
    .io_result(x572_x8_1_io_result)
  );
  x534_x7 x573_x7_1 ( // @[Math.scala 150:24:@62677.4]
    .clock(x573_x7_1_clock),
    .reset(x573_x7_1_reset),
    .io_a(x573_x7_1_io_a),
    .io_b(x573_x7_1_io_b),
    .io_flow(x573_x7_1_io_flow),
    .io_result(x573_x7_1_io_result)
  );
  x534_x7 x574_x8_1 ( // @[Math.scala 150:24:@62687.4]
    .clock(x574_x8_1_clock),
    .reset(x574_x8_1_reset),
    .io_a(x574_x8_1_io_a),
    .io_b(x574_x8_1_io_b),
    .io_flow(x574_x8_1_io_flow),
    .io_result(x574_x8_1_io_result)
  );
  x534_x7 x575_x7_1 ( // @[Math.scala 150:24:@62697.4]
    .clock(x575_x7_1_clock),
    .reset(x575_x7_1_reset),
    .io_a(x575_x7_1_io_a),
    .io_b(x575_x7_1_io_b),
    .io_flow(x575_x7_1_io_flow),
    .io_result(x575_x7_1_io_result)
  );
  x534_x7 x576_x8_1 ( // @[Math.scala 150:24:@62707.4]
    .clock(x576_x8_1_clock),
    .reset(x576_x8_1_reset),
    .io_a(x576_x8_1_io_a),
    .io_b(x576_x8_1_io_b),
    .io_flow(x576_x8_1_io_flow),
    .io_result(x576_x8_1_io_result)
  );
  x534_x7 x577_x7_1 ( // @[Math.scala 150:24:@62717.4]
    .clock(x577_x7_1_clock),
    .reset(x577_x7_1_reset),
    .io_a(x577_x7_1_io_a),
    .io_b(x577_x7_1_io_b),
    .io_flow(x577_x7_1_io_flow),
    .io_result(x577_x7_1_io_result)
  );
  RetimeWrapper_443 RetimeWrapper_106 ( // @[package.scala 93:22:@62727.4]
    .clock(RetimeWrapper_106_clock),
    .reset(RetimeWrapper_106_reset),
    .io_flow(RetimeWrapper_106_io_flow),
    .io_in(RetimeWrapper_106_io_in),
    .io_out(RetimeWrapper_106_io_out)
  );
  x534_x7 x578_sum_1 ( // @[Math.scala 150:24:@62736.4]
    .clock(x578_sum_1_clock),
    .reset(x578_sum_1_reset),
    .io_a(x578_sum_1_io_a),
    .io_b(x578_sum_1_io_b),
    .io_flow(x578_sum_1_io_flow),
    .io_result(x578_sum_1_io_result)
  );
  x542 x579_1 ( // @[Math.scala 720:24:@62746.4]
    .io_b(x579_1_io_b),
    .io_result(x579_1_io_result)
  );
  x543_mul x580_mul_1 ( // @[Math.scala 262:24:@62757.4]
    .clock(x580_mul_1_clock),
    .io_a(x580_mul_1_io_a),
    .io_b(x580_mul_1_io_b),
    .io_flow(x580_mul_1_io_flow),
    .io_result(x580_mul_1_io_result)
  );
  x544 x581_1 ( // @[Math.scala 720:24:@62767.4]
    .io_b(x581_1_io_b),
    .io_result(x581_1_io_result)
  );
  x525 x582_1 ( // @[Math.scala 262:24:@62778.4]
    .clock(x582_1_clock),
    .io_a(x582_1_io_a),
    .io_b(x582_1_io_b),
    .io_flow(x582_1_io_flow),
    .io_result(x582_1_io_result)
  );
  x525 x583_1 ( // @[Math.scala 262:24:@62790.4]
    .clock(x583_1_clock),
    .io_a(x583_1_io_a),
    .io_b(x583_1_io_b),
    .io_flow(x583_1_io_flow),
    .io_result(x583_1_io_result)
  );
  x525 x584_1 ( // @[Math.scala 262:24:@62802.4]
    .clock(x584_1_clock),
    .io_a(x584_1_io_a),
    .io_b(x584_1_io_b),
    .io_flow(x584_1_io_flow),
    .io_result(x584_1_io_result)
  );
  x525 x585_1 ( // @[Math.scala 262:24:@62814.4]
    .clock(x585_1_clock),
    .io_a(x585_1_io_a),
    .io_b(x585_1_io_b),
    .io_flow(x585_1_io_flow),
    .io_result(x585_1_io_result)
  );
  x525 x586_1 ( // @[Math.scala 262:24:@62826.4]
    .clock(x586_1_clock),
    .io_a(x586_1_io_a),
    .io_b(x586_1_io_b),
    .io_flow(x586_1_io_flow),
    .io_result(x586_1_io_result)
  );
  x525 x587_1 ( // @[Math.scala 262:24:@62838.4]
    .clock(x587_1_clock),
    .io_a(x587_1_io_a),
    .io_b(x587_1_io_b),
    .io_flow(x587_1_io_flow),
    .io_result(x587_1_io_result)
  );
  x534_x7 x588_x7_1 ( // @[Math.scala 150:24:@62848.4]
    .clock(x588_x7_1_clock),
    .reset(x588_x7_1_reset),
    .io_a(x588_x7_1_io_a),
    .io_b(x588_x7_1_io_b),
    .io_flow(x588_x7_1_io_flow),
    .io_result(x588_x7_1_io_result)
  );
  x534_x7 x589_x8_1 ( // @[Math.scala 150:24:@62858.4]
    .clock(x589_x8_1_clock),
    .reset(x589_x8_1_reset),
    .io_a(x589_x8_1_io_a),
    .io_b(x589_x8_1_io_b),
    .io_flow(x589_x8_1_io_flow),
    .io_result(x589_x8_1_io_result)
  );
  x534_x7 x590_x7_1 ( // @[Math.scala 150:24:@62868.4]
    .clock(x590_x7_1_clock),
    .reset(x590_x7_1_reset),
    .io_a(x590_x7_1_io_a),
    .io_b(x590_x7_1_io_b),
    .io_flow(x590_x7_1_io_flow),
    .io_result(x590_x7_1_io_result)
  );
  x534_x7 x591_x8_1 ( // @[Math.scala 150:24:@62878.4]
    .clock(x591_x8_1_clock),
    .reset(x591_x8_1_reset),
    .io_a(x591_x8_1_io_a),
    .io_b(x591_x8_1_io_b),
    .io_flow(x591_x8_1_io_flow),
    .io_result(x591_x8_1_io_result)
  );
  x534_x7 x592_x7_1 ( // @[Math.scala 150:24:@62888.4]
    .clock(x592_x7_1_clock),
    .reset(x592_x7_1_reset),
    .io_a(x592_x7_1_io_a),
    .io_b(x592_x7_1_io_b),
    .io_flow(x592_x7_1_io_flow),
    .io_result(x592_x7_1_io_result)
  );
  x534_x7 x593_x8_1 ( // @[Math.scala 150:24:@62898.4]
    .clock(x593_x8_1_clock),
    .reset(x593_x8_1_reset),
    .io_a(x593_x8_1_io_a),
    .io_b(x593_x8_1_io_b),
    .io_flow(x593_x8_1_io_flow),
    .io_result(x593_x8_1_io_result)
  );
  x534_x7 x594_x7_1 ( // @[Math.scala 150:24:@62908.4]
    .clock(x594_x7_1_clock),
    .reset(x594_x7_1_reset),
    .io_a(x594_x7_1_io_a),
    .io_b(x594_x7_1_io_b),
    .io_flow(x594_x7_1_io_flow),
    .io_result(x594_x7_1_io_result)
  );
  RetimeWrapper_443 RetimeWrapper_107 ( // @[package.scala 93:22:@62918.4]
    .clock(RetimeWrapper_107_clock),
    .reset(RetimeWrapper_107_reset),
    .io_flow(RetimeWrapper_107_io_flow),
    .io_in(RetimeWrapper_107_io_in),
    .io_out(RetimeWrapper_107_io_out)
  );
  x534_x7 x595_sum_1 ( // @[Math.scala 150:24:@62927.4]
    .clock(x595_sum_1_clock),
    .reset(x595_sum_1_reset),
    .io_a(x595_sum_1_io_a),
    .io_b(x595_sum_1_io_b),
    .io_flow(x595_sum_1_io_flow),
    .io_result(x595_sum_1_io_result)
  );
  x542 x596_1 ( // @[Math.scala 720:24:@62939.4]
    .io_b(x596_1_io_b),
    .io_result(x596_1_io_result)
  );
  x543_mul x597_mul_1 ( // @[Math.scala 262:24:@62950.4]
    .clock(x597_mul_1_clock),
    .io_a(x597_mul_1_io_a),
    .io_b(x597_mul_1_io_b),
    .io_flow(x597_mul_1_io_flow),
    .io_result(x597_mul_1_io_result)
  );
  x544 x598_1 ( // @[Math.scala 720:24:@62960.4]
    .io_b(x598_1_io_b),
    .io_result(x598_1_io_result)
  );
  RetimeWrapper_604 RetimeWrapper_108 ( // @[package.scala 93:22:@62969.4]
    .clock(RetimeWrapper_108_clock),
    .reset(RetimeWrapper_108_reset),
    .io_flow(RetimeWrapper_108_io_flow),
    .io_in(RetimeWrapper_108_io_in),
    .io_out(RetimeWrapper_108_io_out)
  );
  RetimeWrapper_605 RetimeWrapper_109 ( // @[package.scala 93:22:@62978.4]
    .clock(RetimeWrapper_109_clock),
    .reset(RetimeWrapper_109_reset),
    .io_flow(RetimeWrapper_109_io_flow),
    .io_in(RetimeWrapper_109_io_in),
    .io_out(RetimeWrapper_109_io_out)
  );
  RetimeWrapper_604 RetimeWrapper_110 ( // @[package.scala 93:22:@62987.4]
    .clock(RetimeWrapper_110_clock),
    .reset(RetimeWrapper_110_reset),
    .io_flow(RetimeWrapper_110_io_flow),
    .io_in(RetimeWrapper_110_io_in),
    .io_out(RetimeWrapper_110_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_111 ( // @[package.scala 93:22:@62996.4]
    .clock(RetimeWrapper_111_clock),
    .reset(RetimeWrapper_111_reset),
    .io_flow(RetimeWrapper_111_io_flow),
    .io_in(RetimeWrapper_111_io_in),
    .io_out(RetimeWrapper_111_io_out)
  );
  RetimeWrapper_498 RetimeWrapper_112 ( // @[package.scala 93:22:@63005.4]
    .clock(RetimeWrapper_112_clock),
    .reset(RetimeWrapper_112_reset),
    .io_flow(RetimeWrapper_112_io_flow),
    .io_in(RetimeWrapper_112_io_in),
    .io_out(RetimeWrapper_112_io_out)
  );
  RetimeWrapper_609 RetimeWrapper_113 ( // @[package.scala 93:22:@63014.4]
    .clock(RetimeWrapper_113_clock),
    .reset(RetimeWrapper_113_reset),
    .io_flow(RetimeWrapper_113_io_flow),
    .io_in(RetimeWrapper_113_io_in),
    .io_out(RetimeWrapper_113_io_out)
  );
  RetimeWrapper_604 RetimeWrapper_114 ( // @[package.scala 93:22:@63025.4]
    .clock(RetimeWrapper_114_clock),
    .reset(RetimeWrapper_114_reset),
    .io_flow(RetimeWrapper_114_io_flow),
    .io_in(RetimeWrapper_114_io_in),
    .io_out(RetimeWrapper_114_io_out)
  );
  RetimeWrapper_611 RetimeWrapper_115 ( // @[package.scala 93:22:@63046.4]
    .clock(RetimeWrapper_115_clock),
    .reset(RetimeWrapper_115_reset),
    .io_flow(RetimeWrapper_115_io_flow),
    .io_in(RetimeWrapper_115_io_in),
    .io_out(RetimeWrapper_115_io_out)
  );
  RetimeWrapper_612 RetimeWrapper_116 ( // @[package.scala 93:22:@63055.4]
    .clock(RetimeWrapper_116_clock),
    .reset(RetimeWrapper_116_reset),
    .io_flow(RetimeWrapper_116_io_flow),
    .io_in(RetimeWrapper_116_io_in),
    .io_out(RetimeWrapper_116_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_117 ( // @[package.scala 93:22:@63064.4]
    .clock(RetimeWrapper_117_clock),
    .reset(RetimeWrapper_117_reset),
    .io_flow(RetimeWrapper_117_io_flow),
    .io_in(RetimeWrapper_117_io_in),
    .io_out(RetimeWrapper_117_io_out)
  );
  RetimeWrapper_604 RetimeWrapper_118 ( // @[package.scala 93:22:@63075.4]
    .clock(RetimeWrapper_118_clock),
    .reset(RetimeWrapper_118_reset),
    .io_flow(RetimeWrapper_118_io_flow),
    .io_in(RetimeWrapper_118_io_in),
    .io_out(RetimeWrapper_118_io_out)
  );
  RetimeWrapper_611 RetimeWrapper_119 ( // @[package.scala 93:22:@63096.4]
    .clock(RetimeWrapper_119_clock),
    .reset(RetimeWrapper_119_reset),
    .io_flow(RetimeWrapper_119_io_flow),
    .io_in(RetimeWrapper_119_io_in),
    .io_out(RetimeWrapper_119_io_out)
  );
  RetimeWrapper_612 RetimeWrapper_120 ( // @[package.scala 93:22:@63105.4]
    .clock(RetimeWrapper_120_clock),
    .reset(RetimeWrapper_120_reset),
    .io_flow(RetimeWrapper_120_io_flow),
    .io_in(RetimeWrapper_120_io_in),
    .io_out(RetimeWrapper_120_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_121 ( // @[package.scala 93:22:@63114.4]
    .clock(RetimeWrapper_121_clock),
    .reset(RetimeWrapper_121_reset),
    .io_flow(RetimeWrapper_121_io_flow),
    .io_in(RetimeWrapper_121_io_in),
    .io_out(RetimeWrapper_121_io_out)
  );
  RetimeWrapper_604 RetimeWrapper_122 ( // @[package.scala 93:22:@63125.4]
    .clock(RetimeWrapper_122_clock),
    .reset(RetimeWrapper_122_reset),
    .io_flow(RetimeWrapper_122_io_flow),
    .io_in(RetimeWrapper_122_io_in),
    .io_out(RetimeWrapper_122_io_out)
  );
  RetimeWrapper_612 RetimeWrapper_123 ( // @[package.scala 93:22:@63146.4]
    .clock(RetimeWrapper_123_clock),
    .reset(RetimeWrapper_123_reset),
    .io_flow(RetimeWrapper_123_io_flow),
    .io_in(RetimeWrapper_123_io_in),
    .io_out(RetimeWrapper_123_io_out)
  );
  RetimeWrapper_611 RetimeWrapper_124 ( // @[package.scala 93:22:@63155.4]
    .clock(RetimeWrapper_124_clock),
    .reset(RetimeWrapper_124_reset),
    .io_flow(RetimeWrapper_124_io_flow),
    .io_in(RetimeWrapper_124_io_in),
    .io_out(RetimeWrapper_124_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_125 ( // @[package.scala 93:22:@63164.4]
    .clock(RetimeWrapper_125_clock),
    .reset(RetimeWrapper_125_reset),
    .io_flow(RetimeWrapper_125_io_flow),
    .io_in(RetimeWrapper_125_io_in),
    .io_out(RetimeWrapper_125_io_out)
  );
  RetimeWrapper_604 RetimeWrapper_126 ( // @[package.scala 93:22:@63175.4]
    .clock(RetimeWrapper_126_clock),
    .reset(RetimeWrapper_126_reset),
    .io_flow(RetimeWrapper_126_io_flow),
    .io_in(RetimeWrapper_126_io_in),
    .io_out(RetimeWrapper_126_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_127 ( // @[package.scala 93:22:@63196.4]
    .clock(RetimeWrapper_127_clock),
    .reset(RetimeWrapper_127_reset),
    .io_flow(RetimeWrapper_127_io_flow),
    .io_in(RetimeWrapper_127_io_in),
    .io_out(RetimeWrapper_127_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_128 ( // @[package.scala 93:22:@63205.4]
    .clock(RetimeWrapper_128_clock),
    .reset(RetimeWrapper_128_reset),
    .io_flow(RetimeWrapper_128_io_flow),
    .io_in(RetimeWrapper_128_io_in),
    .io_out(RetimeWrapper_128_io_out)
  );
  RetimeWrapper_498 RetimeWrapper_129 ( // @[package.scala 93:22:@63214.4]
    .clock(RetimeWrapper_129_clock),
    .reset(RetimeWrapper_129_reset),
    .io_flow(RetimeWrapper_129_io_flow),
    .io_in(RetimeWrapper_129_io_in),
    .io_out(RetimeWrapper_129_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_130 ( // @[package.scala 93:22:@63223.4]
    .clock(RetimeWrapper_130_clock),
    .reset(RetimeWrapper_130_reset),
    .io_flow(RetimeWrapper_130_io_flow),
    .io_in(RetimeWrapper_130_io_in),
    .io_out(RetimeWrapper_130_io_out)
  );
  RetimeWrapper_627 RetimeWrapper_131 ( // @[package.scala 93:22:@63232.4]
    .clock(RetimeWrapper_131_clock),
    .reset(RetimeWrapper_131_reset),
    .io_flow(RetimeWrapper_131_io_flow),
    .io_in(RetimeWrapper_131_io_in),
    .io_out(RetimeWrapper_131_io_out)
  );
  RetimeWrapper_605 RetimeWrapper_132 ( // @[package.scala 93:22:@63241.4]
    .clock(RetimeWrapper_132_clock),
    .reset(RetimeWrapper_132_reset),
    .io_flow(RetimeWrapper_132_io_flow),
    .io_in(RetimeWrapper_132_io_in),
    .io_out(RetimeWrapper_132_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_133 ( // @[package.scala 93:22:@63253.4]
    .clock(RetimeWrapper_133_clock),
    .reset(RetimeWrapper_133_reset),
    .io_flow(RetimeWrapper_133_io_flow),
    .io_in(RetimeWrapper_133_io_in),
    .io_out(RetimeWrapper_133_io_out)
  );
  RetimeWrapper_605 RetimeWrapper_134 ( // @[package.scala 93:22:@63274.4]
    .clock(RetimeWrapper_134_clock),
    .reset(RetimeWrapper_134_reset),
    .io_flow(RetimeWrapper_134_io_flow),
    .io_in(RetimeWrapper_134_io_in),
    .io_out(RetimeWrapper_134_io_out)
  );
  RetimeWrapper_498 RetimeWrapper_135 ( // @[package.scala 93:22:@63283.4]
    .clock(RetimeWrapper_135_clock),
    .reset(RetimeWrapper_135_reset),
    .io_flow(RetimeWrapper_135_io_flow),
    .io_in(RetimeWrapper_135_io_in),
    .io_out(RetimeWrapper_135_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_136 ( // @[package.scala 93:22:@63292.4]
    .clock(RetimeWrapper_136_clock),
    .reset(RetimeWrapper_136_reset),
    .io_flow(RetimeWrapper_136_io_flow),
    .io_in(RetimeWrapper_136_io_in),
    .io_out(RetimeWrapper_136_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_137 ( // @[package.scala 93:22:@63304.4]
    .clock(RetimeWrapper_137_clock),
    .reset(RetimeWrapper_137_reset),
    .io_flow(RetimeWrapper_137_io_flow),
    .io_in(RetimeWrapper_137_io_in),
    .io_out(RetimeWrapper_137_io_out)
  );
  RetimeWrapper_605 RetimeWrapper_138 ( // @[package.scala 93:22:@63325.4]
    .clock(RetimeWrapper_138_clock),
    .reset(RetimeWrapper_138_reset),
    .io_flow(RetimeWrapper_138_io_flow),
    .io_in(RetimeWrapper_138_io_in),
    .io_out(RetimeWrapper_138_io_out)
  );
  RetimeWrapper_498 RetimeWrapper_139 ( // @[package.scala 93:22:@63334.4]
    .clock(RetimeWrapper_139_clock),
    .reset(RetimeWrapper_139_reset),
    .io_flow(RetimeWrapper_139_io_flow),
    .io_in(RetimeWrapper_139_io_in),
    .io_out(RetimeWrapper_139_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_140 ( // @[package.scala 93:22:@63343.4]
    .clock(RetimeWrapper_140_clock),
    .reset(RetimeWrapper_140_reset),
    .io_flow(RetimeWrapper_140_io_flow),
    .io_in(RetimeWrapper_140_io_in),
    .io_out(RetimeWrapper_140_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_141 ( // @[package.scala 93:22:@63355.4]
    .clock(RetimeWrapper_141_clock),
    .reset(RetimeWrapper_141_reset),
    .io_flow(RetimeWrapper_141_io_flow),
    .io_in(RetimeWrapper_141_io_in),
    .io_out(RetimeWrapper_141_io_out)
  );
  RetimeWrapper_638 RetimeWrapper_142 ( // @[package.scala 93:22:@63376.4]
    .clock(RetimeWrapper_142_clock),
    .reset(RetimeWrapper_142_reset),
    .io_flow(RetimeWrapper_142_io_flow),
    .io_in(RetimeWrapper_142_io_in),
    .io_out(RetimeWrapper_142_io_out)
  );
  RetimeWrapper_639 RetimeWrapper_143 ( // @[package.scala 93:22:@63385.4]
    .clock(RetimeWrapper_143_clock),
    .reset(RetimeWrapper_143_reset),
    .io_flow(RetimeWrapper_143_io_flow),
    .io_in(RetimeWrapper_143_io_in),
    .io_out(RetimeWrapper_143_io_out)
  );
  RetimeWrapper_640 RetimeWrapper_144 ( // @[package.scala 93:22:@63394.4]
    .clock(RetimeWrapper_144_clock),
    .reset(RetimeWrapper_144_reset),
    .io_flow(RetimeWrapper_144_io_flow),
    .io_in(RetimeWrapper_144_io_in),
    .io_out(RetimeWrapper_144_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_145 ( // @[package.scala 93:22:@63406.4]
    .clock(RetimeWrapper_145_clock),
    .reset(RetimeWrapper_145_reset),
    .io_flow(RetimeWrapper_145_io_flow),
    .io_in(RetimeWrapper_145_io_in),
    .io_out(RetimeWrapper_145_io_out)
  );
  RetimeWrapper_642 RetimeWrapper_146 ( // @[package.scala 93:22:@63427.4]
    .clock(RetimeWrapper_146_clock),
    .reset(RetimeWrapper_146_reset),
    .io_flow(RetimeWrapper_146_io_flow),
    .io_in(RetimeWrapper_146_io_in),
    .io_out(RetimeWrapper_146_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_147 ( // @[package.scala 93:22:@63436.4]
    .clock(RetimeWrapper_147_clock),
    .reset(RetimeWrapper_147_reset),
    .io_flow(RetimeWrapper_147_io_flow),
    .io_in(RetimeWrapper_147_io_in),
    .io_out(RetimeWrapper_147_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_148 ( // @[package.scala 93:22:@63445.4]
    .clock(RetimeWrapper_148_clock),
    .reset(RetimeWrapper_148_reset),
    .io_flow(RetimeWrapper_148_io_flow),
    .io_in(RetimeWrapper_148_io_in),
    .io_out(RetimeWrapper_148_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_149 ( // @[package.scala 93:22:@63457.4]
    .clock(RetimeWrapper_149_clock),
    .reset(RetimeWrapper_149_reset),
    .io_flow(RetimeWrapper_149_io_flow),
    .io_in(RetimeWrapper_149_io_in),
    .io_out(RetimeWrapper_149_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_150 ( // @[package.scala 93:22:@63478.4]
    .clock(RetimeWrapper_150_clock),
    .reset(RetimeWrapper_150_reset),
    .io_flow(RetimeWrapper_150_io_flow),
    .io_in(RetimeWrapper_150_io_in),
    .io_out(RetimeWrapper_150_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_151 ( // @[package.scala 93:22:@63487.4]
    .clock(RetimeWrapper_151_clock),
    .reset(RetimeWrapper_151_reset),
    .io_flow(RetimeWrapper_151_io_flow),
    .io_in(RetimeWrapper_151_io_in),
    .io_out(RetimeWrapper_151_io_out)
  );
  RetimeWrapper_648 RetimeWrapper_152 ( // @[package.scala 93:22:@63496.4]
    .clock(RetimeWrapper_152_clock),
    .reset(RetimeWrapper_152_reset),
    .io_flow(RetimeWrapper_152_io_flow),
    .io_in(RetimeWrapper_152_io_in),
    .io_out(RetimeWrapper_152_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_153 ( // @[package.scala 93:22:@63508.4]
    .clock(RetimeWrapper_153_clock),
    .reset(RetimeWrapper_153_reset),
    .io_flow(RetimeWrapper_153_io_flow),
    .io_in(RetimeWrapper_153_io_in),
    .io_out(RetimeWrapper_153_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_154 ( // @[package.scala 93:22:@63529.4]
    .clock(RetimeWrapper_154_clock),
    .reset(RetimeWrapper_154_reset),
    .io_flow(RetimeWrapper_154_io_flow),
    .io_in(RetimeWrapper_154_io_in),
    .io_out(RetimeWrapper_154_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_155 ( // @[package.scala 93:22:@63538.4]
    .clock(RetimeWrapper_155_clock),
    .reset(RetimeWrapper_155_reset),
    .io_flow(RetimeWrapper_155_io_flow),
    .io_in(RetimeWrapper_155_io_in),
    .io_out(RetimeWrapper_155_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_156 ( // @[package.scala 93:22:@63550.4]
    .clock(RetimeWrapper_156_clock),
    .reset(RetimeWrapper_156_reset),
    .io_flow(RetimeWrapper_156_io_flow),
    .io_in(RetimeWrapper_156_io_in),
    .io_out(RetimeWrapper_156_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_157 ( // @[package.scala 93:22:@63571.4]
    .clock(RetimeWrapper_157_clock),
    .reset(RetimeWrapper_157_reset),
    .io_flow(RetimeWrapper_157_io_flow),
    .io_in(RetimeWrapper_157_io_in),
    .io_out(RetimeWrapper_157_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_158 ( // @[package.scala 93:22:@63580.4]
    .clock(RetimeWrapper_158_clock),
    .reset(RetimeWrapper_158_reset),
    .io_flow(RetimeWrapper_158_io_flow),
    .io_in(RetimeWrapper_158_io_in),
    .io_out(RetimeWrapper_158_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_159 ( // @[package.scala 93:22:@63592.4]
    .clock(RetimeWrapper_159_clock),
    .reset(RetimeWrapper_159_reset),
    .io_flow(RetimeWrapper_159_io_flow),
    .io_in(RetimeWrapper_159_io_in),
    .io_out(RetimeWrapper_159_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_160 ( // @[package.scala 93:22:@63613.4]
    .clock(RetimeWrapper_160_clock),
    .reset(RetimeWrapper_160_reset),
    .io_flow(RetimeWrapper_160_io_flow),
    .io_in(RetimeWrapper_160_io_in),
    .io_out(RetimeWrapper_160_io_out)
  );
  RetimeWrapper_657 RetimeWrapper_161 ( // @[package.scala 93:22:@63622.4]
    .clock(RetimeWrapper_161_clock),
    .reset(RetimeWrapper_161_reset),
    .io_flow(RetimeWrapper_161_io_flow),
    .io_in(RetimeWrapper_161_io_in),
    .io_out(RetimeWrapper_161_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_162 ( // @[package.scala 93:22:@63634.4]
    .clock(RetimeWrapper_162_clock),
    .reset(RetimeWrapper_162_reset),
    .io_flow(RetimeWrapper_162_io_flow),
    .io_in(RetimeWrapper_162_io_in),
    .io_out(RetimeWrapper_162_io_out)
  );
  RetimeWrapper_448 RetimeWrapper_163 ( // @[package.scala 93:22:@63655.4]
    .clock(RetimeWrapper_163_clock),
    .reset(RetimeWrapper_163_reset),
    .io_flow(RetimeWrapper_163_io_flow),
    .io_in(RetimeWrapper_163_io_in),
    .io_out(RetimeWrapper_163_io_out)
  );
  RetimeWrapper_624 RetimeWrapper_164 ( // @[package.scala 93:22:@63664.4]
    .clock(RetimeWrapper_164_clock),
    .reset(RetimeWrapper_164_reset),
    .io_flow(RetimeWrapper_164_io_flow),
    .io_in(RetimeWrapper_164_io_in),
    .io_out(RetimeWrapper_164_io_out)
  );
  RetimeWrapper_623 RetimeWrapper_165 ( // @[package.scala 93:22:@63676.4]
    .clock(RetimeWrapper_165_clock),
    .reset(RetimeWrapper_165_reset),
    .io_flow(RetimeWrapper_165_io_flow),
    .io_in(RetimeWrapper_165_io_in),
    .io_out(RetimeWrapper_165_io_out)
  );
  x525 x625_1 ( // @[Math.scala 262:24:@63701.4]
    .clock(x625_1_clock),
    .io_a(x625_1_io_a),
    .io_b(x625_1_io_b),
    .io_flow(x625_1_io_flow),
    .io_result(x625_1_io_result)
  );
  x525 x626_1 ( // @[Math.scala 262:24:@63713.4]
    .clock(x626_1_clock),
    .io_a(x626_1_io_a),
    .io_b(x626_1_io_b),
    .io_flow(x626_1_io_flow),
    .io_result(x626_1_io_result)
  );
  x525 x627_1 ( // @[Math.scala 262:24:@63725.4]
    .clock(x627_1_clock),
    .io_a(x627_1_io_a),
    .io_b(x627_1_io_b),
    .io_flow(x627_1_io_flow),
    .io_result(x627_1_io_result)
  );
  x525 x628_1 ( // @[Math.scala 262:24:@63737.4]
    .clock(x628_1_clock),
    .io_a(x628_1_io_a),
    .io_b(x628_1_io_b),
    .io_flow(x628_1_io_flow),
    .io_result(x628_1_io_result)
  );
  x534_x7 x629_x9_1 ( // @[Math.scala 150:24:@63747.4]
    .clock(x629_x9_1_clock),
    .reset(x629_x9_1_reset),
    .io_a(x629_x9_1_io_a),
    .io_b(x629_x9_1_io_b),
    .io_flow(x629_x9_1_io_flow),
    .io_result(x629_x9_1_io_result)
  );
  x534_x7 x630_x10_1 ( // @[Math.scala 150:24:@63757.4]
    .clock(x630_x10_1_clock),
    .reset(x630_x10_1_reset),
    .io_a(x630_x10_1_io_a),
    .io_b(x630_x10_1_io_b),
    .io_flow(x630_x10_1_io_flow),
    .io_result(x630_x10_1_io_result)
  );
  x534_x7 x631_sum_1 ( // @[Math.scala 150:24:@63767.4]
    .clock(x631_sum_1_clock),
    .reset(x631_sum_1_reset),
    .io_a(x631_sum_1_io_a),
    .io_b(x631_sum_1_io_b),
    .io_flow(x631_sum_1_io_flow),
    .io_result(x631_sum_1_io_result)
  );
  x542 x632_1 ( // @[Math.scala 720:24:@63777.4]
    .io_b(x632_1_io_b),
    .io_result(x632_1_io_result)
  );
  x543_mul x633_mul_1 ( // @[Math.scala 262:24:@63788.4]
    .clock(x633_mul_1_clock),
    .io_a(x633_mul_1_io_a),
    .io_b(x633_mul_1_io_b),
    .io_flow(x633_mul_1_io_flow),
    .io_result(x633_mul_1_io_result)
  );
  x544 x634_1 ( // @[Math.scala 720:24:@63798.4]
    .io_b(x634_1_io_b),
    .io_result(x634_1_io_result)
  );
  x525 x635_1 ( // @[Math.scala 262:24:@63809.4]
    .clock(x635_1_clock),
    .io_a(x635_1_io_a),
    .io_b(x635_1_io_b),
    .io_flow(x635_1_io_flow),
    .io_result(x635_1_io_result)
  );
  x525 x636_1 ( // @[Math.scala 262:24:@63821.4]
    .clock(x636_1_clock),
    .io_a(x636_1_io_a),
    .io_b(x636_1_io_b),
    .io_flow(x636_1_io_flow),
    .io_result(x636_1_io_result)
  );
  x525 x637_1 ( // @[Math.scala 262:24:@63833.4]
    .clock(x637_1_clock),
    .io_a(x637_1_io_a),
    .io_b(x637_1_io_b),
    .io_flow(x637_1_io_flow),
    .io_result(x637_1_io_result)
  );
  x525 x638_1 ( // @[Math.scala 262:24:@63845.4]
    .clock(x638_1_clock),
    .io_a(x638_1_io_a),
    .io_b(x638_1_io_b),
    .io_flow(x638_1_io_flow),
    .io_result(x638_1_io_result)
  );
  x534_x7 x639_x9_1 ( // @[Math.scala 150:24:@63855.4]
    .clock(x639_x9_1_clock),
    .reset(x639_x9_1_reset),
    .io_a(x639_x9_1_io_a),
    .io_b(x639_x9_1_io_b),
    .io_flow(x639_x9_1_io_flow),
    .io_result(x639_x9_1_io_result)
  );
  x534_x7 x640_x10_1 ( // @[Math.scala 150:24:@63865.4]
    .clock(x640_x10_1_clock),
    .reset(x640_x10_1_reset),
    .io_a(x640_x10_1_io_a),
    .io_b(x640_x10_1_io_b),
    .io_flow(x640_x10_1_io_flow),
    .io_result(x640_x10_1_io_result)
  );
  x534_x7 x641_sum_1 ( // @[Math.scala 150:24:@63875.4]
    .clock(x641_sum_1_clock),
    .reset(x641_sum_1_reset),
    .io_a(x641_sum_1_io_a),
    .io_b(x641_sum_1_io_b),
    .io_flow(x641_sum_1_io_flow),
    .io_result(x641_sum_1_io_result)
  );
  x542 x642_1 ( // @[Math.scala 720:24:@63885.4]
    .io_b(x642_1_io_b),
    .io_result(x642_1_io_result)
  );
  x543_mul x643_mul_1 ( // @[Math.scala 262:24:@63896.4]
    .clock(x643_mul_1_clock),
    .io_a(x643_mul_1_io_a),
    .io_b(x643_mul_1_io_b),
    .io_flow(x643_mul_1_io_flow),
    .io_result(x643_mul_1_io_result)
  );
  x544 x644_1 ( // @[Math.scala 720:24:@63906.4]
    .io_b(x644_1_io_b),
    .io_result(x644_1_io_result)
  );
  x525 x645_1 ( // @[Math.scala 262:24:@63917.4]
    .clock(x645_1_clock),
    .io_a(x645_1_io_a),
    .io_b(x645_1_io_b),
    .io_flow(x645_1_io_flow),
    .io_result(x645_1_io_result)
  );
  x525 x646_1 ( // @[Math.scala 262:24:@63929.4]
    .clock(x646_1_clock),
    .io_a(x646_1_io_a),
    .io_b(x646_1_io_b),
    .io_flow(x646_1_io_flow),
    .io_result(x646_1_io_result)
  );
  x525 x647_1 ( // @[Math.scala 262:24:@63941.4]
    .clock(x647_1_clock),
    .io_a(x647_1_io_a),
    .io_b(x647_1_io_b),
    .io_flow(x647_1_io_flow),
    .io_result(x647_1_io_result)
  );
  x525 x648_1 ( // @[Math.scala 262:24:@63953.4]
    .clock(x648_1_clock),
    .io_a(x648_1_io_a),
    .io_b(x648_1_io_b),
    .io_flow(x648_1_io_flow),
    .io_result(x648_1_io_result)
  );
  x534_x7 x649_x9_1 ( // @[Math.scala 150:24:@63963.4]
    .clock(x649_x9_1_clock),
    .reset(x649_x9_1_reset),
    .io_a(x649_x9_1_io_a),
    .io_b(x649_x9_1_io_b),
    .io_flow(x649_x9_1_io_flow),
    .io_result(x649_x9_1_io_result)
  );
  x534_x7 x650_x10_1 ( // @[Math.scala 150:24:@63975.4]
    .clock(x650_x10_1_clock),
    .reset(x650_x10_1_reset),
    .io_a(x650_x10_1_io_a),
    .io_b(x650_x10_1_io_b),
    .io_flow(x650_x10_1_io_flow),
    .io_result(x650_x10_1_io_result)
  );
  x534_x7 x651_sum_1 ( // @[Math.scala 150:24:@63985.4]
    .clock(x651_sum_1_clock),
    .reset(x651_sum_1_reset),
    .io_a(x651_sum_1_io_a),
    .io_b(x651_sum_1_io_b),
    .io_flow(x651_sum_1_io_flow),
    .io_result(x651_sum_1_io_result)
  );
  x542 x652_1 ( // @[Math.scala 720:24:@63995.4]
    .io_b(x652_1_io_b),
    .io_result(x652_1_io_result)
  );
  x543_mul x653_mul_1 ( // @[Math.scala 262:24:@64006.4]
    .clock(x653_mul_1_clock),
    .io_a(x653_mul_1_io_a),
    .io_b(x653_mul_1_io_b),
    .io_flow(x653_mul_1_io_flow),
    .io_result(x653_mul_1_io_result)
  );
  x544 x654_1 ( // @[Math.scala 720:24:@64016.4]
    .io_b(x654_1_io_b),
    .io_result(x654_1_io_result)
  );
  x525 x655_1 ( // @[Math.scala 262:24:@64027.4]
    .clock(x655_1_clock),
    .io_a(x655_1_io_a),
    .io_b(x655_1_io_b),
    .io_flow(x655_1_io_flow),
    .io_result(x655_1_io_result)
  );
  x525 x656_1 ( // @[Math.scala 262:24:@64039.4]
    .clock(x656_1_clock),
    .io_a(x656_1_io_a),
    .io_b(x656_1_io_b),
    .io_flow(x656_1_io_flow),
    .io_result(x656_1_io_result)
  );
  x525 x657_1 ( // @[Math.scala 262:24:@64051.4]
    .clock(x657_1_clock),
    .io_a(x657_1_io_a),
    .io_b(x657_1_io_b),
    .io_flow(x657_1_io_flow),
    .io_result(x657_1_io_result)
  );
  x525 x658_1 ( // @[Math.scala 262:24:@64063.4]
    .clock(x658_1_clock),
    .io_a(x658_1_io_a),
    .io_b(x658_1_io_b),
    .io_flow(x658_1_io_flow),
    .io_result(x658_1_io_result)
  );
  x534_x7 x659_x9_1 ( // @[Math.scala 150:24:@64073.4]
    .clock(x659_x9_1_clock),
    .reset(x659_x9_1_reset),
    .io_a(x659_x9_1_io_a),
    .io_b(x659_x9_1_io_b),
    .io_flow(x659_x9_1_io_flow),
    .io_result(x659_x9_1_io_result)
  );
  x534_x7 x660_x10_1 ( // @[Math.scala 150:24:@64083.4]
    .clock(x660_x10_1_clock),
    .reset(x660_x10_1_reset),
    .io_a(x660_x10_1_io_a),
    .io_b(x660_x10_1_io_b),
    .io_flow(x660_x10_1_io_flow),
    .io_result(x660_x10_1_io_result)
  );
  x534_x7 x661_sum_1 ( // @[Math.scala 150:24:@64093.4]
    .clock(x661_sum_1_clock),
    .reset(x661_sum_1_reset),
    .io_a(x661_sum_1_io_a),
    .io_b(x661_sum_1_io_b),
    .io_flow(x661_sum_1_io_flow),
    .io_result(x661_sum_1_io_result)
  );
  x542 x662_1 ( // @[Math.scala 720:24:@64103.4]
    .io_b(x662_1_io_b),
    .io_result(x662_1_io_result)
  );
  x543_mul x663_mul_1 ( // @[Math.scala 262:24:@64114.4]
    .clock(x663_mul_1_clock),
    .io_a(x663_mul_1_io_a),
    .io_b(x663_mul_1_io_b),
    .io_flow(x663_mul_1_io_flow),
    .io_result(x663_mul_1_io_result)
  );
  x544 x664_1 ( // @[Math.scala 720:24:@64124.4]
    .io_b(x664_1_io_b),
    .io_result(x664_1_io_result)
  );
  RetimeWrapper_674 RetimeWrapper_166 ( // @[package.scala 93:22:@64143.4]
    .clock(RetimeWrapper_166_clock),
    .reset(RetimeWrapper_166_reset),
    .io_flow(RetimeWrapper_166_io_flow),
    .io_in(RetimeWrapper_166_io_in),
    .io_out(RetimeWrapper_166_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_167 ( // @[package.scala 93:22:@64152.4]
    .clock(RetimeWrapper_167_clock),
    .reset(RetimeWrapper_167_reset),
    .io_flow(RetimeWrapper_167_io_flow),
    .io_in(RetimeWrapper_167_io_in),
    .io_out(RetimeWrapper_167_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_168 ( // @[package.scala 93:22:@64161.4]
    .clock(RetimeWrapper_168_clock),
    .reset(RetimeWrapper_168_reset),
    .io_flow(RetimeWrapper_168_io_flow),
    .io_in(RetimeWrapper_168_io_in),
    .io_out(RetimeWrapper_168_io_out)
  );
  RetimeWrapper_675 RetimeWrapper_169 ( // @[package.scala 93:22:@64170.4]
    .clock(RetimeWrapper_169_clock),
    .reset(RetimeWrapper_169_reset),
    .io_flow(RetimeWrapper_169_io_flow),
    .io_in(RetimeWrapper_169_io_in),
    .io_out(RetimeWrapper_169_io_out)
  );
  assign b379 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 62:18:@59847.4]
  assign b380 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 63:18:@59848.4]
  assign _T_205 = b379 & b380; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 67:30:@59850.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 67:37:@59851.4]
  assign _T_210 = io_in_x342_TID == 8'h0; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 69:76:@59856.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 69:62:@59857.4]
  assign _T_213 = io_in_x342_TDEST == 8'h0; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 69:101:@59858.4]
  assign x745_x381_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@59867.4 package.scala 96:25:@59868.4]
  assign b377_number = __io_result; // @[Math.scala 723:22:@59832.4 Math.scala 724:14:@59833.4]
  assign _T_248 = $signed(b377_number); // @[Math.scala 406:49:@60129.4]
  assign _T_250 = $signed(_T_248) & $signed(32'sh3); // @[Math.scala 406:56:@60131.4]
  assign _T_251 = $signed(_T_250); // @[Math.scala 406:56:@60132.4]
  assign x725_number = $unsigned(_T_251); // @[implicits.scala 133:21:@60133.4]
  assign _T_261 = $signed(x725_number); // @[Math.scala 406:49:@60142.4]
  assign _T_263 = $signed(_T_261) & $signed(32'sh3); // @[Math.scala 406:56:@60144.4]
  assign _T_264 = $signed(_T_263); // @[Math.scala 406:56:@60145.4]
  assign _T_275 = x725_number[31]; // @[FixedPoint.scala 50:25:@60163.4]
  assign _T_279 = _T_275 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@60165.4]
  assign _T_280 = x725_number[31:2]; // @[FixedPoint.scala 18:52:@60166.4]
  assign _T_286 = _T_280 == 30'h3fffffff; // @[Math.scala 451:55:@60168.4]
  assign _T_287 = x725_number[1:0]; // @[FixedPoint.scala 18:52:@60169.4]
  assign _T_293 = _T_287 != 2'h0; // @[Math.scala 451:110:@60171.4]
  assign _T_294 = _T_286 & _T_293; // @[Math.scala 451:94:@60172.4]
  assign _T_296 = {_T_279,_T_280}; // @[Cat.scala 30:58:@60174.4]
  assign x390_1_number = _T_294 ? 32'h0 : _T_296; // @[Math.scala 454:20:@60175.4]
  assign _GEN_0 = {{8'd0}, x390_1_number}; // @[Math.scala 461:32:@60180.4]
  assign _T_301 = _GEN_0 << 8; // @[Math.scala 461:32:@60180.4]
  assign _GEN_1 = {{6'd0}, x390_1_number}; // @[Math.scala 461:32:@60185.4]
  assign _T_304 = _GEN_1 << 6; // @[Math.scala 461:32:@60185.4]
  assign _T_340 = ~ io_sigsIn_break; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:101:@60283.4]
  assign _T_344 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@60291.4 package.scala 96:25:@60292.4]
  assign _T_346 = io_rr ? _T_344 : 1'h0; // @[implicits.scala 55:10:@60293.4]
  assign _T_347 = _T_340 & _T_346; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:118:@60294.4]
  assign _T_349 = _T_347 & _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:207:@60296.4]
  assign _T_350 = _T_349 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:226:@60297.4]
  assign x747_b379_D24 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@60235.4 package.scala 96:25:@60236.4]
  assign _T_351 = _T_350 & x747_b379_D24; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 118:252:@60298.4]
  assign x749_b380_D24 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@60253.4 package.scala 96:25:@60254.4]
  assign _T_395 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@60398.4 package.scala 96:25:@60399.4]
  assign _T_397 = io_rr ? _T_395 : 1'h0; // @[implicits.scala 55:10:@60400.4]
  assign _T_398 = _T_340 & _T_397; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 141:118:@60401.4]
  assign _T_400 = _T_398 & _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 141:207:@60403.4]
  assign _T_401 = _T_400 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 141:226:@60404.4]
  assign _T_402 = _T_401 & x747_b379_D24; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 141:252:@60405.4]
  assign _T_443 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@60496.4 package.scala 96:25:@60497.4]
  assign _T_445 = io_rr ? _T_443 : 1'h0; // @[implicits.scala 55:10:@60498.4]
  assign _T_446 = _T_340 & _T_445; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 162:118:@60499.4]
  assign _T_448 = _T_446 & _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 162:207:@60501.4]
  assign _T_449 = _T_448 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 162:226:@60502.4]
  assign _T_450 = _T_449 & x747_b379_D24; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 162:252:@60503.4]
  assign _T_491 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@60594.4 package.scala 96:25:@60595.4]
  assign _T_493 = io_rr ? _T_491 : 1'h0; // @[implicits.scala 55:10:@60596.4]
  assign _T_494 = _T_340 & _T_493; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 189:166:@60597.4]
  assign _T_496 = _T_494 & _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 189:255:@60599.4]
  assign _T_497 = _T_496 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 189:274:@60600.4]
  assign _T_498 = _T_497 & x747_b379_D24; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 189:300:@60601.4]
  assign x763_b377_D26_number = RetimeWrapper_22_io_out; // @[package.scala 96:25:@60615.4 package.scala 96:25:@60616.4]
  assign _T_510 = $signed(x763_b377_D26_number); // @[Math.scala 476:37:@60623.4]
  assign x764_x407_rdcol_D26_number = RetimeWrapper_24_io_out; // @[package.scala 96:25:@60640.4 package.scala 96:25:@60641.4]
  assign _T_523 = $signed(x764_x407_rdcol_D26_number); // @[Math.scala 476:37:@60646.4]
  assign x765_x414_D1 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@60663.4 package.scala 96:25:@60664.4]
  assign x415 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@60654.4 package.scala 96:25:@60655.4]
  assign x416 = x765_x414_D1 | x415; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 204:24:@60667.4]
  assign _T_564 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@60735.4 package.scala 96:25:@60736.4]
  assign _T_566 = io_rr ? _T_564 : 1'h0; // @[implicits.scala 55:10:@60737.4]
  assign _T_567 = _T_340 & _T_566; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 223:194:@60738.4]
  assign x767_x417_D20 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@60687.4 package.scala 96:25:@60688.4]
  assign _T_568 = _T_567 & x767_x417_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 223:283:@60739.4]
  assign x766_b379_D48 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@60678.4 package.scala 96:25:@60679.4]
  assign _T_569 = _T_568 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 223:291:@60740.4]
  assign x769_b380_D48 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@60705.4 package.scala 96:25:@60706.4]
  assign x772_x401_rdcol_D26_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@60756.4 package.scala 96:25:@60757.4]
  assign _T_580 = $signed(x772_x401_rdcol_D26_number); // @[Math.scala 476:37:@60762.4]
  assign x420 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@60770.4 package.scala 96:25:@60771.4]
  assign x421 = x765_x414_D1 | x420; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 231:24:@60774.4]
  assign _T_609 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@60815.4 package.scala 96:25:@60816.4]
  assign _T_611 = io_rr ? _T_609 : 1'h0; // @[implicits.scala 55:10:@60817.4]
  assign _T_612 = _T_340 & _T_611; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 244:194:@60818.4]
  assign x775_x422_D20 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@60803.4 package.scala 96:25:@60804.4]
  assign _T_613 = _T_612 & x775_x422_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 244:283:@60819.4]
  assign _T_614 = _T_613 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 244:291:@60820.4]
  assign x776_x395_rdcol_D26_number = RetimeWrapper_40_io_out; // @[package.scala 96:25:@60836.4 package.scala 96:25:@60837.4]
  assign _T_625 = $signed(x776_x395_rdcol_D26_number); // @[Math.scala 476:37:@60842.4]
  assign x425 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@60850.4 package.scala 96:25:@60851.4]
  assign x426 = x765_x414_D1 | x425; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 252:24:@60854.4]
  assign _T_654 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@60895.4 package.scala 96:25:@60896.4]
  assign _T_656 = io_rr ? _T_654 : 1'h0; // @[implicits.scala 55:10:@60897.4]
  assign _T_657 = _T_340 & _T_656; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 265:194:@60898.4]
  assign x779_x427_D20 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@60883.4 package.scala 96:25:@60884.4]
  assign _T_658 = _T_657 & x779_x427_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 265:283:@60899.4]
  assign _T_659 = _T_658 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 265:291:@60900.4]
  assign x780_b378_D26_number = RetimeWrapper_46_io_out; // @[package.scala 96:25:@60916.4 package.scala 96:25:@60917.4]
  assign _T_670 = $signed(x780_b378_D26_number); // @[Math.scala 476:37:@60922.4]
  assign x414 = RetimeWrapper_23_io_out; // @[package.scala 96:25:@60631.4 package.scala 96:25:@60632.4]
  assign x430 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@60930.4 package.scala 96:25:@60931.4]
  assign x431 = x414 | x430; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 273:24:@60934.4]
  assign _T_699 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@60975.4 package.scala 96:25:@60976.4]
  assign _T_701 = io_rr ? _T_699 : 1'h0; // @[implicits.scala 55:10:@60977.4]
  assign _T_702 = _T_340 & _T_701; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 286:194:@60978.4]
  assign x783_x432_D21 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@60963.4 package.scala 96:25:@60964.4]
  assign _T_703 = _T_702 & x783_x432_D21; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 286:283:@60979.4]
  assign _T_704 = _T_703 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 286:291:@60980.4]
  assign x435_rdcol_number = x435_rdcol_1_io_result; // @[Math.scala 154:22:@60999.4 Math.scala 155:14:@61000.4]
  assign _T_719 = $signed(x435_rdcol_number); // @[Math.scala 476:37:@61005.4]
  assign x436 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@61013.4 package.scala 96:25:@61014.4]
  assign x437 = x765_x414_D1 | x436; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 294:24:@61017.4]
  assign _T_767 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@61094.4 package.scala 96:25:@61095.4]
  assign _T_769 = io_rr ? _T_767 : 1'h0; // @[implicits.scala 55:10:@61096.4]
  assign _T_770 = _T_340 & _T_769; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 321:194:@61097.4]
  assign x786_x438_D20 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@61082.4 package.scala 96:25:@61083.4]
  assign _T_771 = _T_770 & x786_x438_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 321:283:@61098.4]
  assign _T_772 = _T_771 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 321:291:@61099.4]
  assign x444_rdcol_number = x444_rdcol_1_io_result; // @[Math.scala 154:22:@61118.4 Math.scala 155:14:@61119.4]
  assign _T_787 = $signed(x444_rdcol_number); // @[Math.scala 476:37:@61124.4]
  assign x445 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@61132.4 package.scala 96:25:@61133.4]
  assign x446 = x765_x414_D1 | x445; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 329:59:@61136.4]
  assign _T_830 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@61202.4 package.scala 96:25:@61203.4]
  assign _T_832 = io_rr ? _T_830 : 1'h0; // @[implicits.scala 55:10:@61204.4]
  assign _T_833 = _T_340 & _T_832; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 346:194:@61205.4]
  assign x788_x447_D20 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@61190.4 package.scala 96:25:@61191.4]
  assign _T_834 = _T_833 & x788_x447_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 346:283:@61206.4]
  assign _T_835 = _T_834 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 346:291:@61207.4]
  assign x453_rdrow_number = x453_rdrow_1_io_result; // @[Math.scala 195:22:@61226.4 Math.scala 196:14:@61227.4]
  assign _T_852 = $signed(x453_rdrow_number); // @[Math.scala 406:49:@61233.4]
  assign _T_854 = $signed(_T_852) & $signed(32'sh3); // @[Math.scala 406:56:@61235.4]
  assign _T_855 = $signed(_T_854); // @[Math.scala 406:56:@61236.4]
  assign x730_number = $unsigned(_T_855); // @[implicits.scala 133:21:@61237.4]
  assign x455 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@61251.4 package.scala 96:25:@61252.4]
  assign x456 = x455 | x415; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 356:24:@61255.4]
  assign _T_878 = $signed(x730_number); // @[Math.scala 406:49:@61264.4]
  assign _T_880 = $signed(_T_878) & $signed(32'sh3); // @[Math.scala 406:56:@61266.4]
  assign _T_881 = $signed(_T_880); // @[Math.scala 406:56:@61267.4]
  assign _T_885 = $signed(RetimeWrapper_62_io_out); // @[package.scala 96:25:@61275.4]
  assign _T_889 = x730_number[31]; // @[FixedPoint.scala 50:25:@61282.4]
  assign _T_893 = _T_889 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@61284.4]
  assign _T_894 = x730_number[31:2]; // @[FixedPoint.scala 18:52:@61285.4]
  assign _T_900 = _T_894 == 30'h3fffffff; // @[Math.scala 451:55:@61287.4]
  assign _T_901 = x730_number[1:0]; // @[FixedPoint.scala 18:52:@61288.4]
  assign _T_907 = _T_901 != 2'h0; // @[Math.scala 451:110:@61290.4]
  assign _T_908 = _T_900 & _T_907; // @[Math.scala 451:94:@61291.4]
  assign _T_912 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@61299.4 package.scala 96:25:@61300.4]
  assign x459_1_number = _T_908 ? 32'h0 : _T_912; // @[Math.scala 454:20:@61301.4]
  assign _GEN_2 = {{8'd0}, x459_1_number}; // @[Math.scala 461:32:@61306.4]
  assign _T_917 = _GEN_2 << 8; // @[Math.scala 461:32:@61306.4]
  assign _GEN_3 = {{6'd0}, x459_1_number}; // @[Math.scala 461:32:@61311.4]
  assign _T_920 = _GEN_3 << 6; // @[Math.scala 461:32:@61311.4]
  assign _T_950 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@61379.4 package.scala 96:25:@61380.4]
  assign _T_952 = io_rr ? _T_950 : 1'h0; // @[implicits.scala 55:10:@61381.4]
  assign _T_953 = _T_340 & _T_952; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 383:194:@61382.4]
  assign x791_x457_D20 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@61358.4 package.scala 96:25:@61359.4]
  assign _T_954 = _T_953 & x791_x457_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 383:283:@61383.4]
  assign _T_955 = _T_954 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 383:291:@61384.4]
  assign x464 = x455 | x420; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 387:24:@61395.4]
  assign _T_982 = RetimeWrapper_71_io_out; // @[package.scala 96:25:@61437.4 package.scala 96:25:@61438.4]
  assign _T_984 = io_rr ? _T_982 : 1'h0; // @[implicits.scala 55:10:@61439.4]
  assign _T_985 = _T_340 & _T_984; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 400:194:@61440.4]
  assign x794_x465_D20 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@61425.4 package.scala 96:25:@61426.4]
  assign _T_986 = _T_985 & x794_x465_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 400:283:@61441.4]
  assign _T_987 = _T_986 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 400:291:@61442.4]
  assign x469 = x455 | x425; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 404:24:@61453.4]
  assign _T_1014 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@61495.4 package.scala 96:25:@61496.4]
  assign _T_1016 = io_rr ? _T_1014 : 1'h0; // @[implicits.scala 55:10:@61497.4]
  assign _T_1017 = _T_340 & _T_1016; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 423:194:@61498.4]
  assign x796_x470_D20 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@61483.4 package.scala 96:25:@61484.4]
  assign _T_1018 = _T_1017 & x796_x470_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 423:283:@61499.4]
  assign _T_1019 = _T_1018 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 423:326:@61500.4]
  assign x797_x430_D1 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@61516.4 package.scala 96:25:@61517.4]
  assign x474 = x455 | x797_x430_D1; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 429:59:@61520.4]
  assign _T_1057 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@61582.4 package.scala 96:25:@61583.4]
  assign _T_1059 = io_rr ? _T_1057 : 1'h0; // @[implicits.scala 55:10:@61584.4]
  assign _T_1060 = _T_340 & _T_1059; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 448:194:@61585.4]
  assign x800_x475_D20 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@61561.4 package.scala 96:25:@61562.4]
  assign _T_1061 = _T_1060 & x800_x475_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 448:283:@61586.4]
  assign _T_1062 = _T_1061 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 448:291:@61587.4]
  assign x479 = x455 | x436; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 452:59:@61598.4]
  assign _T_1086 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@61631.4 package.scala 96:25:@61632.4]
  assign _T_1088 = io_rr ? _T_1086 : 1'h0; // @[implicits.scala 55:10:@61633.4]
  assign _T_1089 = _T_340 & _T_1088; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 463:194:@61634.4]
  assign x802_x480_D20 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@61619.4 package.scala 96:25:@61620.4]
  assign _T_1090 = _T_1089 & x802_x480_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 463:283:@61635.4]
  assign _T_1091 = _T_1090 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 463:291:@61636.4]
  assign x484 = x455 | x445; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 467:59:@61647.4]
  assign _T_1115 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@61680.4 package.scala 96:25:@61681.4]
  assign _T_1117 = io_rr ? _T_1115 : 1'h0; // @[implicits.scala 55:10:@61682.4]
  assign _T_1118 = _T_340 & _T_1117; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 478:194:@61683.4]
  assign x803_x485_D20 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@61668.4 package.scala 96:25:@61669.4]
  assign _T_1119 = _T_1118 & x803_x485_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 478:283:@61684.4]
  assign _T_1120 = _T_1119 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 478:291:@61685.4]
  assign x489_rdrow_number = x489_rdrow_1_io_result; // @[Math.scala 195:22:@61704.4 Math.scala 196:14:@61705.4]
  assign _T_1137 = $signed(x489_rdrow_number); // @[Math.scala 406:49:@61711.4]
  assign _T_1139 = $signed(_T_1137) & $signed(32'sh3); // @[Math.scala 406:56:@61713.4]
  assign _T_1140 = $signed(_T_1139); // @[Math.scala 406:56:@61714.4]
  assign x735_number = $unsigned(_T_1140); // @[implicits.scala 133:21:@61715.4]
  assign x491 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@61729.4 package.scala 96:25:@61730.4]
  assign x492 = x491 | x415; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 488:24:@61733.4]
  assign _T_1163 = $signed(x735_number); // @[Math.scala 406:49:@61742.4]
  assign _T_1165 = $signed(_T_1163) & $signed(32'sh3); // @[Math.scala 406:56:@61744.4]
  assign _T_1166 = $signed(_T_1165); // @[Math.scala 406:56:@61745.4]
  assign _T_1170 = $signed(RetimeWrapper_86_io_out); // @[package.scala 96:25:@61753.4]
  assign _T_1174 = x735_number[31]; // @[FixedPoint.scala 50:25:@61760.4]
  assign _T_1178 = _T_1174 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@61762.4]
  assign _T_1179 = x735_number[31:2]; // @[FixedPoint.scala 18:52:@61763.4]
  assign _T_1185 = _T_1179 == 30'h3fffffff; // @[Math.scala 451:55:@61765.4]
  assign _T_1186 = x735_number[1:0]; // @[FixedPoint.scala 18:52:@61766.4]
  assign _T_1192 = _T_1186 != 2'h0; // @[Math.scala 451:110:@61768.4]
  assign _T_1193 = _T_1185 & _T_1192; // @[Math.scala 451:94:@61769.4]
  assign _T_1197 = RetimeWrapper_87_io_out; // @[package.scala 96:25:@61777.4 package.scala 96:25:@61778.4]
  assign x495_1_number = _T_1193 ? 32'h0 : _T_1197; // @[Math.scala 454:20:@61779.4]
  assign _GEN_4 = {{8'd0}, x495_1_number}; // @[Math.scala 461:32:@61784.4]
  assign _T_1202 = _GEN_4 << 8; // @[Math.scala 461:32:@61784.4]
  assign _GEN_5 = {{6'd0}, x495_1_number}; // @[Math.scala 461:32:@61789.4]
  assign _T_1205 = _GEN_5 << 6; // @[Math.scala 461:32:@61789.4]
  assign _T_1232 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@61848.4 package.scala 96:25:@61849.4]
  assign _T_1234 = io_rr ? _T_1232 : 1'h0; // @[implicits.scala 55:10:@61850.4]
  assign _T_1235 = _T_340 & _T_1234; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 513:194:@61851.4]
  assign x805_x493_D20 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@61827.4 package.scala 96:25:@61828.4]
  assign _T_1236 = _T_1235 & x805_x493_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 513:283:@61852.4]
  assign _T_1237 = _T_1236 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 513:291:@61853.4]
  assign x500 = x491 | x420; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 517:24:@61864.4]
  assign _T_1261 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@61897.4 package.scala 96:25:@61898.4]
  assign _T_1263 = io_rr ? _T_1261 : 1'h0; // @[implicits.scala 55:10:@61899.4]
  assign _T_1264 = _T_340 & _T_1263; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 528:194:@61900.4]
  assign x807_x501_D20 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@61885.4 package.scala 96:25:@61886.4]
  assign _T_1265 = _T_1264 & x807_x501_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 528:283:@61901.4]
  assign _T_1266 = _T_1265 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 528:291:@61902.4]
  assign x505 = x491 | x425; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 532:24:@61913.4]
  assign _T_1290 = RetimeWrapper_95_io_out; // @[package.scala 96:25:@61946.4 package.scala 96:25:@61947.4]
  assign _T_1292 = io_rr ? _T_1290 : 1'h0; // @[implicits.scala 55:10:@61948.4]
  assign _T_1293 = _T_340 & _T_1292; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 549:194:@61949.4]
  assign x808_x506_D20 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@61934.4 package.scala 96:25:@61935.4]
  assign _T_1294 = _T_1293 & x808_x506_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 549:283:@61950.4]
  assign _T_1295 = _T_1294 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 549:291:@61951.4]
  assign x510 = x491 | x797_x430_D1; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 553:59:@61962.4]
  assign _T_1327 = RetimeWrapper_99_io_out; // @[package.scala 96:25:@62015.4 package.scala 96:25:@62016.4]
  assign _T_1329 = io_rr ? _T_1327 : 1'h0; // @[implicits.scala 55:10:@62017.4]
  assign _T_1330 = _T_340 & _T_1329; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 570:194:@62018.4]
  assign x810_x511_D20 = RetimeWrapper_97_io_out; // @[package.scala 96:25:@61994.4 package.scala 96:25:@61995.4]
  assign _T_1331 = _T_1330 & x810_x511_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 570:283:@62019.4]
  assign _T_1332 = _T_1331 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 570:291:@62020.4]
  assign x515 = x491 | x436; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 574:59:@62031.4]
  assign _T_1356 = RetimeWrapper_101_io_out; // @[package.scala 96:25:@62064.4 package.scala 96:25:@62065.4]
  assign _T_1358 = io_rr ? _T_1356 : 1'h0; // @[implicits.scala 55:10:@62066.4]
  assign _T_1359 = _T_340 & _T_1358; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 585:194:@62067.4]
  assign x812_x516_D20 = RetimeWrapper_100_io_out; // @[package.scala 96:25:@62052.4 package.scala 96:25:@62053.4]
  assign _T_1360 = _T_1359 & x812_x516_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 585:283:@62068.4]
  assign _T_1361 = _T_1360 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 585:291:@62069.4]
  assign x520 = x491 | x445; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 589:59:@62080.4]
  assign _T_1385 = RetimeWrapper_103_io_out; // @[package.scala 96:25:@62113.4 package.scala 96:25:@62114.4]
  assign _T_1387 = io_rr ? _T_1385 : 1'h0; // @[implicits.scala 55:10:@62115.4]
  assign _T_1388 = _T_340 & _T_1387; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 600:194:@62116.4]
  assign x813_x521_D20 = RetimeWrapper_102_io_out; // @[package.scala 96:25:@62101.4 package.scala 96:25:@62102.4]
  assign _T_1389 = _T_1388 & x813_x521_D20; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 600:283:@62117.4]
  assign _T_1390 = _T_1389 & x766_b379_D48; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 600:291:@62118.4]
  assign _T_1790 = RetimeWrapper_114_io_out; // @[package.scala 96:25:@63030.4 package.scala 96:25:@63031.4]
  assign _T_1792 = io_rr ? _T_1790 : 1'h0; // @[implicits.scala 55:10:@63032.4]
  assign _T_1793 = _T_340 & _T_1792; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 792:167:@63033.4]
  assign _T_1795 = _T_1793 & _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 792:256:@63035.4]
  assign _T_1796 = _T_1795 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 792:275:@63036.4]
  assign x818_b379_D67 = RetimeWrapper_108_io_out; // @[package.scala 96:25:@62974.4 package.scala 96:25:@62975.4]
  assign _T_1797 = _T_1796 & x818_b379_D67; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 792:301:@63037.4]
  assign x820_b380_D67 = RetimeWrapper_110_io_out; // @[package.scala 96:25:@62992.4 package.scala 96:25:@62993.4]
  assign _T_1813 = RetimeWrapper_118_io_out; // @[package.scala 96:25:@63080.4 package.scala 96:25:@63081.4]
  assign _T_1815 = io_rr ? _T_1813 : 1'h0; // @[implicits.scala 55:10:@63082.4]
  assign _T_1816 = _T_340 & _T_1815; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 803:167:@63083.4]
  assign _T_1818 = _T_1816 & _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 803:256:@63085.4]
  assign _T_1819 = _T_1818 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 803:275:@63086.4]
  assign _T_1820 = _T_1819 & x818_b379_D67; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 803:301:@63087.4]
  assign _T_1836 = RetimeWrapper_122_io_out; // @[package.scala 96:25:@63130.4 package.scala 96:25:@63131.4]
  assign _T_1838 = io_rr ? _T_1836 : 1'h0; // @[implicits.scala 55:10:@63132.4]
  assign _T_1839 = _T_340 & _T_1838; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 814:167:@63133.4]
  assign _T_1841 = _T_1839 & _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 814:256:@63135.4]
  assign _T_1842 = _T_1841 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 814:275:@63136.4]
  assign _T_1843 = _T_1842 & x818_b379_D67; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 814:301:@63137.4]
  assign _T_1859 = RetimeWrapper_126_io_out; // @[package.scala 96:25:@63180.4 package.scala 96:25:@63181.4]
  assign _T_1861 = io_rr ? _T_1859 : 1'h0; // @[implicits.scala 55:10:@63182.4]
  assign _T_1862 = _T_340 & _T_1861; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 825:167:@63183.4]
  assign _T_1864 = _T_1862 & _T_340; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 825:256:@63185.4]
  assign _T_1865 = _T_1864 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 825:275:@63186.4]
  assign _T_1866 = _T_1865 & x818_b379_D67; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 825:301:@63187.4]
  assign _T_1897 = RetimeWrapper_133_io_out; // @[package.scala 96:25:@63258.4 package.scala 96:25:@63259.4]
  assign _T_1899 = io_rr ? _T_1897 : 1'h0; // @[implicits.scala 55:10:@63260.4]
  assign _T_1900 = _T_340 & _T_1899; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 843:195:@63261.4]
  assign x834_x417_D40 = RetimeWrapper_128_io_out; // @[package.scala 96:25:@63210.4 package.scala 96:25:@63211.4]
  assign _T_1901 = _T_1900 & x834_x417_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 843:284:@63262.4]
  assign x833_b379_D68 = RetimeWrapper_127_io_out; // @[package.scala 96:25:@63201.4 package.scala 96:25:@63202.4]
  assign _T_1902 = _T_1901 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 843:292:@63263.4]
  assign x836_b380_D68 = RetimeWrapper_130_io_out; // @[package.scala 96:25:@63228.4 package.scala 96:25:@63229.4]
  assign _T_1925 = RetimeWrapper_137_io_out; // @[package.scala 96:25:@63309.4 package.scala 96:25:@63310.4]
  assign _T_1927 = io_rr ? _T_1925 : 1'h0; // @[implicits.scala 55:10:@63311.4]
  assign _T_1928 = _T_340 & _T_1927; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 856:195:@63312.4]
  assign x841_x422_D40 = RetimeWrapper_136_io_out; // @[package.scala 96:25:@63297.4 package.scala 96:25:@63298.4]
  assign _T_1929 = _T_1928 & x841_x422_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 856:284:@63313.4]
  assign _T_1930 = _T_1929 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 856:292:@63314.4]
  assign _T_1953 = RetimeWrapper_141_io_out; // @[package.scala 96:25:@63360.4 package.scala 96:25:@63361.4]
  assign _T_1955 = io_rr ? _T_1953 : 1'h0; // @[implicits.scala 55:10:@63362.4]
  assign _T_1956 = _T_340 & _T_1955; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 869:195:@63363.4]
  assign x844_x427_D40 = RetimeWrapper_140_io_out; // @[package.scala 96:25:@63348.4 package.scala 96:25:@63349.4]
  assign _T_1957 = _T_1956 & x844_x427_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 869:284:@63364.4]
  assign _T_1958 = _T_1957 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 869:292:@63365.4]
  assign _T_1981 = RetimeWrapper_145_io_out; // @[package.scala 96:25:@63411.4 package.scala 96:25:@63412.4]
  assign _T_1983 = io_rr ? _T_1981 : 1'h0; // @[implicits.scala 55:10:@63413.4]
  assign _T_1984 = _T_340 & _T_1983; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 882:195:@63414.4]
  assign x847_x432_D41 = RetimeWrapper_144_io_out; // @[package.scala 96:25:@63399.4 package.scala 96:25:@63400.4]
  assign _T_1985 = _T_1984 & x847_x432_D41; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 882:284:@63415.4]
  assign _T_1986 = _T_1985 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 882:292:@63416.4]
  assign _T_2009 = RetimeWrapper_149_io_out; // @[package.scala 96:25:@63462.4 package.scala 96:25:@63463.4]
  assign _T_2011 = io_rr ? _T_2009 : 1'h0; // @[implicits.scala 55:10:@63464.4]
  assign _T_2012 = _T_340 & _T_2011; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 901:195:@63465.4]
  assign x849_x438_D40 = RetimeWrapper_147_io_out; // @[package.scala 96:25:@63441.4 package.scala 96:25:@63442.4]
  assign _T_2013 = _T_2012 & x849_x438_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 901:284:@63466.4]
  assign _T_2014 = _T_2013 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 901:327:@63467.4]
  assign _T_2037 = RetimeWrapper_153_io_out; // @[package.scala 96:25:@63513.4 package.scala 96:25:@63514.4]
  assign _T_2039 = io_rr ? _T_2037 : 1'h0; // @[implicits.scala 55:10:@63515.4]
  assign _T_2040 = _T_340 & _T_2039; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 914:195:@63516.4]
  assign x852_x457_D40 = RetimeWrapper_151_io_out; // @[package.scala 96:25:@63492.4 package.scala 96:25:@63493.4]
  assign _T_2041 = _T_2040 & x852_x457_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 914:284:@63517.4]
  assign _T_2042 = _T_2041 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 914:292:@63518.4]
  assign _T_2062 = RetimeWrapper_156_io_out; // @[package.scala 96:25:@63555.4 package.scala 96:25:@63556.4]
  assign _T_2064 = io_rr ? _T_2062 : 1'h0; // @[implicits.scala 55:10:@63557.4]
  assign _T_2065 = _T_340 & _T_2064; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 925:195:@63558.4]
  assign x855_x465_D40 = RetimeWrapper_155_io_out; // @[package.scala 96:25:@63543.4 package.scala 96:25:@63544.4]
  assign _T_2066 = _T_2065 & x855_x465_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 925:284:@63559.4]
  assign _T_2067 = _T_2066 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 925:292:@63560.4]
  assign _T_2087 = RetimeWrapper_159_io_out; // @[package.scala 96:25:@63597.4 package.scala 96:25:@63598.4]
  assign _T_2089 = io_rr ? _T_2087 : 1'h0; // @[implicits.scala 55:10:@63599.4]
  assign _T_2090 = _T_340 & _T_2089; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 936:195:@63600.4]
  assign x857_x470_D40 = RetimeWrapper_158_io_out; // @[package.scala 96:25:@63585.4 package.scala 96:25:@63586.4]
  assign _T_2091 = _T_2090 & x857_x470_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 936:284:@63601.4]
  assign _T_2092 = _T_2091 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 936:292:@63602.4]
  assign _T_2112 = RetimeWrapper_162_io_out; // @[package.scala 96:25:@63639.4 package.scala 96:25:@63640.4]
  assign _T_2114 = io_rr ? _T_2112 : 1'h0; // @[implicits.scala 55:10:@63641.4]
  assign _T_2115 = _T_340 & _T_2114; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 947:195:@63642.4]
  assign x858_x475_D40 = RetimeWrapper_160_io_out; // @[package.scala 96:25:@63618.4 package.scala 96:25:@63619.4]
  assign _T_2116 = _T_2115 & x858_x475_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 947:284:@63643.4]
  assign _T_2117 = _T_2116 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 947:292:@63644.4]
  assign _T_2137 = RetimeWrapper_165_io_out; // @[package.scala 96:25:@63681.4 package.scala 96:25:@63682.4]
  assign _T_2139 = io_rr ? _T_2137 : 1'h0; // @[implicits.scala 55:10:@63683.4]
  assign _T_2140 = _T_340 & _T_2139; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 958:195:@63684.4]
  assign x861_x480_D40 = RetimeWrapper_164_io_out; // @[package.scala 96:25:@63669.4 package.scala 96:25:@63670.4]
  assign _T_2141 = _T_2140 & x861_x480_D40; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 958:284:@63685.4]
  assign _T_2142 = _T_2141 & x833_b379_D68; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 958:292:@63686.4]
  assign x654_number = x654_1_io_result; // @[Math.scala 723:22:@64021.4 Math.scala 724:14:@64022.4]
  assign x664_number = x664_1_io_result; // @[Math.scala 723:22:@64129.4 Math.scala 724:14:@64130.4]
  assign _T_2360 = {x654_number,x664_number}; // @[Cat.scala 30:58:@64138.4]
  assign x634_number = x634_1_io_result; // @[Math.scala 723:22:@63803.4 Math.scala 724:14:@63804.4]
  assign x644_number = x644_1_io_result; // @[Math.scala 723:22:@63911.4 Math.scala 724:14:@63912.4]
  assign _T_2361 = {x634_number,x644_number}; // @[Cat.scala 30:58:@64139.4]
  assign _T_2374 = RetimeWrapper_169_io_out; // @[package.scala 96:25:@64175.4 package.scala 96:25:@64176.4]
  assign _T_2376 = io_rr ? _T_2374 : 1'h0; // @[implicits.scala 55:10:@64177.4]
  assign x863_b379_D87 = RetimeWrapper_168_io_out; // @[package.scala 96:25:@64166.4 package.scala 96:25:@64167.4]
  assign _T_2377 = _T_2376 & x863_b379_D87; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1060:117:@64178.4]
  assign x862_b380_D87 = RetimeWrapper_167_io_out; // @[package.scala 96:25:@64157.4 package.scala 96:25:@64158.4]
  assign _T_2378 = _T_2377 & x862_b380_D87; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1060:123:@64179.4]
  assign x748_x389_D8_number = RetimeWrapper_3_io_out; // @[package.scala 96:25:@60244.4 package.scala 96:25:@60245.4]
  assign x750_x393_sum_D3_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@60262.4 package.scala 96:25:@60263.4]
  assign x752_x726_D24_number = RetimeWrapper_7_io_out; // @[package.scala 96:25:@60280.4 package.scala 96:25:@60281.4]
  assign x754_x397_D7_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@60369.4 package.scala 96:25:@60370.4]
  assign x756_x399_sum_D2_number = RetimeWrapper_12_io_out; // @[package.scala 96:25:@60387.4 package.scala 96:25:@60388.4]
  assign x757_x403_D7_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@60467.4 package.scala 96:25:@60468.4]
  assign x759_x405_sum_D2_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@60485.4 package.scala 96:25:@60486.4]
  assign x761_x411_sum_D2_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@60574.4 package.scala 96:25:@60575.4]
  assign x762_x409_D7_number = RetimeWrapper_20_io_out; // @[package.scala 96:25:@60583.4 package.scala 96:25:@60584.4]
  assign x768_x411_sum_D26_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@60696.4 package.scala 96:25:@60697.4]
  assign x770_x726_D48_number = RetimeWrapper_31_io_out; // @[package.scala 96:25:@60714.4 package.scala 96:25:@60715.4]
  assign x771_x409_D31_number = RetimeWrapper_32_io_out; // @[package.scala 96:25:@60723.4 package.scala 96:25:@60724.4]
  assign x773_x403_D31_number = RetimeWrapper_36_io_out; // @[package.scala 96:25:@60785.4 package.scala 96:25:@60786.4]
  assign x774_x405_sum_D26_number = RetimeWrapper_37_io_out; // @[package.scala 96:25:@60794.4 package.scala 96:25:@60795.4]
  assign x777_x397_D31_number = RetimeWrapper_42_io_out; // @[package.scala 96:25:@60865.4 package.scala 96:25:@60866.4]
  assign x778_x399_sum_D26_number = RetimeWrapper_43_io_out; // @[package.scala 96:25:@60874.4 package.scala 96:25:@60875.4]
  assign x781_x389_D32_number = RetimeWrapper_48_io_out; // @[package.scala 96:25:@60945.4 package.scala 96:25:@60946.4]
  assign x782_x393_sum_D27_number = RetimeWrapper_49_io_out; // @[package.scala 96:25:@60954.4 package.scala 96:25:@60955.4]
  assign x441_sum_number = x441_sum_1_io_result; // @[Math.scala 154:22:@61064.4 Math.scala 155:14:@61065.4]
  assign x785_x439_D5_number = RetimeWrapper_54_io_out; // @[package.scala 96:25:@61073.4 package.scala 96:25:@61074.4]
  assign x450_sum_number = x450_sum_1_io_result; // @[Math.scala 154:22:@61172.4 Math.scala 155:14:@61173.4]
  assign x787_x448_D5_number = RetimeWrapper_58_io_out; // @[package.scala 96:25:@61181.4 package.scala 96:25:@61182.4]
  assign x461_sum_number = x461_sum_1_io_result; // @[Math.scala 154:22:@61349.4 Math.scala 155:14:@61350.4]
  assign x792_x731_D20_number = RetimeWrapper_67_io_out; // @[package.scala 96:25:@61367.4 package.scala 96:25:@61368.4]
  assign x466_sum_number = x466_sum_1_io_result; // @[Math.scala 154:22:@61416.4 Math.scala 155:14:@61417.4]
  assign x471_sum_number = x471_sum_1_io_result; // @[Math.scala 154:22:@61474.4 Math.scala 155:14:@61475.4]
  assign x801_x476_sum_D1_number = RetimeWrapper_79_io_out; // @[package.scala 96:25:@61570.4 package.scala 96:25:@61571.4]
  assign x481_sum_number = x481_sum_1_io_result; // @[Math.scala 154:22:@61610.4 Math.scala 155:14:@61611.4]
  assign x486_sum_number = x486_sum_1_io_result; // @[Math.scala 154:22:@61659.4 Math.scala 155:14:@61660.4]
  assign x497_sum_number = x497_sum_1_io_result; // @[Math.scala 154:22:@61818.4 Math.scala 155:14:@61819.4]
  assign x806_x736_D20_number = RetimeWrapper_90_io_out; // @[package.scala 96:25:@61836.4 package.scala 96:25:@61837.4]
  assign x502_sum_number = x502_sum_1_io_result; // @[Math.scala 154:22:@61876.4 Math.scala 155:14:@61877.4]
  assign x507_sum_number = x507_sum_1_io_result; // @[Math.scala 154:22:@61925.4 Math.scala 155:14:@61926.4]
  assign x811_x512_sum_D1_number = RetimeWrapper_98_io_out; // @[package.scala 96:25:@62003.4 package.scala 96:25:@62004.4]
  assign x517_sum_number = x517_sum_1_io_result; // @[Math.scala 154:22:@62043.4 Math.scala 155:14:@62044.4]
  assign x522_sum_number = x522_sum_1_io_result; // @[Math.scala 154:22:@62092.4 Math.scala 155:14:@62093.4]
  assign x819_x389_D51_number = RetimeWrapper_109_io_out; // @[package.scala 96:25:@62983.4 package.scala 96:25:@62984.4]
  assign x822_x393_sum_D46_number = RetimeWrapper_112_io_out; // @[package.scala 96:25:@63010.4 package.scala 96:25:@63011.4]
  assign x823_x726_D67_number = RetimeWrapper_113_io_out; // @[package.scala 96:25:@63019.4 package.scala 96:25:@63020.4]
  assign x824_x397_D50_number = RetimeWrapper_115_io_out; // @[package.scala 96:25:@63051.4 package.scala 96:25:@63052.4]
  assign x825_x399_sum_D45_number = RetimeWrapper_116_io_out; // @[package.scala 96:25:@63060.4 package.scala 96:25:@63061.4]
  assign x827_x403_D50_number = RetimeWrapper_119_io_out; // @[package.scala 96:25:@63101.4 package.scala 96:25:@63102.4]
  assign x828_x405_sum_D45_number = RetimeWrapper_120_io_out; // @[package.scala 96:25:@63110.4 package.scala 96:25:@63111.4]
  assign x830_x411_sum_D45_number = RetimeWrapper_123_io_out; // @[package.scala 96:25:@63151.4 package.scala 96:25:@63152.4]
  assign x831_x409_D50_number = RetimeWrapper_124_io_out; // @[package.scala 96:25:@63160.4 package.scala 96:25:@63161.4]
  assign x835_x411_sum_D46_number = RetimeWrapper_129_io_out; // @[package.scala 96:25:@63219.4 package.scala 96:25:@63220.4]
  assign x837_x726_D68_number = RetimeWrapper_131_io_out; // @[package.scala 96:25:@63237.4 package.scala 96:25:@63238.4]
  assign x838_x409_D51_number = RetimeWrapper_132_io_out; // @[package.scala 96:25:@63246.4 package.scala 96:25:@63247.4]
  assign x839_x403_D51_number = RetimeWrapper_134_io_out; // @[package.scala 96:25:@63279.4 package.scala 96:25:@63280.4]
  assign x840_x405_sum_D46_number = RetimeWrapper_135_io_out; // @[package.scala 96:25:@63288.4 package.scala 96:25:@63289.4]
  assign x842_x397_D51_number = RetimeWrapper_138_io_out; // @[package.scala 96:25:@63330.4 package.scala 96:25:@63331.4]
  assign x843_x399_sum_D46_number = RetimeWrapper_139_io_out; // @[package.scala 96:25:@63339.4 package.scala 96:25:@63340.4]
  assign x845_x389_D52_number = RetimeWrapper_142_io_out; // @[package.scala 96:25:@63381.4 package.scala 96:25:@63382.4]
  assign x846_x393_sum_D47_number = RetimeWrapper_143_io_out; // @[package.scala 96:25:@63390.4 package.scala 96:25:@63391.4]
  assign x848_x439_D25_number = RetimeWrapper_146_io_out; // @[package.scala 96:25:@63432.4 package.scala 96:25:@63433.4]
  assign x850_x441_sum_D20_number = RetimeWrapper_148_io_out; // @[package.scala 96:25:@63450.4 package.scala 96:25:@63451.4]
  assign x851_x461_sum_D20_number = RetimeWrapper_150_io_out; // @[package.scala 96:25:@63483.4 package.scala 96:25:@63484.4]
  assign x853_x731_D40_number = RetimeWrapper_152_io_out; // @[package.scala 96:25:@63501.4 package.scala 96:25:@63502.4]
  assign x854_x466_sum_D20_number = RetimeWrapper_154_io_out; // @[package.scala 96:25:@63534.4 package.scala 96:25:@63535.4]
  assign x856_x471_sum_D20_number = RetimeWrapper_157_io_out; // @[package.scala 96:25:@63576.4 package.scala 96:25:@63577.4]
  assign x859_x476_sum_D21_number = RetimeWrapper_161_io_out; // @[package.scala 96:25:@63627.4 package.scala 96:25:@63628.4]
  assign x860_x481_sum_D20_number = RetimeWrapper_163_io_out; // @[package.scala 96:25:@63660.4 package.scala 96:25:@63661.4]
  assign io_in_x343_TVALID = _T_2378 & io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1060:22:@64181.4]
  assign io_in_x343_TDATA = {{128'd0}, RetimeWrapper_166_io_out}; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1061:24:@64182.4]
  assign io_in_x342_TREADY = _T_211 & _T_213; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 67:22:@59852.4 sm_x669_inr_Foreach_SAMPLER_BOX.scala 69:22:@59860.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@59830.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@59842.4]
  assign RetimeWrapper_clock = clock; // @[:@59863.4]
  assign RetimeWrapper_reset = reset; // @[:@59864.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@59866.4]
  assign RetimeWrapper_io_in = io_in_x342_TDATA[127:0]; // @[package.scala 94:16:@59865.4]
  assign x383_lb_0_clock = clock; // @[:@59873.4]
  assign x383_lb_0_reset = reset; // @[:@59874.4]
  assign x383_lb_0_io_rPort_17_banks_1 = x785_x439_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@61102.4]
  assign x383_lb_0_io_rPort_17_banks_0 = x770_x726_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@61101.4]
  assign x383_lb_0_io_rPort_17_ofs_0 = x441_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61103.4]
  assign x383_lb_0_io_rPort_17_en_0 = _T_772 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61105.4]
  assign x383_lb_0_io_rPort_17_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61104.4]
  assign x383_lb_0_io_rPort_16_banks_1 = x781_x389_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@60983.4]
  assign x383_lb_0_io_rPort_16_banks_0 = x770_x726_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@60982.4]
  assign x383_lb_0_io_rPort_16_ofs_0 = x782_x393_sum_D27_number[8:0]; // @[MemInterfaceType.scala 107:54:@60984.4]
  assign x383_lb_0_io_rPort_16_en_0 = _T_704 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@60986.4]
  assign x383_lb_0_io_rPort_16_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@60985.4]
  assign x383_lb_0_io_rPort_15_banks_1 = x771_x409_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@60743.4]
  assign x383_lb_0_io_rPort_15_banks_0 = x770_x726_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@60742.4]
  assign x383_lb_0_io_rPort_15_ofs_0 = x768_x411_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@60744.4]
  assign x383_lb_0_io_rPort_15_en_0 = _T_569 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@60746.4]
  assign x383_lb_0_io_rPort_15_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@60745.4]
  assign x383_lb_0_io_rPort_14_banks_1 = x785_x439_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@61639.4]
  assign x383_lb_0_io_rPort_14_banks_0 = x792_x731_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61638.4]
  assign x383_lb_0_io_rPort_14_ofs_0 = x481_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61640.4]
  assign x383_lb_0_io_rPort_14_en_0 = _T_1091 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61642.4]
  assign x383_lb_0_io_rPort_14_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61641.4]
  assign x383_lb_0_io_rPort_13_banks_1 = x787_x448_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@61688.4]
  assign x383_lb_0_io_rPort_13_banks_0 = x792_x731_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61687.4]
  assign x383_lb_0_io_rPort_13_ofs_0 = x486_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61689.4]
  assign x383_lb_0_io_rPort_13_en_0 = _T_1120 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61691.4]
  assign x383_lb_0_io_rPort_13_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61690.4]
  assign x383_lb_0_io_rPort_12_banks_1 = x771_x409_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@61387.4]
  assign x383_lb_0_io_rPort_12_banks_0 = x792_x731_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61386.4]
  assign x383_lb_0_io_rPort_12_ofs_0 = x461_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61388.4]
  assign x383_lb_0_io_rPort_12_en_0 = _T_955 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61390.4]
  assign x383_lb_0_io_rPort_12_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61389.4]
  assign x383_lb_0_io_rPort_11_banks_1 = x781_x389_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@61590.4]
  assign x383_lb_0_io_rPort_11_banks_0 = x792_x731_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61589.4]
  assign x383_lb_0_io_rPort_11_ofs_0 = x801_x476_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@61591.4]
  assign x383_lb_0_io_rPort_11_en_0 = _T_1062 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61593.4]
  assign x383_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61592.4]
  assign x383_lb_0_io_rPort_10_banks_1 = x787_x448_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@61210.4]
  assign x383_lb_0_io_rPort_10_banks_0 = x770_x726_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@61209.4]
  assign x383_lb_0_io_rPort_10_ofs_0 = x450_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61211.4]
  assign x383_lb_0_io_rPort_10_en_0 = _T_835 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61213.4]
  assign x383_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61212.4]
  assign x383_lb_0_io_rPort_9_banks_1 = x771_x409_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@61856.4]
  assign x383_lb_0_io_rPort_9_banks_0 = x806_x736_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61855.4]
  assign x383_lb_0_io_rPort_9_ofs_0 = x497_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61857.4]
  assign x383_lb_0_io_rPort_9_en_0 = _T_1237 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61859.4]
  assign x383_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61858.4]
  assign x383_lb_0_io_rPort_8_banks_1 = x773_x403_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@60823.4]
  assign x383_lb_0_io_rPort_8_banks_0 = x770_x726_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@60822.4]
  assign x383_lb_0_io_rPort_8_ofs_0 = x774_x405_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@60824.4]
  assign x383_lb_0_io_rPort_8_en_0 = _T_614 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@60826.4]
  assign x383_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@60825.4]
  assign x383_lb_0_io_rPort_7_banks_1 = x781_x389_D32_number[2:0]; // @[MemInterfaceType.scala 106:58:@62023.4]
  assign x383_lb_0_io_rPort_7_banks_0 = x806_x736_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@62022.4]
  assign x383_lb_0_io_rPort_7_ofs_0 = x811_x512_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@62024.4]
  assign x383_lb_0_io_rPort_7_en_0 = _T_1332 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@62026.4]
  assign x383_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@62025.4]
  assign x383_lb_0_io_rPort_6_banks_1 = x777_x397_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@61954.4]
  assign x383_lb_0_io_rPort_6_banks_0 = x806_x736_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61953.4]
  assign x383_lb_0_io_rPort_6_ofs_0 = x507_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61955.4]
  assign x383_lb_0_io_rPort_6_en_0 = _T_1295 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61957.4]
  assign x383_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61956.4]
  assign x383_lb_0_io_rPort_5_banks_1 = x773_x403_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@61905.4]
  assign x383_lb_0_io_rPort_5_banks_0 = x806_x736_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61904.4]
  assign x383_lb_0_io_rPort_5_ofs_0 = x502_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61906.4]
  assign x383_lb_0_io_rPort_5_en_0 = _T_1266 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61908.4]
  assign x383_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61907.4]
  assign x383_lb_0_io_rPort_4_banks_1 = x773_x403_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@61445.4]
  assign x383_lb_0_io_rPort_4_banks_0 = x792_x731_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61444.4]
  assign x383_lb_0_io_rPort_4_ofs_0 = x466_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61446.4]
  assign x383_lb_0_io_rPort_4_en_0 = _T_987 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61448.4]
  assign x383_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61447.4]
  assign x383_lb_0_io_rPort_3_banks_1 = x777_x397_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@60903.4]
  assign x383_lb_0_io_rPort_3_banks_0 = x770_x726_D48_number[2:0]; // @[MemInterfaceType.scala 106:58:@60902.4]
  assign x383_lb_0_io_rPort_3_ofs_0 = x778_x399_sum_D26_number[8:0]; // @[MemInterfaceType.scala 107:54:@60904.4]
  assign x383_lb_0_io_rPort_3_en_0 = _T_659 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@60906.4]
  assign x383_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@60905.4]
  assign x383_lb_0_io_rPort_2_banks_1 = x777_x397_D31_number[2:0]; // @[MemInterfaceType.scala 106:58:@61503.4]
  assign x383_lb_0_io_rPort_2_banks_0 = x792_x731_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@61502.4]
  assign x383_lb_0_io_rPort_2_ofs_0 = x471_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@61504.4]
  assign x383_lb_0_io_rPort_2_en_0 = _T_1019 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@61506.4]
  assign x383_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@61505.4]
  assign x383_lb_0_io_rPort_1_banks_1 = x787_x448_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@62121.4]
  assign x383_lb_0_io_rPort_1_banks_0 = x806_x736_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@62120.4]
  assign x383_lb_0_io_rPort_1_ofs_0 = x522_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@62122.4]
  assign x383_lb_0_io_rPort_1_en_0 = _T_1390 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@62124.4]
  assign x383_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@62123.4]
  assign x383_lb_0_io_rPort_0_banks_1 = x785_x439_D5_number[2:0]; // @[MemInterfaceType.scala 106:58:@62072.4]
  assign x383_lb_0_io_rPort_0_banks_0 = x806_x736_D20_number[2:0]; // @[MemInterfaceType.scala 106:58:@62071.4]
  assign x383_lb_0_io_rPort_0_ofs_0 = x517_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@62073.4]
  assign x383_lb_0_io_rPort_0_en_0 = _T_1361 & x769_b380_D48; // @[MemInterfaceType.scala 110:79:@62075.4]
  assign x383_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@62074.4]
  assign x383_lb_0_io_wPort_3_banks_1 = x762_x409_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@60604.4]
  assign x383_lb_0_io_wPort_3_banks_0 = x752_x726_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@60603.4]
  assign x383_lb_0_io_wPort_3_ofs_0 = x761_x411_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@60605.4]
  assign x383_lb_0_io_wPort_3_data_0 = RetimeWrapper_18_io_out; // @[MemInterfaceType.scala 90:56:@60606.4]
  assign x383_lb_0_io_wPort_3_en_0 = _T_498 & x749_b380_D24; // @[MemInterfaceType.scala 93:57:@60608.4]
  assign x383_lb_0_io_wPort_2_banks_1 = x757_x403_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@60506.4]
  assign x383_lb_0_io_wPort_2_banks_0 = x752_x726_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@60505.4]
  assign x383_lb_0_io_wPort_2_ofs_0 = x759_x405_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@60507.4]
  assign x383_lb_0_io_wPort_2_data_0 = RetimeWrapper_15_io_out; // @[MemInterfaceType.scala 90:56:@60508.4]
  assign x383_lb_0_io_wPort_2_en_0 = _T_450 & x749_b380_D24; // @[MemInterfaceType.scala 93:57:@60510.4]
  assign x383_lb_0_io_wPort_1_banks_1 = x754_x397_D7_number[2:0]; // @[MemInterfaceType.scala 88:58:@60408.4]
  assign x383_lb_0_io_wPort_1_banks_0 = x752_x726_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@60407.4]
  assign x383_lb_0_io_wPort_1_ofs_0 = x756_x399_sum_D2_number[8:0]; // @[MemInterfaceType.scala 89:54:@60409.4]
  assign x383_lb_0_io_wPort_1_data_0 = RetimeWrapper_11_io_out; // @[MemInterfaceType.scala 90:56:@60410.4]
  assign x383_lb_0_io_wPort_1_en_0 = _T_402 & x749_b380_D24; // @[MemInterfaceType.scala 93:57:@60412.4]
  assign x383_lb_0_io_wPort_0_banks_1 = x748_x389_D8_number[2:0]; // @[MemInterfaceType.scala 88:58:@60301.4]
  assign x383_lb_0_io_wPort_0_banks_0 = x752_x726_D24_number[2:0]; // @[MemInterfaceType.scala 88:58:@60300.4]
  assign x383_lb_0_io_wPort_0_ofs_0 = x750_x393_sum_D3_number[8:0]; // @[MemInterfaceType.scala 89:54:@60302.4]
  assign x383_lb_0_io_wPort_0_data_0 = RetimeWrapper_6_io_out; // @[MemInterfaceType.scala 90:56:@60303.4]
  assign x383_lb_0_io_wPort_0_en_0 = _T_351 & x749_b380_D24; // @[MemInterfaceType.scala 93:57:@60305.4]
  assign x384_lb2_0_clock = clock; // @[:@60018.4]
  assign x384_lb2_0_reset = reset; // @[:@60019.4]
  assign x384_lb2_0_io_rPort_9_banks_1 = x839_x403_D51_number[2:0]; // @[MemInterfaceType.scala 106:58:@63317.4]
  assign x384_lb2_0_io_rPort_9_banks_0 = x837_x726_D68_number[2:0]; // @[MemInterfaceType.scala 106:58:@63316.4]
  assign x384_lb2_0_io_rPort_9_ofs_0 = x840_x405_sum_D46_number[8:0]; // @[MemInterfaceType.scala 107:54:@63318.4]
  assign x384_lb2_0_io_rPort_9_en_0 = _T_1930 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63320.4]
  assign x384_lb2_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63319.4]
  assign x384_lb2_0_io_rPort_8_banks_1 = x848_x439_D25_number[2:0]; // @[MemInterfaceType.scala 106:58:@63470.4]
  assign x384_lb2_0_io_rPort_8_banks_0 = x837_x726_D68_number[2:0]; // @[MemInterfaceType.scala 106:58:@63469.4]
  assign x384_lb2_0_io_rPort_8_ofs_0 = x850_x441_sum_D20_number[8:0]; // @[MemInterfaceType.scala 107:54:@63471.4]
  assign x384_lb2_0_io_rPort_8_en_0 = _T_2014 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63473.4]
  assign x384_lb2_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63472.4]
  assign x384_lb2_0_io_rPort_7_banks_1 = x839_x403_D51_number[2:0]; // @[MemInterfaceType.scala 106:58:@63563.4]
  assign x384_lb2_0_io_rPort_7_banks_0 = x853_x731_D40_number[2:0]; // @[MemInterfaceType.scala 106:58:@63562.4]
  assign x384_lb2_0_io_rPort_7_ofs_0 = x854_x466_sum_D20_number[8:0]; // @[MemInterfaceType.scala 107:54:@63564.4]
  assign x384_lb2_0_io_rPort_7_en_0 = _T_2067 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63566.4]
  assign x384_lb2_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63565.4]
  assign x384_lb2_0_io_rPort_6_banks_1 = x845_x389_D52_number[2:0]; // @[MemInterfaceType.scala 106:58:@63647.4]
  assign x384_lb2_0_io_rPort_6_banks_0 = x853_x731_D40_number[2:0]; // @[MemInterfaceType.scala 106:58:@63646.4]
  assign x384_lb2_0_io_rPort_6_ofs_0 = x859_x476_sum_D21_number[8:0]; // @[MemInterfaceType.scala 107:54:@63648.4]
  assign x384_lb2_0_io_rPort_6_en_0 = _T_2117 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63650.4]
  assign x384_lb2_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63649.4]
  assign x384_lb2_0_io_rPort_5_banks_1 = x842_x397_D51_number[2:0]; // @[MemInterfaceType.scala 106:58:@63368.4]
  assign x384_lb2_0_io_rPort_5_banks_0 = x837_x726_D68_number[2:0]; // @[MemInterfaceType.scala 106:58:@63367.4]
  assign x384_lb2_0_io_rPort_5_ofs_0 = x843_x399_sum_D46_number[8:0]; // @[MemInterfaceType.scala 107:54:@63369.4]
  assign x384_lb2_0_io_rPort_5_en_0 = _T_1958 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63371.4]
  assign x384_lb2_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63370.4]
  assign x384_lb2_0_io_rPort_4_banks_1 = x845_x389_D52_number[2:0]; // @[MemInterfaceType.scala 106:58:@63419.4]
  assign x384_lb2_0_io_rPort_4_banks_0 = x837_x726_D68_number[2:0]; // @[MemInterfaceType.scala 106:58:@63418.4]
  assign x384_lb2_0_io_rPort_4_ofs_0 = x846_x393_sum_D47_number[8:0]; // @[MemInterfaceType.scala 107:54:@63420.4]
  assign x384_lb2_0_io_rPort_4_en_0 = _T_1986 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63422.4]
  assign x384_lb2_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63421.4]
  assign x384_lb2_0_io_rPort_3_banks_1 = x838_x409_D51_number[2:0]; // @[MemInterfaceType.scala 106:58:@63266.4]
  assign x384_lb2_0_io_rPort_3_banks_0 = x837_x726_D68_number[2:0]; // @[MemInterfaceType.scala 106:58:@63265.4]
  assign x384_lb2_0_io_rPort_3_ofs_0 = x835_x411_sum_D46_number[8:0]; // @[MemInterfaceType.scala 107:54:@63267.4]
  assign x384_lb2_0_io_rPort_3_en_0 = _T_1902 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63269.4]
  assign x384_lb2_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63268.4]
  assign x384_lb2_0_io_rPort_2_banks_1 = x838_x409_D51_number[2:0]; // @[MemInterfaceType.scala 106:58:@63521.4]
  assign x384_lb2_0_io_rPort_2_banks_0 = x853_x731_D40_number[2:0]; // @[MemInterfaceType.scala 106:58:@63520.4]
  assign x384_lb2_0_io_rPort_2_ofs_0 = x851_x461_sum_D20_number[8:0]; // @[MemInterfaceType.scala 107:54:@63522.4]
  assign x384_lb2_0_io_rPort_2_en_0 = _T_2042 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63524.4]
  assign x384_lb2_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63523.4]
  assign x384_lb2_0_io_rPort_1_banks_1 = x848_x439_D25_number[2:0]; // @[MemInterfaceType.scala 106:58:@63689.4]
  assign x384_lb2_0_io_rPort_1_banks_0 = x853_x731_D40_number[2:0]; // @[MemInterfaceType.scala 106:58:@63688.4]
  assign x384_lb2_0_io_rPort_1_ofs_0 = x860_x481_sum_D20_number[8:0]; // @[MemInterfaceType.scala 107:54:@63690.4]
  assign x384_lb2_0_io_rPort_1_en_0 = _T_2142 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63692.4]
  assign x384_lb2_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63691.4]
  assign x384_lb2_0_io_rPort_0_banks_1 = x842_x397_D51_number[2:0]; // @[MemInterfaceType.scala 106:58:@63605.4]
  assign x384_lb2_0_io_rPort_0_banks_0 = x853_x731_D40_number[2:0]; // @[MemInterfaceType.scala 106:58:@63604.4]
  assign x384_lb2_0_io_rPort_0_ofs_0 = x856_x471_sum_D20_number[8:0]; // @[MemInterfaceType.scala 107:54:@63606.4]
  assign x384_lb2_0_io_rPort_0_en_0 = _T_2092 & x836_b380_D68; // @[MemInterfaceType.scala 110:79:@63608.4]
  assign x384_lb2_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@63607.4]
  assign x384_lb2_0_io_wPort_3_banks_1 = x831_x409_D50_number[2:0]; // @[MemInterfaceType.scala 88:58:@63190.4]
  assign x384_lb2_0_io_wPort_3_banks_0 = x823_x726_D67_number[2:0]; // @[MemInterfaceType.scala 88:58:@63189.4]
  assign x384_lb2_0_io_wPort_3_ofs_0 = x830_x411_sum_D45_number[8:0]; // @[MemInterfaceType.scala 89:54:@63191.4]
  assign x384_lb2_0_io_wPort_3_data_0 = RetimeWrapper_125_io_out; // @[MemInterfaceType.scala 90:56:@63192.4]
  assign x384_lb2_0_io_wPort_3_en_0 = _T_1866 & x820_b380_D67; // @[MemInterfaceType.scala 93:57:@63194.4]
  assign x384_lb2_0_io_wPort_2_banks_1 = x827_x403_D50_number[2:0]; // @[MemInterfaceType.scala 88:58:@63140.4]
  assign x384_lb2_0_io_wPort_2_banks_0 = x823_x726_D67_number[2:0]; // @[MemInterfaceType.scala 88:58:@63139.4]
  assign x384_lb2_0_io_wPort_2_ofs_0 = x828_x405_sum_D45_number[8:0]; // @[MemInterfaceType.scala 89:54:@63141.4]
  assign x384_lb2_0_io_wPort_2_data_0 = RetimeWrapper_121_io_out; // @[MemInterfaceType.scala 90:56:@63142.4]
  assign x384_lb2_0_io_wPort_2_en_0 = _T_1843 & x820_b380_D67; // @[MemInterfaceType.scala 93:57:@63144.4]
  assign x384_lb2_0_io_wPort_1_banks_1 = x824_x397_D50_number[2:0]; // @[MemInterfaceType.scala 88:58:@63090.4]
  assign x384_lb2_0_io_wPort_1_banks_0 = x823_x726_D67_number[2:0]; // @[MemInterfaceType.scala 88:58:@63089.4]
  assign x384_lb2_0_io_wPort_1_ofs_0 = x825_x399_sum_D45_number[8:0]; // @[MemInterfaceType.scala 89:54:@63091.4]
  assign x384_lb2_0_io_wPort_1_data_0 = RetimeWrapper_117_io_out; // @[MemInterfaceType.scala 90:56:@63092.4]
  assign x384_lb2_0_io_wPort_1_en_0 = _T_1820 & x820_b380_D67; // @[MemInterfaceType.scala 93:57:@63094.4]
  assign x384_lb2_0_io_wPort_0_banks_1 = x819_x389_D51_number[2:0]; // @[MemInterfaceType.scala 88:58:@63040.4]
  assign x384_lb2_0_io_wPort_0_banks_0 = x823_x726_D67_number[2:0]; // @[MemInterfaceType.scala 88:58:@63039.4]
  assign x384_lb2_0_io_wPort_0_ofs_0 = x822_x393_sum_D46_number[8:0]; // @[MemInterfaceType.scala 89:54:@63041.4]
  assign x384_lb2_0_io_wPort_0_data_0 = RetimeWrapper_111_io_out; // @[MemInterfaceType.scala 90:56:@63042.4]
  assign x384_lb2_0_io_wPort_0_en_0 = _T_1797 & x820_b380_D67; // @[MemInterfaceType.scala 93:57:@63044.4]
  assign x389_1_clock = clock; // @[:@60153.4]
  assign x389_1_io_a = __1_io_result; // @[Math.scala 367:17:@60155.4]
  assign x389_1_io_flow = io_in_x343_TREADY; // @[Math.scala 369:20:@60157.4]
  assign x729_sum_1_clock = clock; // @[:@60190.4]
  assign x729_sum_1_reset = reset; // @[:@60191.4]
  assign x729_sum_1_io_a = _T_301[31:0]; // @[Math.scala 151:17:@60192.4]
  assign x729_sum_1_io_b = _T_304[31:0]; // @[Math.scala 152:17:@60193.4]
  assign x729_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60194.4]
  assign x392_div_1_clock = clock; // @[:@60202.4]
  assign x392_div_1_io_a = __1_io_result; // @[Math.scala 328:17:@60204.4]
  assign x392_div_1_io_flow = io_in_x343_TREADY; // @[Math.scala 330:20:@60206.4]
  assign RetimeWrapper_1_clock = clock; // @[:@60212.4]
  assign RetimeWrapper_1_reset = reset; // @[:@60213.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60215.4]
  assign RetimeWrapper_1_io_in = x729_sum_1_io_result; // @[package.scala 94:16:@60214.4]
  assign x393_sum_1_clock = clock; // @[:@60221.4]
  assign x393_sum_1_reset = reset; // @[:@60222.4]
  assign x393_sum_1_io_a = RetimeWrapper_1_io_out; // @[Math.scala 151:17:@60223.4]
  assign x393_sum_1_io_b = x392_div_1_io_result; // @[Math.scala 152:17:@60224.4]
  assign x393_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60225.4]
  assign RetimeWrapper_2_clock = clock; // @[:@60231.4]
  assign RetimeWrapper_2_reset = reset; // @[:@60232.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60234.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@60233.4]
  assign RetimeWrapper_3_clock = clock; // @[:@60240.4]
  assign RetimeWrapper_3_reset = reset; // @[:@60241.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60243.4]
  assign RetimeWrapper_3_io_in = x389_1_io_result; // @[package.scala 94:16:@60242.4]
  assign RetimeWrapper_4_clock = clock; // @[:@60249.4]
  assign RetimeWrapper_4_reset = reset; // @[:@60250.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60252.4]
  assign RetimeWrapper_4_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@60251.4]
  assign RetimeWrapper_5_clock = clock; // @[:@60258.4]
  assign RetimeWrapper_5_reset = reset; // @[:@60259.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60261.4]
  assign RetimeWrapper_5_io_in = x393_sum_1_io_result; // @[package.scala 94:16:@60260.4]
  assign RetimeWrapper_6_clock = clock; // @[:@60267.4]
  assign RetimeWrapper_6_reset = reset; // @[:@60268.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60270.4]
  assign RetimeWrapper_6_io_in = x745_x381_D1_0_number[31:0]; // @[package.scala 94:16:@60269.4]
  assign RetimeWrapper_7_clock = clock; // @[:@60276.4]
  assign RetimeWrapper_7_reset = reset; // @[:@60277.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60279.4]
  assign RetimeWrapper_7_io_in = $unsigned(_T_264); // @[package.scala 94:16:@60278.4]
  assign RetimeWrapper_8_clock = clock; // @[:@60287.4]
  assign RetimeWrapper_8_reset = reset; // @[:@60288.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60290.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60289.4]
  assign x395_rdcol_1_clock = clock; // @[:@60310.4]
  assign x395_rdcol_1_reset = reset; // @[:@60311.4]
  assign x395_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@60312.4]
  assign x395_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@60313.4]
  assign x395_rdcol_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60314.4]
  assign x397_1_clock = clock; // @[:@60324.4]
  assign x397_1_io_a = x395_rdcol_1_io_result; // @[Math.scala 367:17:@60326.4]
  assign x397_1_io_flow = io_in_x343_TREADY; // @[Math.scala 369:20:@60328.4]
  assign x398_div_1_clock = clock; // @[:@60336.4]
  assign x398_div_1_io_a = x395_rdcol_1_io_result; // @[Math.scala 328:17:@60338.4]
  assign x398_div_1_io_flow = io_in_x343_TREADY; // @[Math.scala 330:20:@60340.4]
  assign RetimeWrapper_9_clock = clock; // @[:@60346.4]
  assign RetimeWrapper_9_reset = reset; // @[:@60347.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60349.4]
  assign RetimeWrapper_9_io_in = x729_sum_1_io_result; // @[package.scala 94:16:@60348.4]
  assign x399_sum_1_clock = clock; // @[:@60355.4]
  assign x399_sum_1_reset = reset; // @[:@60356.4]
  assign x399_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@60357.4]
  assign x399_sum_1_io_b = x398_div_1_io_result; // @[Math.scala 152:17:@60358.4]
  assign x399_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60359.4]
  assign RetimeWrapper_10_clock = clock; // @[:@60365.4]
  assign RetimeWrapper_10_reset = reset; // @[:@60366.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60368.4]
  assign RetimeWrapper_10_io_in = x397_1_io_result; // @[package.scala 94:16:@60367.4]
  assign RetimeWrapper_11_clock = clock; // @[:@60374.4]
  assign RetimeWrapper_11_reset = reset; // @[:@60375.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60377.4]
  assign RetimeWrapper_11_io_in = x745_x381_D1_0_number[63:32]; // @[package.scala 94:16:@60376.4]
  assign RetimeWrapper_12_clock = clock; // @[:@60383.4]
  assign RetimeWrapper_12_reset = reset; // @[:@60384.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60386.4]
  assign RetimeWrapper_12_io_in = x399_sum_1_io_result; // @[package.scala 94:16:@60385.4]
  assign RetimeWrapper_13_clock = clock; // @[:@60394.4]
  assign RetimeWrapper_13_reset = reset; // @[:@60395.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60397.4]
  assign RetimeWrapper_13_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60396.4]
  assign x401_rdcol_1_clock = clock; // @[:@60417.4]
  assign x401_rdcol_1_reset = reset; // @[:@60418.4]
  assign x401_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@60419.4]
  assign x401_rdcol_1_io_b = 32'h2; // @[Math.scala 152:17:@60420.4]
  assign x401_rdcol_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60421.4]
  assign x403_1_clock = clock; // @[:@60431.4]
  assign x403_1_io_a = x401_rdcol_1_io_result; // @[Math.scala 367:17:@60433.4]
  assign x403_1_io_flow = io_in_x343_TREADY; // @[Math.scala 369:20:@60435.4]
  assign x404_div_1_clock = clock; // @[:@60443.4]
  assign x404_div_1_io_a = x401_rdcol_1_io_result; // @[Math.scala 328:17:@60445.4]
  assign x404_div_1_io_flow = io_in_x343_TREADY; // @[Math.scala 330:20:@60447.4]
  assign x405_sum_1_clock = clock; // @[:@60453.4]
  assign x405_sum_1_reset = reset; // @[:@60454.4]
  assign x405_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@60455.4]
  assign x405_sum_1_io_b = x404_div_1_io_result; // @[Math.scala 152:17:@60456.4]
  assign x405_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60457.4]
  assign RetimeWrapper_14_clock = clock; // @[:@60463.4]
  assign RetimeWrapper_14_reset = reset; // @[:@60464.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60466.4]
  assign RetimeWrapper_14_io_in = x403_1_io_result; // @[package.scala 94:16:@60465.4]
  assign RetimeWrapper_15_clock = clock; // @[:@60472.4]
  assign RetimeWrapper_15_reset = reset; // @[:@60473.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60475.4]
  assign RetimeWrapper_15_io_in = x745_x381_D1_0_number[95:64]; // @[package.scala 94:16:@60474.4]
  assign RetimeWrapper_16_clock = clock; // @[:@60481.4]
  assign RetimeWrapper_16_reset = reset; // @[:@60482.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60484.4]
  assign RetimeWrapper_16_io_in = x405_sum_1_io_result; // @[package.scala 94:16:@60483.4]
  assign RetimeWrapper_17_clock = clock; // @[:@60492.4]
  assign RetimeWrapper_17_reset = reset; // @[:@60493.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60495.4]
  assign RetimeWrapper_17_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60494.4]
  assign x407_rdcol_1_clock = clock; // @[:@60515.4]
  assign x407_rdcol_1_reset = reset; // @[:@60516.4]
  assign x407_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@60517.4]
  assign x407_rdcol_1_io_b = 32'h3; // @[Math.scala 152:17:@60518.4]
  assign x407_rdcol_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60519.4]
  assign x409_1_clock = clock; // @[:@60529.4]
  assign x409_1_io_a = x407_rdcol_1_io_result; // @[Math.scala 367:17:@60531.4]
  assign x409_1_io_flow = io_in_x343_TREADY; // @[Math.scala 369:20:@60533.4]
  assign x410_div_1_clock = clock; // @[:@60541.4]
  assign x410_div_1_io_a = x407_rdcol_1_io_result; // @[Math.scala 328:17:@60543.4]
  assign x410_div_1_io_flow = io_in_x343_TREADY; // @[Math.scala 330:20:@60545.4]
  assign x411_sum_1_clock = clock; // @[:@60551.4]
  assign x411_sum_1_reset = reset; // @[:@60552.4]
  assign x411_sum_1_io_a = RetimeWrapper_9_io_out; // @[Math.scala 151:17:@60553.4]
  assign x411_sum_1_io_b = x410_div_1_io_result; // @[Math.scala 152:17:@60554.4]
  assign x411_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60555.4]
  assign RetimeWrapper_18_clock = clock; // @[:@60561.4]
  assign RetimeWrapper_18_reset = reset; // @[:@60562.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60564.4]
  assign RetimeWrapper_18_io_in = x745_x381_D1_0_number[127:96]; // @[package.scala 94:16:@60563.4]
  assign RetimeWrapper_19_clock = clock; // @[:@60570.4]
  assign RetimeWrapper_19_reset = reset; // @[:@60571.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60573.4]
  assign RetimeWrapper_19_io_in = x411_sum_1_io_result; // @[package.scala 94:16:@60572.4]
  assign RetimeWrapper_20_clock = clock; // @[:@60579.4]
  assign RetimeWrapper_20_reset = reset; // @[:@60580.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60582.4]
  assign RetimeWrapper_20_io_in = x409_1_io_result; // @[package.scala 94:16:@60581.4]
  assign RetimeWrapper_21_clock = clock; // @[:@60590.4]
  assign RetimeWrapper_21_reset = reset; // @[:@60591.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60593.4]
  assign RetimeWrapper_21_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60592.4]
  assign RetimeWrapper_22_clock = clock; // @[:@60611.4]
  assign RetimeWrapper_22_reset = reset; // @[:@60612.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60614.4]
  assign RetimeWrapper_22_io_in = __io_result; // @[package.scala 94:16:@60613.4]
  assign RetimeWrapper_23_clock = clock; // @[:@60627.4]
  assign RetimeWrapper_23_reset = reset; // @[:@60628.4]
  assign RetimeWrapper_23_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@60630.4]
  assign RetimeWrapper_23_io_in = $signed(_T_510) < $signed(32'sh0); // @[package.scala 94:16:@60629.4]
  assign RetimeWrapper_24_clock = clock; // @[:@60636.4]
  assign RetimeWrapper_24_reset = reset; // @[:@60637.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60639.4]
  assign RetimeWrapper_24_io_in = x407_rdcol_1_io_result; // @[package.scala 94:16:@60638.4]
  assign RetimeWrapper_25_clock = clock; // @[:@60650.4]
  assign RetimeWrapper_25_reset = reset; // @[:@60651.4]
  assign RetimeWrapper_25_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@60653.4]
  assign RetimeWrapper_25_io_in = $signed(_T_523) < $signed(32'sh0); // @[package.scala 94:16:@60652.4]
  assign RetimeWrapper_26_clock = clock; // @[:@60659.4]
  assign RetimeWrapper_26_reset = reset; // @[:@60660.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60662.4]
  assign RetimeWrapper_26_io_in = RetimeWrapper_23_io_out; // @[package.scala 94:16:@60661.4]
  assign RetimeWrapper_27_clock = clock; // @[:@60674.4]
  assign RetimeWrapper_27_reset = reset; // @[:@60675.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60677.4]
  assign RetimeWrapper_27_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@60676.4]
  assign RetimeWrapper_28_clock = clock; // @[:@60683.4]
  assign RetimeWrapper_28_reset = reset; // @[:@60684.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60686.4]
  assign RetimeWrapper_28_io_in = ~ x416; // @[package.scala 94:16:@60685.4]
  assign RetimeWrapper_29_clock = clock; // @[:@60692.4]
  assign RetimeWrapper_29_reset = reset; // @[:@60693.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60695.4]
  assign RetimeWrapper_29_io_in = x411_sum_1_io_result; // @[package.scala 94:16:@60694.4]
  assign RetimeWrapper_30_clock = clock; // @[:@60701.4]
  assign RetimeWrapper_30_reset = reset; // @[:@60702.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60704.4]
  assign RetimeWrapper_30_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@60703.4]
  assign RetimeWrapper_31_clock = clock; // @[:@60710.4]
  assign RetimeWrapper_31_reset = reset; // @[:@60711.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60713.4]
  assign RetimeWrapper_31_io_in = $unsigned(_T_264); // @[package.scala 94:16:@60712.4]
  assign RetimeWrapper_32_clock = clock; // @[:@60719.4]
  assign RetimeWrapper_32_reset = reset; // @[:@60720.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60722.4]
  assign RetimeWrapper_32_io_in = x409_1_io_result; // @[package.scala 94:16:@60721.4]
  assign RetimeWrapper_33_clock = clock; // @[:@60731.4]
  assign RetimeWrapper_33_reset = reset; // @[:@60732.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60734.4]
  assign RetimeWrapper_33_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60733.4]
  assign RetimeWrapper_34_clock = clock; // @[:@60752.4]
  assign RetimeWrapper_34_reset = reset; // @[:@60753.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60755.4]
  assign RetimeWrapper_34_io_in = x401_rdcol_1_io_result; // @[package.scala 94:16:@60754.4]
  assign RetimeWrapper_35_clock = clock; // @[:@60766.4]
  assign RetimeWrapper_35_reset = reset; // @[:@60767.4]
  assign RetimeWrapper_35_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@60769.4]
  assign RetimeWrapper_35_io_in = $signed(_T_580) < $signed(32'sh0); // @[package.scala 94:16:@60768.4]
  assign RetimeWrapper_36_clock = clock; // @[:@60781.4]
  assign RetimeWrapper_36_reset = reset; // @[:@60782.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60784.4]
  assign RetimeWrapper_36_io_in = x403_1_io_result; // @[package.scala 94:16:@60783.4]
  assign RetimeWrapper_37_clock = clock; // @[:@60790.4]
  assign RetimeWrapper_37_reset = reset; // @[:@60791.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60793.4]
  assign RetimeWrapper_37_io_in = x405_sum_1_io_result; // @[package.scala 94:16:@60792.4]
  assign RetimeWrapper_38_clock = clock; // @[:@60799.4]
  assign RetimeWrapper_38_reset = reset; // @[:@60800.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60802.4]
  assign RetimeWrapper_38_io_in = ~ x421; // @[package.scala 94:16:@60801.4]
  assign RetimeWrapper_39_clock = clock; // @[:@60811.4]
  assign RetimeWrapper_39_reset = reset; // @[:@60812.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60814.4]
  assign RetimeWrapper_39_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60813.4]
  assign RetimeWrapper_40_clock = clock; // @[:@60832.4]
  assign RetimeWrapper_40_reset = reset; // @[:@60833.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60835.4]
  assign RetimeWrapper_40_io_in = x395_rdcol_1_io_result; // @[package.scala 94:16:@60834.4]
  assign RetimeWrapper_41_clock = clock; // @[:@60846.4]
  assign RetimeWrapper_41_reset = reset; // @[:@60847.4]
  assign RetimeWrapper_41_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@60849.4]
  assign RetimeWrapper_41_io_in = $signed(_T_625) < $signed(32'sh0); // @[package.scala 94:16:@60848.4]
  assign RetimeWrapper_42_clock = clock; // @[:@60861.4]
  assign RetimeWrapper_42_reset = reset; // @[:@60862.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60864.4]
  assign RetimeWrapper_42_io_in = x397_1_io_result; // @[package.scala 94:16:@60863.4]
  assign RetimeWrapper_43_clock = clock; // @[:@60870.4]
  assign RetimeWrapper_43_reset = reset; // @[:@60871.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60873.4]
  assign RetimeWrapper_43_io_in = x399_sum_1_io_result; // @[package.scala 94:16:@60872.4]
  assign RetimeWrapper_44_clock = clock; // @[:@60879.4]
  assign RetimeWrapper_44_reset = reset; // @[:@60880.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60882.4]
  assign RetimeWrapper_44_io_in = ~ x426; // @[package.scala 94:16:@60881.4]
  assign RetimeWrapper_45_clock = clock; // @[:@60891.4]
  assign RetimeWrapper_45_reset = reset; // @[:@60892.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60894.4]
  assign RetimeWrapper_45_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60893.4]
  assign RetimeWrapper_46_clock = clock; // @[:@60912.4]
  assign RetimeWrapper_46_reset = reset; // @[:@60913.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60915.4]
  assign RetimeWrapper_46_io_in = __1_io_result; // @[package.scala 94:16:@60914.4]
  assign RetimeWrapper_47_clock = clock; // @[:@60926.4]
  assign RetimeWrapper_47_reset = reset; // @[:@60927.4]
  assign RetimeWrapper_47_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@60929.4]
  assign RetimeWrapper_47_io_in = $signed(_T_670) < $signed(32'sh0); // @[package.scala 94:16:@60928.4]
  assign RetimeWrapper_48_clock = clock; // @[:@60941.4]
  assign RetimeWrapper_48_reset = reset; // @[:@60942.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60944.4]
  assign RetimeWrapper_48_io_in = x389_1_io_result; // @[package.scala 94:16:@60943.4]
  assign RetimeWrapper_49_clock = clock; // @[:@60950.4]
  assign RetimeWrapper_49_reset = reset; // @[:@60951.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60953.4]
  assign RetimeWrapper_49_io_in = x393_sum_1_io_result; // @[package.scala 94:16:@60952.4]
  assign RetimeWrapper_50_clock = clock; // @[:@60959.4]
  assign RetimeWrapper_50_reset = reset; // @[:@60960.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60962.4]
  assign RetimeWrapper_50_io_in = ~ x431; // @[package.scala 94:16:@60961.4]
  assign RetimeWrapper_51_clock = clock; // @[:@60971.4]
  assign RetimeWrapper_51_reset = reset; // @[:@60972.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@60974.4]
  assign RetimeWrapper_51_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@60973.4]
  assign x435_rdcol_1_clock = clock; // @[:@60994.4]
  assign x435_rdcol_1_reset = reset; // @[:@60995.4]
  assign x435_rdcol_1_io_a = RetimeWrapper_46_io_out; // @[Math.scala 151:17:@60996.4]
  assign x435_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@60997.4]
  assign x435_rdcol_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@60998.4]
  assign RetimeWrapper_52_clock = clock; // @[:@61009.4]
  assign RetimeWrapper_52_reset = reset; // @[:@61010.4]
  assign RetimeWrapper_52_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@61012.4]
  assign RetimeWrapper_52_io_in = $signed(_T_719) < $signed(32'sh0); // @[package.scala 94:16:@61011.4]
  assign x439_1_clock = clock; // @[:@61028.4]
  assign x439_1_io_a = x435_rdcol_1_io_result; // @[Math.scala 367:17:@61030.4]
  assign x439_1_io_flow = io_in_x343_TREADY; // @[Math.scala 369:20:@61032.4]
  assign x440_div_1_clock = clock; // @[:@61040.4]
  assign x440_div_1_io_a = x435_rdcol_1_io_result; // @[Math.scala 328:17:@61042.4]
  assign x440_div_1_io_flow = io_in_x343_TREADY; // @[Math.scala 330:20:@61044.4]
  assign RetimeWrapper_53_clock = clock; // @[:@61050.4]
  assign RetimeWrapper_53_reset = reset; // @[:@61051.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61053.4]
  assign RetimeWrapper_53_io_in = x729_sum_1_io_result; // @[package.scala 94:16:@61052.4]
  assign x441_sum_1_clock = clock; // @[:@61059.4]
  assign x441_sum_1_reset = reset; // @[:@61060.4]
  assign x441_sum_1_io_a = RetimeWrapper_53_io_out; // @[Math.scala 151:17:@61061.4]
  assign x441_sum_1_io_b = x440_div_1_io_result; // @[Math.scala 152:17:@61062.4]
  assign x441_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61063.4]
  assign RetimeWrapper_54_clock = clock; // @[:@61069.4]
  assign RetimeWrapper_54_reset = reset; // @[:@61070.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61072.4]
  assign RetimeWrapper_54_io_in = x439_1_io_result; // @[package.scala 94:16:@61071.4]
  assign RetimeWrapper_55_clock = clock; // @[:@61078.4]
  assign RetimeWrapper_55_reset = reset; // @[:@61079.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61081.4]
  assign RetimeWrapper_55_io_in = ~ x437; // @[package.scala 94:16:@61080.4]
  assign RetimeWrapper_56_clock = clock; // @[:@61090.4]
  assign RetimeWrapper_56_reset = reset; // @[:@61091.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61093.4]
  assign RetimeWrapper_56_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61092.4]
  assign x444_rdcol_1_clock = clock; // @[:@61113.4]
  assign x444_rdcol_1_reset = reset; // @[:@61114.4]
  assign x444_rdcol_1_io_a = RetimeWrapper_46_io_out; // @[Math.scala 151:17:@61115.4]
  assign x444_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@61116.4]
  assign x444_rdcol_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61117.4]
  assign RetimeWrapper_57_clock = clock; // @[:@61128.4]
  assign RetimeWrapper_57_reset = reset; // @[:@61129.4]
  assign RetimeWrapper_57_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@61131.4]
  assign RetimeWrapper_57_io_in = $signed(_T_787) < $signed(32'sh0); // @[package.scala 94:16:@61130.4]
  assign x448_1_clock = clock; // @[:@61145.4]
  assign x448_1_io_a = x444_rdcol_1_io_result; // @[Math.scala 367:17:@61147.4]
  assign x448_1_io_flow = io_in_x343_TREADY; // @[Math.scala 369:20:@61149.4]
  assign x449_div_1_clock = clock; // @[:@61157.4]
  assign x449_div_1_io_a = x444_rdcol_1_io_result; // @[Math.scala 328:17:@61159.4]
  assign x449_div_1_io_flow = io_in_x343_TREADY; // @[Math.scala 330:20:@61161.4]
  assign x450_sum_1_clock = clock; // @[:@61167.4]
  assign x450_sum_1_reset = reset; // @[:@61168.4]
  assign x450_sum_1_io_a = RetimeWrapper_53_io_out; // @[Math.scala 151:17:@61169.4]
  assign x450_sum_1_io_b = x449_div_1_io_result; // @[Math.scala 152:17:@61170.4]
  assign x450_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61171.4]
  assign RetimeWrapper_58_clock = clock; // @[:@61177.4]
  assign RetimeWrapper_58_reset = reset; // @[:@61178.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61180.4]
  assign RetimeWrapper_58_io_in = x448_1_io_result; // @[package.scala 94:16:@61179.4]
  assign RetimeWrapper_59_clock = clock; // @[:@61186.4]
  assign RetimeWrapper_59_reset = reset; // @[:@61187.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61189.4]
  assign RetimeWrapper_59_io_in = ~ x446; // @[package.scala 94:16:@61188.4]
  assign RetimeWrapper_60_clock = clock; // @[:@61198.4]
  assign RetimeWrapper_60_reset = reset; // @[:@61199.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61201.4]
  assign RetimeWrapper_60_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61200.4]
  assign x453_rdrow_1_clock = clock; // @[:@61221.4]
  assign x453_rdrow_1_reset = reset; // @[:@61222.4]
  assign x453_rdrow_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 192:17:@61223.4]
  assign x453_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@61224.4]
  assign x453_rdrow_1_io_flow = io_in_x343_TREADY; // @[Math.scala 194:20:@61225.4]
  assign RetimeWrapper_61_clock = clock; // @[:@61247.4]
  assign RetimeWrapper_61_reset = reset; // @[:@61248.4]
  assign RetimeWrapper_61_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@61250.4]
  assign RetimeWrapper_61_io_in = $signed(_T_852) < $signed(32'sh0); // @[package.scala 94:16:@61249.4]
  assign RetimeWrapper_62_clock = clock; // @[:@61269.4]
  assign RetimeWrapper_62_reset = reset; // @[:@61270.4]
  assign RetimeWrapper_62_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@61273.4]
  assign RetimeWrapper_62_io_in = $unsigned(_T_881); // @[package.scala 94:16:@61272.4]
  assign RetimeWrapper_63_clock = clock; // @[:@61295.4]
  assign RetimeWrapper_63_reset = reset; // @[:@61296.4]
  assign RetimeWrapper_63_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@61298.4]
  assign RetimeWrapper_63_io_in = {_T_893,_T_894}; // @[package.scala 94:16:@61297.4]
  assign x734_sum_1_clock = clock; // @[:@61316.4]
  assign x734_sum_1_reset = reset; // @[:@61317.4]
  assign x734_sum_1_io_a = _T_917[31:0]; // @[Math.scala 151:17:@61318.4]
  assign x734_sum_1_io_b = _T_920[31:0]; // @[Math.scala 152:17:@61319.4]
  assign x734_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61320.4]
  assign RetimeWrapper_64_clock = clock; // @[:@61326.4]
  assign RetimeWrapper_64_reset = reset; // @[:@61327.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61329.4]
  assign RetimeWrapper_64_io_in = x410_div_1_io_result; // @[package.scala 94:16:@61328.4]
  assign RetimeWrapper_65_clock = clock; // @[:@61335.4]
  assign RetimeWrapper_65_reset = reset; // @[:@61336.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61338.4]
  assign RetimeWrapper_65_io_in = x734_sum_1_io_result; // @[package.scala 94:16:@61337.4]
  assign x461_sum_1_clock = clock; // @[:@61344.4]
  assign x461_sum_1_reset = reset; // @[:@61345.4]
  assign x461_sum_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@61346.4]
  assign x461_sum_1_io_b = RetimeWrapper_64_io_out; // @[Math.scala 152:17:@61347.4]
  assign x461_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61348.4]
  assign RetimeWrapper_66_clock = clock; // @[:@61354.4]
  assign RetimeWrapper_66_reset = reset; // @[:@61355.4]
  assign RetimeWrapper_66_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61357.4]
  assign RetimeWrapper_66_io_in = ~ x456; // @[package.scala 94:16:@61356.4]
  assign RetimeWrapper_67_clock = clock; // @[:@61363.4]
  assign RetimeWrapper_67_reset = reset; // @[:@61364.4]
  assign RetimeWrapper_67_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61366.4]
  assign RetimeWrapper_67_io_in = $unsigned(_T_885); // @[package.scala 94:16:@61365.4]
  assign RetimeWrapper_68_clock = clock; // @[:@61375.4]
  assign RetimeWrapper_68_reset = reset; // @[:@61376.4]
  assign RetimeWrapper_68_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61378.4]
  assign RetimeWrapper_68_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61377.4]
  assign RetimeWrapper_69_clock = clock; // @[:@61402.4]
  assign RetimeWrapper_69_reset = reset; // @[:@61403.4]
  assign RetimeWrapper_69_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61405.4]
  assign RetimeWrapper_69_io_in = x404_div_1_io_result; // @[package.scala 94:16:@61404.4]
  assign x466_sum_1_clock = clock; // @[:@61411.4]
  assign x466_sum_1_reset = reset; // @[:@61412.4]
  assign x466_sum_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@61413.4]
  assign x466_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@61414.4]
  assign x466_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61415.4]
  assign RetimeWrapper_70_clock = clock; // @[:@61421.4]
  assign RetimeWrapper_70_reset = reset; // @[:@61422.4]
  assign RetimeWrapper_70_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61424.4]
  assign RetimeWrapper_70_io_in = ~ x464; // @[package.scala 94:16:@61423.4]
  assign RetimeWrapper_71_clock = clock; // @[:@61433.4]
  assign RetimeWrapper_71_reset = reset; // @[:@61434.4]
  assign RetimeWrapper_71_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61436.4]
  assign RetimeWrapper_71_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61435.4]
  assign RetimeWrapper_72_clock = clock; // @[:@61460.4]
  assign RetimeWrapper_72_reset = reset; // @[:@61461.4]
  assign RetimeWrapper_72_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61463.4]
  assign RetimeWrapper_72_io_in = x398_div_1_io_result; // @[package.scala 94:16:@61462.4]
  assign x471_sum_1_clock = clock; // @[:@61469.4]
  assign x471_sum_1_reset = reset; // @[:@61470.4]
  assign x471_sum_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@61471.4]
  assign x471_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@61472.4]
  assign x471_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61473.4]
  assign RetimeWrapper_73_clock = clock; // @[:@61479.4]
  assign RetimeWrapper_73_reset = reset; // @[:@61480.4]
  assign RetimeWrapper_73_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61482.4]
  assign RetimeWrapper_73_io_in = ~ x469; // @[package.scala 94:16:@61481.4]
  assign RetimeWrapper_74_clock = clock; // @[:@61491.4]
  assign RetimeWrapper_74_reset = reset; // @[:@61492.4]
  assign RetimeWrapper_74_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61494.4]
  assign RetimeWrapper_74_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61493.4]
  assign RetimeWrapper_75_clock = clock; // @[:@61512.4]
  assign RetimeWrapper_75_reset = reset; // @[:@61513.4]
  assign RetimeWrapper_75_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61515.4]
  assign RetimeWrapper_75_io_in = RetimeWrapper_47_io_out; // @[package.scala 94:16:@61514.4]
  assign RetimeWrapper_76_clock = clock; // @[:@61527.4]
  assign RetimeWrapper_76_reset = reset; // @[:@61528.4]
  assign RetimeWrapper_76_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61530.4]
  assign RetimeWrapper_76_io_in = x392_div_1_io_result; // @[package.scala 94:16:@61529.4]
  assign RetimeWrapper_77_clock = clock; // @[:@61536.4]
  assign RetimeWrapper_77_reset = reset; // @[:@61537.4]
  assign RetimeWrapper_77_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61539.4]
  assign RetimeWrapper_77_io_in = x734_sum_1_io_result; // @[package.scala 94:16:@61538.4]
  assign x476_sum_1_clock = clock; // @[:@61547.4]
  assign x476_sum_1_reset = reset; // @[:@61548.4]
  assign x476_sum_1_io_a = RetimeWrapper_77_io_out; // @[Math.scala 151:17:@61549.4]
  assign x476_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@61550.4]
  assign x476_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61551.4]
  assign RetimeWrapper_78_clock = clock; // @[:@61557.4]
  assign RetimeWrapper_78_reset = reset; // @[:@61558.4]
  assign RetimeWrapper_78_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61560.4]
  assign RetimeWrapper_78_io_in = ~ x474; // @[package.scala 94:16:@61559.4]
  assign RetimeWrapper_79_clock = clock; // @[:@61566.4]
  assign RetimeWrapper_79_reset = reset; // @[:@61567.4]
  assign RetimeWrapper_79_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61569.4]
  assign RetimeWrapper_79_io_in = x476_sum_1_io_result; // @[package.scala 94:16:@61568.4]
  assign RetimeWrapper_80_clock = clock; // @[:@61578.4]
  assign RetimeWrapper_80_reset = reset; // @[:@61579.4]
  assign RetimeWrapper_80_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61581.4]
  assign RetimeWrapper_80_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61580.4]
  assign x481_sum_1_clock = clock; // @[:@61605.4]
  assign x481_sum_1_reset = reset; // @[:@61606.4]
  assign x481_sum_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@61607.4]
  assign x481_sum_1_io_b = x440_div_1_io_result; // @[Math.scala 152:17:@61608.4]
  assign x481_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61609.4]
  assign RetimeWrapper_81_clock = clock; // @[:@61615.4]
  assign RetimeWrapper_81_reset = reset; // @[:@61616.4]
  assign RetimeWrapper_81_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61618.4]
  assign RetimeWrapper_81_io_in = ~ x479; // @[package.scala 94:16:@61617.4]
  assign RetimeWrapper_82_clock = clock; // @[:@61627.4]
  assign RetimeWrapper_82_reset = reset; // @[:@61628.4]
  assign RetimeWrapper_82_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61630.4]
  assign RetimeWrapper_82_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61629.4]
  assign x486_sum_1_clock = clock; // @[:@61654.4]
  assign x486_sum_1_reset = reset; // @[:@61655.4]
  assign x486_sum_1_io_a = RetimeWrapper_65_io_out; // @[Math.scala 151:17:@61656.4]
  assign x486_sum_1_io_b = x449_div_1_io_result; // @[Math.scala 152:17:@61657.4]
  assign x486_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61658.4]
  assign RetimeWrapper_83_clock = clock; // @[:@61664.4]
  assign RetimeWrapper_83_reset = reset; // @[:@61665.4]
  assign RetimeWrapper_83_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61667.4]
  assign RetimeWrapper_83_io_in = ~ x484; // @[package.scala 94:16:@61666.4]
  assign RetimeWrapper_84_clock = clock; // @[:@61676.4]
  assign RetimeWrapper_84_reset = reset; // @[:@61677.4]
  assign RetimeWrapper_84_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61679.4]
  assign RetimeWrapper_84_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61678.4]
  assign x489_rdrow_1_clock = clock; // @[:@61699.4]
  assign x489_rdrow_1_reset = reset; // @[:@61700.4]
  assign x489_rdrow_1_io_a = RetimeWrapper_22_io_out; // @[Math.scala 192:17:@61701.4]
  assign x489_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@61702.4]
  assign x489_rdrow_1_io_flow = io_in_x343_TREADY; // @[Math.scala 194:20:@61703.4]
  assign RetimeWrapper_85_clock = clock; // @[:@61725.4]
  assign RetimeWrapper_85_reset = reset; // @[:@61726.4]
  assign RetimeWrapper_85_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@61728.4]
  assign RetimeWrapper_85_io_in = $signed(_T_1137) < $signed(32'sh0); // @[package.scala 94:16:@61727.4]
  assign RetimeWrapper_86_clock = clock; // @[:@61747.4]
  assign RetimeWrapper_86_reset = reset; // @[:@61748.4]
  assign RetimeWrapper_86_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@61751.4]
  assign RetimeWrapper_86_io_in = $unsigned(_T_1166); // @[package.scala 94:16:@61750.4]
  assign RetimeWrapper_87_clock = clock; // @[:@61773.4]
  assign RetimeWrapper_87_reset = reset; // @[:@61774.4]
  assign RetimeWrapper_87_io_flow = io_in_x343_TREADY; // @[package.scala 95:18:@61776.4]
  assign RetimeWrapper_87_io_in = {_T_1178,_T_1179}; // @[package.scala 94:16:@61775.4]
  assign x739_sum_1_clock = clock; // @[:@61794.4]
  assign x739_sum_1_reset = reset; // @[:@61795.4]
  assign x739_sum_1_io_a = _T_1202[31:0]; // @[Math.scala 151:17:@61796.4]
  assign x739_sum_1_io_b = _T_1205[31:0]; // @[Math.scala 152:17:@61797.4]
  assign x739_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61798.4]
  assign RetimeWrapper_88_clock = clock; // @[:@61804.4]
  assign RetimeWrapper_88_reset = reset; // @[:@61805.4]
  assign RetimeWrapper_88_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61807.4]
  assign RetimeWrapper_88_io_in = x739_sum_1_io_result; // @[package.scala 94:16:@61806.4]
  assign x497_sum_1_clock = clock; // @[:@61813.4]
  assign x497_sum_1_reset = reset; // @[:@61814.4]
  assign x497_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@61815.4]
  assign x497_sum_1_io_b = RetimeWrapper_64_io_out; // @[Math.scala 152:17:@61816.4]
  assign x497_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61817.4]
  assign RetimeWrapper_89_clock = clock; // @[:@61823.4]
  assign RetimeWrapper_89_reset = reset; // @[:@61824.4]
  assign RetimeWrapper_89_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61826.4]
  assign RetimeWrapper_89_io_in = ~ x492; // @[package.scala 94:16:@61825.4]
  assign RetimeWrapper_90_clock = clock; // @[:@61832.4]
  assign RetimeWrapper_90_reset = reset; // @[:@61833.4]
  assign RetimeWrapper_90_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61835.4]
  assign RetimeWrapper_90_io_in = $unsigned(_T_1170); // @[package.scala 94:16:@61834.4]
  assign RetimeWrapper_91_clock = clock; // @[:@61844.4]
  assign RetimeWrapper_91_reset = reset; // @[:@61845.4]
  assign RetimeWrapper_91_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61847.4]
  assign RetimeWrapper_91_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61846.4]
  assign x502_sum_1_clock = clock; // @[:@61871.4]
  assign x502_sum_1_reset = reset; // @[:@61872.4]
  assign x502_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@61873.4]
  assign x502_sum_1_io_b = RetimeWrapper_69_io_out; // @[Math.scala 152:17:@61874.4]
  assign x502_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61875.4]
  assign RetimeWrapper_92_clock = clock; // @[:@61881.4]
  assign RetimeWrapper_92_reset = reset; // @[:@61882.4]
  assign RetimeWrapper_92_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61884.4]
  assign RetimeWrapper_92_io_in = ~ x500; // @[package.scala 94:16:@61883.4]
  assign RetimeWrapper_93_clock = clock; // @[:@61893.4]
  assign RetimeWrapper_93_reset = reset; // @[:@61894.4]
  assign RetimeWrapper_93_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61896.4]
  assign RetimeWrapper_93_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61895.4]
  assign x507_sum_1_clock = clock; // @[:@61920.4]
  assign x507_sum_1_reset = reset; // @[:@61921.4]
  assign x507_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@61922.4]
  assign x507_sum_1_io_b = RetimeWrapper_72_io_out; // @[Math.scala 152:17:@61923.4]
  assign x507_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61924.4]
  assign RetimeWrapper_94_clock = clock; // @[:@61930.4]
  assign RetimeWrapper_94_reset = reset; // @[:@61931.4]
  assign RetimeWrapper_94_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61933.4]
  assign RetimeWrapper_94_io_in = ~ x505; // @[package.scala 94:16:@61932.4]
  assign RetimeWrapper_95_clock = clock; // @[:@61942.4]
  assign RetimeWrapper_95_reset = reset; // @[:@61943.4]
  assign RetimeWrapper_95_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61945.4]
  assign RetimeWrapper_95_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@61944.4]
  assign RetimeWrapper_96_clock = clock; // @[:@61969.4]
  assign RetimeWrapper_96_reset = reset; // @[:@61970.4]
  assign RetimeWrapper_96_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61972.4]
  assign RetimeWrapper_96_io_in = x739_sum_1_io_result; // @[package.scala 94:16:@61971.4]
  assign x512_sum_1_clock = clock; // @[:@61980.4]
  assign x512_sum_1_reset = reset; // @[:@61981.4]
  assign x512_sum_1_io_a = RetimeWrapper_96_io_out; // @[Math.scala 151:17:@61982.4]
  assign x512_sum_1_io_b = RetimeWrapper_76_io_out; // @[Math.scala 152:17:@61983.4]
  assign x512_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@61984.4]
  assign RetimeWrapper_97_clock = clock; // @[:@61990.4]
  assign RetimeWrapper_97_reset = reset; // @[:@61991.4]
  assign RetimeWrapper_97_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@61993.4]
  assign RetimeWrapper_97_io_in = ~ x510; // @[package.scala 94:16:@61992.4]
  assign RetimeWrapper_98_clock = clock; // @[:@61999.4]
  assign RetimeWrapper_98_reset = reset; // @[:@62000.4]
  assign RetimeWrapper_98_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62002.4]
  assign RetimeWrapper_98_io_in = x512_sum_1_io_result; // @[package.scala 94:16:@62001.4]
  assign RetimeWrapper_99_clock = clock; // @[:@62011.4]
  assign RetimeWrapper_99_reset = reset; // @[:@62012.4]
  assign RetimeWrapper_99_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62014.4]
  assign RetimeWrapper_99_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@62013.4]
  assign x517_sum_1_clock = clock; // @[:@62038.4]
  assign x517_sum_1_reset = reset; // @[:@62039.4]
  assign x517_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@62040.4]
  assign x517_sum_1_io_b = x440_div_1_io_result; // @[Math.scala 152:17:@62041.4]
  assign x517_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62042.4]
  assign RetimeWrapper_100_clock = clock; // @[:@62048.4]
  assign RetimeWrapper_100_reset = reset; // @[:@62049.4]
  assign RetimeWrapper_100_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62051.4]
  assign RetimeWrapper_100_io_in = ~ x515; // @[package.scala 94:16:@62050.4]
  assign RetimeWrapper_101_clock = clock; // @[:@62060.4]
  assign RetimeWrapper_101_reset = reset; // @[:@62061.4]
  assign RetimeWrapper_101_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62063.4]
  assign RetimeWrapper_101_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@62062.4]
  assign x522_sum_1_clock = clock; // @[:@62087.4]
  assign x522_sum_1_reset = reset; // @[:@62088.4]
  assign x522_sum_1_io_a = RetimeWrapper_88_io_out; // @[Math.scala 151:17:@62089.4]
  assign x522_sum_1_io_b = x449_div_1_io_result; // @[Math.scala 152:17:@62090.4]
  assign x522_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62091.4]
  assign RetimeWrapper_102_clock = clock; // @[:@62097.4]
  assign RetimeWrapper_102_reset = reset; // @[:@62098.4]
  assign RetimeWrapper_102_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62100.4]
  assign RetimeWrapper_102_io_in = ~ x520; // @[package.scala 94:16:@62099.4]
  assign RetimeWrapper_103_clock = clock; // @[:@62109.4]
  assign RetimeWrapper_103_reset = reset; // @[:@62110.4]
  assign RetimeWrapper_103_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62112.4]
  assign RetimeWrapper_103_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@62111.4]
  assign x525_1_clock = clock; // @[:@62132.4]
  assign x525_1_io_a = x383_lb_0_io_rPort_15_output_0; // @[Math.scala 263:17:@62134.4]
  assign x525_1_io_b = 32'h1; // @[Math.scala 264:17:@62135.4]
  assign x525_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62136.4]
  assign x526_1_clock = clock; // @[:@62144.4]
  assign x526_1_io_a = x383_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@62146.4]
  assign x526_1_io_b = 32'h2; // @[Math.scala 264:17:@62147.4]
  assign x526_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62148.4]
  assign x527_1_clock = clock; // @[:@62156.4]
  assign x527_1_io_a = x383_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@62158.4]
  assign x527_1_io_b = 32'h1; // @[Math.scala 264:17:@62159.4]
  assign x527_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62160.4]
  assign x528_1_clock = clock; // @[:@62168.4]
  assign x528_1_io_a = x383_lb_0_io_rPort_12_output_0; // @[Math.scala 263:17:@62170.4]
  assign x528_1_io_b = 32'h2; // @[Math.scala 264:17:@62171.4]
  assign x528_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62172.4]
  assign x529_1_clock = clock; // @[:@62180.4]
  assign x529_1_io_a = x383_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@62182.4]
  assign x529_1_io_b = 32'h4; // @[Math.scala 264:17:@62183.4]
  assign x529_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62184.4]
  assign x530_1_clock = clock; // @[:@62192.4]
  assign x530_1_io_a = x383_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@62194.4]
  assign x530_1_io_b = 32'h2; // @[Math.scala 264:17:@62195.4]
  assign x530_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62196.4]
  assign x531_1_clock = clock; // @[:@62204.4]
  assign x531_1_io_a = x383_lb_0_io_rPort_9_output_0; // @[Math.scala 263:17:@62206.4]
  assign x531_1_io_b = 32'h1; // @[Math.scala 264:17:@62207.4]
  assign x531_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62208.4]
  assign x532_1_clock = clock; // @[:@62216.4]
  assign x532_1_io_a = x383_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@62218.4]
  assign x532_1_io_b = 32'h2; // @[Math.scala 264:17:@62219.4]
  assign x532_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62220.4]
  assign x533_1_clock = clock; // @[:@62228.4]
  assign x533_1_io_a = x383_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@62230.4]
  assign x533_1_io_b = 32'h1; // @[Math.scala 264:17:@62231.4]
  assign x533_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62232.4]
  assign x534_x7_1_clock = clock; // @[:@62238.4]
  assign x534_x7_1_reset = reset; // @[:@62239.4]
  assign x534_x7_1_io_a = x525_1_io_result; // @[Math.scala 151:17:@62240.4]
  assign x534_x7_1_io_b = x526_1_io_result; // @[Math.scala 152:17:@62241.4]
  assign x534_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62242.4]
  assign x535_x8_1_clock = clock; // @[:@62248.4]
  assign x535_x8_1_reset = reset; // @[:@62249.4]
  assign x535_x8_1_io_a = x527_1_io_result; // @[Math.scala 151:17:@62250.4]
  assign x535_x8_1_io_b = x528_1_io_result; // @[Math.scala 152:17:@62251.4]
  assign x535_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62252.4]
  assign x536_x7_1_clock = clock; // @[:@62258.4]
  assign x536_x7_1_reset = reset; // @[:@62259.4]
  assign x536_x7_1_io_a = x529_1_io_result; // @[Math.scala 151:17:@62260.4]
  assign x536_x7_1_io_b = x530_1_io_result; // @[Math.scala 152:17:@62261.4]
  assign x536_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62262.4]
  assign x537_x8_1_clock = clock; // @[:@62268.4]
  assign x537_x8_1_reset = reset; // @[:@62269.4]
  assign x537_x8_1_io_a = x531_1_io_result; // @[Math.scala 151:17:@62270.4]
  assign x537_x8_1_io_b = x532_1_io_result; // @[Math.scala 152:17:@62271.4]
  assign x537_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62272.4]
  assign x538_x7_1_clock = clock; // @[:@62278.4]
  assign x538_x7_1_reset = reset; // @[:@62279.4]
  assign x538_x7_1_io_a = x534_x7_1_io_result; // @[Math.scala 151:17:@62280.4]
  assign x538_x7_1_io_b = x535_x8_1_io_result; // @[Math.scala 152:17:@62281.4]
  assign x538_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62282.4]
  assign x539_x8_1_clock = clock; // @[:@62288.4]
  assign x539_x8_1_reset = reset; // @[:@62289.4]
  assign x539_x8_1_io_a = x536_x7_1_io_result; // @[Math.scala 151:17:@62290.4]
  assign x539_x8_1_io_b = x537_x8_1_io_result; // @[Math.scala 152:17:@62291.4]
  assign x539_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62292.4]
  assign x540_x7_1_clock = clock; // @[:@62298.4]
  assign x540_x7_1_reset = reset; // @[:@62299.4]
  assign x540_x7_1_io_a = x538_x7_1_io_result; // @[Math.scala 151:17:@62300.4]
  assign x540_x7_1_io_b = x539_x8_1_io_result; // @[Math.scala 152:17:@62301.4]
  assign x540_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62302.4]
  assign RetimeWrapper_104_clock = clock; // @[:@62308.4]
  assign RetimeWrapper_104_reset = reset; // @[:@62309.4]
  assign RetimeWrapper_104_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62311.4]
  assign RetimeWrapper_104_io_in = x533_1_io_result; // @[package.scala 94:16:@62310.4]
  assign x541_sum_1_clock = clock; // @[:@62317.4]
  assign x541_sum_1_reset = reset; // @[:@62318.4]
  assign x541_sum_1_io_a = x540_x7_1_io_result; // @[Math.scala 151:17:@62319.4]
  assign x541_sum_1_io_b = RetimeWrapper_104_io_out; // @[Math.scala 152:17:@62320.4]
  assign x541_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62321.4]
  assign x542_1_io_b = x541_sum_1_io_result; // @[Math.scala 721:17:@62329.4]
  assign x543_mul_1_clock = clock; // @[:@62338.4]
  assign x543_mul_1_io_a = x542_1_io_result; // @[Math.scala 263:17:@62340.4]
  assign x543_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@62341.4]
  assign x543_mul_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62342.4]
  assign x544_1_io_b = x543_mul_1_io_result; // @[Math.scala 721:17:@62350.4]
  assign x545_1_clock = clock; // @[:@62359.4]
  assign x545_1_io_a = x383_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@62361.4]
  assign x545_1_io_b = 32'h1; // @[Math.scala 264:17:@62362.4]
  assign x545_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62363.4]
  assign x546_1_clock = clock; // @[:@62371.4]
  assign x546_1_io_a = x383_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@62373.4]
  assign x546_1_io_b = 32'h2; // @[Math.scala 264:17:@62374.4]
  assign x546_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62375.4]
  assign x547_1_clock = clock; // @[:@62383.4]
  assign x547_1_io_a = x383_lb_0_io_rPort_16_output_0; // @[Math.scala 263:17:@62385.4]
  assign x547_1_io_b = 32'h1; // @[Math.scala 264:17:@62386.4]
  assign x547_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62387.4]
  assign x548_1_clock = clock; // @[:@62395.4]
  assign x548_1_io_a = x383_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@62397.4]
  assign x548_1_io_b = 32'h2; // @[Math.scala 264:17:@62398.4]
  assign x548_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62399.4]
  assign x549_1_clock = clock; // @[:@62407.4]
  assign x549_1_io_a = x383_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@62409.4]
  assign x549_1_io_b = 32'h4; // @[Math.scala 264:17:@62410.4]
  assign x549_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62411.4]
  assign x550_1_clock = clock; // @[:@62421.4]
  assign x550_1_io_a = x383_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@62423.4]
  assign x550_1_io_b = 32'h2; // @[Math.scala 264:17:@62424.4]
  assign x550_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62425.4]
  assign x551_1_clock = clock; // @[:@62433.4]
  assign x551_1_io_a = x383_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@62435.4]
  assign x551_1_io_b = 32'h1; // @[Math.scala 264:17:@62436.4]
  assign x551_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62437.4]
  assign x552_1_clock = clock; // @[:@62445.4]
  assign x552_1_io_a = x383_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@62447.4]
  assign x552_1_io_b = 32'h2; // @[Math.scala 264:17:@62448.4]
  assign x552_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62449.4]
  assign x553_1_clock = clock; // @[:@62457.4]
  assign x553_1_io_a = x383_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@62459.4]
  assign x553_1_io_b = 32'h1; // @[Math.scala 264:17:@62460.4]
  assign x553_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62461.4]
  assign x554_x7_1_clock = clock; // @[:@62467.4]
  assign x554_x7_1_reset = reset; // @[:@62468.4]
  assign x554_x7_1_io_a = x545_1_io_result; // @[Math.scala 151:17:@62469.4]
  assign x554_x7_1_io_b = x546_1_io_result; // @[Math.scala 152:17:@62470.4]
  assign x554_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62471.4]
  assign x555_x8_1_clock = clock; // @[:@62477.4]
  assign x555_x8_1_reset = reset; // @[:@62478.4]
  assign x555_x8_1_io_a = x547_1_io_result; // @[Math.scala 151:17:@62479.4]
  assign x555_x8_1_io_b = x548_1_io_result; // @[Math.scala 152:17:@62480.4]
  assign x555_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62481.4]
  assign x556_x7_1_clock = clock; // @[:@62487.4]
  assign x556_x7_1_reset = reset; // @[:@62488.4]
  assign x556_x7_1_io_a = x549_1_io_result; // @[Math.scala 151:17:@62489.4]
  assign x556_x7_1_io_b = x550_1_io_result; // @[Math.scala 152:17:@62490.4]
  assign x556_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62491.4]
  assign x557_x8_1_clock = clock; // @[:@62497.4]
  assign x557_x8_1_reset = reset; // @[:@62498.4]
  assign x557_x8_1_io_a = x551_1_io_result; // @[Math.scala 151:17:@62499.4]
  assign x557_x8_1_io_b = x552_1_io_result; // @[Math.scala 152:17:@62500.4]
  assign x557_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62501.4]
  assign x558_x7_1_clock = clock; // @[:@62507.4]
  assign x558_x7_1_reset = reset; // @[:@62508.4]
  assign x558_x7_1_io_a = x554_x7_1_io_result; // @[Math.scala 151:17:@62509.4]
  assign x558_x7_1_io_b = x555_x8_1_io_result; // @[Math.scala 152:17:@62510.4]
  assign x558_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62511.4]
  assign x559_x8_1_clock = clock; // @[:@62517.4]
  assign x559_x8_1_reset = reset; // @[:@62518.4]
  assign x559_x8_1_io_a = x556_x7_1_io_result; // @[Math.scala 151:17:@62519.4]
  assign x559_x8_1_io_b = x557_x8_1_io_result; // @[Math.scala 152:17:@62520.4]
  assign x559_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62521.4]
  assign x560_x7_1_clock = clock; // @[:@62527.4]
  assign x560_x7_1_reset = reset; // @[:@62528.4]
  assign x560_x7_1_io_a = x558_x7_1_io_result; // @[Math.scala 151:17:@62529.4]
  assign x560_x7_1_io_b = x559_x8_1_io_result; // @[Math.scala 152:17:@62530.4]
  assign x560_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62531.4]
  assign RetimeWrapper_105_clock = clock; // @[:@62537.4]
  assign RetimeWrapper_105_reset = reset; // @[:@62538.4]
  assign RetimeWrapper_105_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62540.4]
  assign RetimeWrapper_105_io_in = x553_1_io_result; // @[package.scala 94:16:@62539.4]
  assign x561_sum_1_clock = clock; // @[:@62546.4]
  assign x561_sum_1_reset = reset; // @[:@62547.4]
  assign x561_sum_1_io_a = x560_x7_1_io_result; // @[Math.scala 151:17:@62548.4]
  assign x561_sum_1_io_b = RetimeWrapper_105_io_out; // @[Math.scala 152:17:@62549.4]
  assign x561_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62550.4]
  assign x562_1_io_b = x561_sum_1_io_result; // @[Math.scala 721:17:@62558.4]
  assign x563_mul_1_clock = clock; // @[:@62567.4]
  assign x563_mul_1_io_a = x562_1_io_result; // @[Math.scala 263:17:@62569.4]
  assign x563_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@62570.4]
  assign x563_mul_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62571.4]
  assign x564_1_io_b = x563_mul_1_io_result; // @[Math.scala 721:17:@62579.4]
  assign x565_1_clock = clock; // @[:@62588.4]
  assign x565_1_io_a = x383_lb_0_io_rPort_16_output_0; // @[Math.scala 263:17:@62590.4]
  assign x565_1_io_b = 32'h2; // @[Math.scala 264:17:@62591.4]
  assign x565_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62592.4]
  assign x566_1_clock = clock; // @[:@62600.4]
  assign x566_1_io_a = x383_lb_0_io_rPort_17_output_0; // @[Math.scala 263:17:@62602.4]
  assign x566_1_io_b = 32'h1; // @[Math.scala 264:17:@62603.4]
  assign x566_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62604.4]
  assign x567_1_clock = clock; // @[:@62612.4]
  assign x567_1_io_a = x383_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@62614.4]
  assign x567_1_io_b = 32'h4; // @[Math.scala 264:17:@62615.4]
  assign x567_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62616.4]
  assign x568_1_clock = clock; // @[:@62624.4]
  assign x568_1_io_a = x383_lb_0_io_rPort_14_output_0; // @[Math.scala 263:17:@62626.4]
  assign x568_1_io_b = 32'h2; // @[Math.scala 264:17:@62627.4]
  assign x568_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62628.4]
  assign x569_1_clock = clock; // @[:@62636.4]
  assign x569_1_io_a = x383_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@62638.4]
  assign x569_1_io_b = 32'h2; // @[Math.scala 264:17:@62639.4]
  assign x569_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62640.4]
  assign x570_1_clock = clock; // @[:@62648.4]
  assign x570_1_io_a = x383_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@62650.4]
  assign x570_1_io_b = 32'h1; // @[Math.scala 264:17:@62651.4]
  assign x570_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62652.4]
  assign x571_x7_1_clock = clock; // @[:@62658.4]
  assign x571_x7_1_reset = reset; // @[:@62659.4]
  assign x571_x7_1_io_a = x527_1_io_result; // @[Math.scala 151:17:@62660.4]
  assign x571_x7_1_io_b = x565_1_io_result; // @[Math.scala 152:17:@62661.4]
  assign x571_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62662.4]
  assign x572_x8_1_clock = clock; // @[:@62668.4]
  assign x572_x8_1_reset = reset; // @[:@62669.4]
  assign x572_x8_1_io_a = x566_1_io_result; // @[Math.scala 151:17:@62670.4]
  assign x572_x8_1_io_b = x530_1_io_result; // @[Math.scala 152:17:@62671.4]
  assign x572_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62672.4]
  assign x573_x7_1_clock = clock; // @[:@62678.4]
  assign x573_x7_1_reset = reset; // @[:@62679.4]
  assign x573_x7_1_io_a = x567_1_io_result; // @[Math.scala 151:17:@62680.4]
  assign x573_x7_1_io_b = x568_1_io_result; // @[Math.scala 152:17:@62681.4]
  assign x573_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62682.4]
  assign x574_x8_1_clock = clock; // @[:@62688.4]
  assign x574_x8_1_reset = reset; // @[:@62689.4]
  assign x574_x8_1_io_a = x533_1_io_result; // @[Math.scala 151:17:@62690.4]
  assign x574_x8_1_io_b = x569_1_io_result; // @[Math.scala 152:17:@62691.4]
  assign x574_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62692.4]
  assign x575_x7_1_clock = clock; // @[:@62698.4]
  assign x575_x7_1_reset = reset; // @[:@62699.4]
  assign x575_x7_1_io_a = x571_x7_1_io_result; // @[Math.scala 151:17:@62700.4]
  assign x575_x7_1_io_b = x572_x8_1_io_result; // @[Math.scala 152:17:@62701.4]
  assign x575_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62702.4]
  assign x576_x8_1_clock = clock; // @[:@62708.4]
  assign x576_x8_1_reset = reset; // @[:@62709.4]
  assign x576_x8_1_io_a = x573_x7_1_io_result; // @[Math.scala 151:17:@62710.4]
  assign x576_x8_1_io_b = x574_x8_1_io_result; // @[Math.scala 152:17:@62711.4]
  assign x576_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62712.4]
  assign x577_x7_1_clock = clock; // @[:@62718.4]
  assign x577_x7_1_reset = reset; // @[:@62719.4]
  assign x577_x7_1_io_a = x575_x7_1_io_result; // @[Math.scala 151:17:@62720.4]
  assign x577_x7_1_io_b = x576_x8_1_io_result; // @[Math.scala 152:17:@62721.4]
  assign x577_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62722.4]
  assign RetimeWrapper_106_clock = clock; // @[:@62728.4]
  assign RetimeWrapper_106_reset = reset; // @[:@62729.4]
  assign RetimeWrapper_106_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62731.4]
  assign RetimeWrapper_106_io_in = x570_1_io_result; // @[package.scala 94:16:@62730.4]
  assign x578_sum_1_clock = clock; // @[:@62737.4]
  assign x578_sum_1_reset = reset; // @[:@62738.4]
  assign x578_sum_1_io_a = x577_x7_1_io_result; // @[Math.scala 151:17:@62739.4]
  assign x578_sum_1_io_b = RetimeWrapper_106_io_out; // @[Math.scala 152:17:@62740.4]
  assign x578_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62741.4]
  assign x579_1_io_b = x578_sum_1_io_result; // @[Math.scala 721:17:@62749.4]
  assign x580_mul_1_clock = clock; // @[:@62758.4]
  assign x580_mul_1_io_a = x579_1_io_result; // @[Math.scala 263:17:@62760.4]
  assign x580_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@62761.4]
  assign x580_mul_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62762.4]
  assign x581_1_io_b = x580_mul_1_io_result; // @[Math.scala 721:17:@62770.4]
  assign x582_1_clock = clock; // @[:@62779.4]
  assign x582_1_io_a = x383_lb_0_io_rPort_17_output_0; // @[Math.scala 263:17:@62781.4]
  assign x582_1_io_b = 32'h2; // @[Math.scala 264:17:@62782.4]
  assign x582_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62783.4]
  assign x583_1_clock = clock; // @[:@62791.4]
  assign x583_1_io_a = x383_lb_0_io_rPort_10_output_0; // @[Math.scala 263:17:@62793.4]
  assign x583_1_io_b = 32'h1; // @[Math.scala 264:17:@62794.4]
  assign x583_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62795.4]
  assign x584_1_clock = clock; // @[:@62803.4]
  assign x584_1_io_a = x383_lb_0_io_rPort_14_output_0; // @[Math.scala 263:17:@62805.4]
  assign x584_1_io_b = 32'h4; // @[Math.scala 264:17:@62806.4]
  assign x584_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62807.4]
  assign x585_1_clock = clock; // @[:@62815.4]
  assign x585_1_io_a = x383_lb_0_io_rPort_13_output_0; // @[Math.scala 263:17:@62817.4]
  assign x585_1_io_b = 32'h2; // @[Math.scala 264:17:@62818.4]
  assign x585_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62819.4]
  assign x586_1_clock = clock; // @[:@62827.4]
  assign x586_1_io_a = x383_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@62829.4]
  assign x586_1_io_b = 32'h2; // @[Math.scala 264:17:@62830.4]
  assign x586_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62831.4]
  assign x587_1_clock = clock; // @[:@62839.4]
  assign x587_1_io_a = x383_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@62841.4]
  assign x587_1_io_b = 32'h1; // @[Math.scala 264:17:@62842.4]
  assign x587_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62843.4]
  assign x588_x7_1_clock = clock; // @[:@62849.4]
  assign x588_x7_1_reset = reset; // @[:@62850.4]
  assign x588_x7_1_io_a = x547_1_io_result; // @[Math.scala 151:17:@62851.4]
  assign x588_x7_1_io_b = x582_1_io_result; // @[Math.scala 152:17:@62852.4]
  assign x588_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62853.4]
  assign x589_x8_1_clock = clock; // @[:@62859.4]
  assign x589_x8_1_reset = reset; // @[:@62860.4]
  assign x589_x8_1_io_a = x583_1_io_result; // @[Math.scala 151:17:@62861.4]
  assign x589_x8_1_io_b = x550_1_io_result; // @[Math.scala 152:17:@62862.4]
  assign x589_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62863.4]
  assign x590_x7_1_clock = clock; // @[:@62869.4]
  assign x590_x7_1_reset = reset; // @[:@62870.4]
  assign x590_x7_1_io_a = x584_1_io_result; // @[Math.scala 151:17:@62871.4]
  assign x590_x7_1_io_b = x585_1_io_result; // @[Math.scala 152:17:@62872.4]
  assign x590_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62873.4]
  assign x591_x8_1_clock = clock; // @[:@62879.4]
  assign x591_x8_1_reset = reset; // @[:@62880.4]
  assign x591_x8_1_io_a = x553_1_io_result; // @[Math.scala 151:17:@62881.4]
  assign x591_x8_1_io_b = x586_1_io_result; // @[Math.scala 152:17:@62882.4]
  assign x591_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62883.4]
  assign x592_x7_1_clock = clock; // @[:@62889.4]
  assign x592_x7_1_reset = reset; // @[:@62890.4]
  assign x592_x7_1_io_a = x588_x7_1_io_result; // @[Math.scala 151:17:@62891.4]
  assign x592_x7_1_io_b = x589_x8_1_io_result; // @[Math.scala 152:17:@62892.4]
  assign x592_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62893.4]
  assign x593_x8_1_clock = clock; // @[:@62899.4]
  assign x593_x8_1_reset = reset; // @[:@62900.4]
  assign x593_x8_1_io_a = x590_x7_1_io_result; // @[Math.scala 151:17:@62901.4]
  assign x593_x8_1_io_b = x591_x8_1_io_result; // @[Math.scala 152:17:@62902.4]
  assign x593_x8_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62903.4]
  assign x594_x7_1_clock = clock; // @[:@62909.4]
  assign x594_x7_1_reset = reset; // @[:@62910.4]
  assign x594_x7_1_io_a = x592_x7_1_io_result; // @[Math.scala 151:17:@62911.4]
  assign x594_x7_1_io_b = x593_x8_1_io_result; // @[Math.scala 152:17:@62912.4]
  assign x594_x7_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62913.4]
  assign RetimeWrapper_107_clock = clock; // @[:@62919.4]
  assign RetimeWrapper_107_reset = reset; // @[:@62920.4]
  assign RetimeWrapper_107_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62922.4]
  assign RetimeWrapper_107_io_in = x587_1_io_result; // @[package.scala 94:16:@62921.4]
  assign x595_sum_1_clock = clock; // @[:@62928.4]
  assign x595_sum_1_reset = reset; // @[:@62929.4]
  assign x595_sum_1_io_a = x594_x7_1_io_result; // @[Math.scala 151:17:@62930.4]
  assign x595_sum_1_io_b = RetimeWrapper_107_io_out; // @[Math.scala 152:17:@62931.4]
  assign x595_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@62932.4]
  assign x596_1_io_b = x595_sum_1_io_result; // @[Math.scala 721:17:@62942.4]
  assign x597_mul_1_clock = clock; // @[:@62951.4]
  assign x597_mul_1_io_a = x596_1_io_result; // @[Math.scala 263:17:@62953.4]
  assign x597_mul_1_io_b = 32'h8; // @[Math.scala 264:17:@62954.4]
  assign x597_mul_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@62955.4]
  assign x598_1_io_b = x597_mul_1_io_result; // @[Math.scala 721:17:@62963.4]
  assign RetimeWrapper_108_clock = clock; // @[:@62970.4]
  assign RetimeWrapper_108_reset = reset; // @[:@62971.4]
  assign RetimeWrapper_108_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62973.4]
  assign RetimeWrapper_108_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@62972.4]
  assign RetimeWrapper_109_clock = clock; // @[:@62979.4]
  assign RetimeWrapper_109_reset = reset; // @[:@62980.4]
  assign RetimeWrapper_109_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62982.4]
  assign RetimeWrapper_109_io_in = x389_1_io_result; // @[package.scala 94:16:@62981.4]
  assign RetimeWrapper_110_clock = clock; // @[:@62988.4]
  assign RetimeWrapper_110_reset = reset; // @[:@62989.4]
  assign RetimeWrapper_110_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@62991.4]
  assign RetimeWrapper_110_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@62990.4]
  assign RetimeWrapper_111_clock = clock; // @[:@62997.4]
  assign RetimeWrapper_111_reset = reset; // @[:@62998.4]
  assign RetimeWrapper_111_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63000.4]
  assign RetimeWrapper_111_io_in = x598_1_io_result; // @[package.scala 94:16:@62999.4]
  assign RetimeWrapper_112_clock = clock; // @[:@63006.4]
  assign RetimeWrapper_112_reset = reset; // @[:@63007.4]
  assign RetimeWrapper_112_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63009.4]
  assign RetimeWrapper_112_io_in = x393_sum_1_io_result; // @[package.scala 94:16:@63008.4]
  assign RetimeWrapper_113_clock = clock; // @[:@63015.4]
  assign RetimeWrapper_113_reset = reset; // @[:@63016.4]
  assign RetimeWrapper_113_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63018.4]
  assign RetimeWrapper_113_io_in = $unsigned(_T_264); // @[package.scala 94:16:@63017.4]
  assign RetimeWrapper_114_clock = clock; // @[:@63026.4]
  assign RetimeWrapper_114_reset = reset; // @[:@63027.4]
  assign RetimeWrapper_114_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63029.4]
  assign RetimeWrapper_114_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63028.4]
  assign RetimeWrapper_115_clock = clock; // @[:@63047.4]
  assign RetimeWrapper_115_reset = reset; // @[:@63048.4]
  assign RetimeWrapper_115_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63050.4]
  assign RetimeWrapper_115_io_in = x397_1_io_result; // @[package.scala 94:16:@63049.4]
  assign RetimeWrapper_116_clock = clock; // @[:@63056.4]
  assign RetimeWrapper_116_reset = reset; // @[:@63057.4]
  assign RetimeWrapper_116_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63059.4]
  assign RetimeWrapper_116_io_in = x399_sum_1_io_result; // @[package.scala 94:16:@63058.4]
  assign RetimeWrapper_117_clock = clock; // @[:@63065.4]
  assign RetimeWrapper_117_reset = reset; // @[:@63066.4]
  assign RetimeWrapper_117_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63068.4]
  assign RetimeWrapper_117_io_in = x581_1_io_result; // @[package.scala 94:16:@63067.4]
  assign RetimeWrapper_118_clock = clock; // @[:@63076.4]
  assign RetimeWrapper_118_reset = reset; // @[:@63077.4]
  assign RetimeWrapper_118_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63079.4]
  assign RetimeWrapper_118_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63078.4]
  assign RetimeWrapper_119_clock = clock; // @[:@63097.4]
  assign RetimeWrapper_119_reset = reset; // @[:@63098.4]
  assign RetimeWrapper_119_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63100.4]
  assign RetimeWrapper_119_io_in = x403_1_io_result; // @[package.scala 94:16:@63099.4]
  assign RetimeWrapper_120_clock = clock; // @[:@63106.4]
  assign RetimeWrapper_120_reset = reset; // @[:@63107.4]
  assign RetimeWrapper_120_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63109.4]
  assign RetimeWrapper_120_io_in = x405_sum_1_io_result; // @[package.scala 94:16:@63108.4]
  assign RetimeWrapper_121_clock = clock; // @[:@63115.4]
  assign RetimeWrapper_121_reset = reset; // @[:@63116.4]
  assign RetimeWrapper_121_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63118.4]
  assign RetimeWrapper_121_io_in = x564_1_io_result; // @[package.scala 94:16:@63117.4]
  assign RetimeWrapper_122_clock = clock; // @[:@63126.4]
  assign RetimeWrapper_122_reset = reset; // @[:@63127.4]
  assign RetimeWrapper_122_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63129.4]
  assign RetimeWrapper_122_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63128.4]
  assign RetimeWrapper_123_clock = clock; // @[:@63147.4]
  assign RetimeWrapper_123_reset = reset; // @[:@63148.4]
  assign RetimeWrapper_123_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63150.4]
  assign RetimeWrapper_123_io_in = x411_sum_1_io_result; // @[package.scala 94:16:@63149.4]
  assign RetimeWrapper_124_clock = clock; // @[:@63156.4]
  assign RetimeWrapper_124_reset = reset; // @[:@63157.4]
  assign RetimeWrapper_124_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63159.4]
  assign RetimeWrapper_124_io_in = x409_1_io_result; // @[package.scala 94:16:@63158.4]
  assign RetimeWrapper_125_clock = clock; // @[:@63165.4]
  assign RetimeWrapper_125_reset = reset; // @[:@63166.4]
  assign RetimeWrapper_125_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63168.4]
  assign RetimeWrapper_125_io_in = x544_1_io_result; // @[package.scala 94:16:@63167.4]
  assign RetimeWrapper_126_clock = clock; // @[:@63176.4]
  assign RetimeWrapper_126_reset = reset; // @[:@63177.4]
  assign RetimeWrapper_126_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63179.4]
  assign RetimeWrapper_126_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63178.4]
  assign RetimeWrapper_127_clock = clock; // @[:@63197.4]
  assign RetimeWrapper_127_reset = reset; // @[:@63198.4]
  assign RetimeWrapper_127_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63200.4]
  assign RetimeWrapper_127_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@63199.4]
  assign RetimeWrapper_128_clock = clock; // @[:@63206.4]
  assign RetimeWrapper_128_reset = reset; // @[:@63207.4]
  assign RetimeWrapper_128_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63209.4]
  assign RetimeWrapper_128_io_in = ~ x416; // @[package.scala 94:16:@63208.4]
  assign RetimeWrapper_129_clock = clock; // @[:@63215.4]
  assign RetimeWrapper_129_reset = reset; // @[:@63216.4]
  assign RetimeWrapper_129_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63218.4]
  assign RetimeWrapper_129_io_in = x411_sum_1_io_result; // @[package.scala 94:16:@63217.4]
  assign RetimeWrapper_130_clock = clock; // @[:@63224.4]
  assign RetimeWrapper_130_reset = reset; // @[:@63225.4]
  assign RetimeWrapper_130_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63227.4]
  assign RetimeWrapper_130_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@63226.4]
  assign RetimeWrapper_131_clock = clock; // @[:@63233.4]
  assign RetimeWrapper_131_reset = reset; // @[:@63234.4]
  assign RetimeWrapper_131_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63236.4]
  assign RetimeWrapper_131_io_in = $unsigned(_T_264); // @[package.scala 94:16:@63235.4]
  assign RetimeWrapper_132_clock = clock; // @[:@63242.4]
  assign RetimeWrapper_132_reset = reset; // @[:@63243.4]
  assign RetimeWrapper_132_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63245.4]
  assign RetimeWrapper_132_io_in = x409_1_io_result; // @[package.scala 94:16:@63244.4]
  assign RetimeWrapper_133_clock = clock; // @[:@63254.4]
  assign RetimeWrapper_133_reset = reset; // @[:@63255.4]
  assign RetimeWrapper_133_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63257.4]
  assign RetimeWrapper_133_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63256.4]
  assign RetimeWrapper_134_clock = clock; // @[:@63275.4]
  assign RetimeWrapper_134_reset = reset; // @[:@63276.4]
  assign RetimeWrapper_134_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63278.4]
  assign RetimeWrapper_134_io_in = x403_1_io_result; // @[package.scala 94:16:@63277.4]
  assign RetimeWrapper_135_clock = clock; // @[:@63284.4]
  assign RetimeWrapper_135_reset = reset; // @[:@63285.4]
  assign RetimeWrapper_135_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63287.4]
  assign RetimeWrapper_135_io_in = x405_sum_1_io_result; // @[package.scala 94:16:@63286.4]
  assign RetimeWrapper_136_clock = clock; // @[:@63293.4]
  assign RetimeWrapper_136_reset = reset; // @[:@63294.4]
  assign RetimeWrapper_136_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63296.4]
  assign RetimeWrapper_136_io_in = ~ x421; // @[package.scala 94:16:@63295.4]
  assign RetimeWrapper_137_clock = clock; // @[:@63305.4]
  assign RetimeWrapper_137_reset = reset; // @[:@63306.4]
  assign RetimeWrapper_137_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63308.4]
  assign RetimeWrapper_137_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63307.4]
  assign RetimeWrapper_138_clock = clock; // @[:@63326.4]
  assign RetimeWrapper_138_reset = reset; // @[:@63327.4]
  assign RetimeWrapper_138_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63329.4]
  assign RetimeWrapper_138_io_in = x397_1_io_result; // @[package.scala 94:16:@63328.4]
  assign RetimeWrapper_139_clock = clock; // @[:@63335.4]
  assign RetimeWrapper_139_reset = reset; // @[:@63336.4]
  assign RetimeWrapper_139_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63338.4]
  assign RetimeWrapper_139_io_in = x399_sum_1_io_result; // @[package.scala 94:16:@63337.4]
  assign RetimeWrapper_140_clock = clock; // @[:@63344.4]
  assign RetimeWrapper_140_reset = reset; // @[:@63345.4]
  assign RetimeWrapper_140_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63347.4]
  assign RetimeWrapper_140_io_in = ~ x426; // @[package.scala 94:16:@63346.4]
  assign RetimeWrapper_141_clock = clock; // @[:@63356.4]
  assign RetimeWrapper_141_reset = reset; // @[:@63357.4]
  assign RetimeWrapper_141_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63359.4]
  assign RetimeWrapper_141_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63358.4]
  assign RetimeWrapper_142_clock = clock; // @[:@63377.4]
  assign RetimeWrapper_142_reset = reset; // @[:@63378.4]
  assign RetimeWrapper_142_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63380.4]
  assign RetimeWrapper_142_io_in = x389_1_io_result; // @[package.scala 94:16:@63379.4]
  assign RetimeWrapper_143_clock = clock; // @[:@63386.4]
  assign RetimeWrapper_143_reset = reset; // @[:@63387.4]
  assign RetimeWrapper_143_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63389.4]
  assign RetimeWrapper_143_io_in = x393_sum_1_io_result; // @[package.scala 94:16:@63388.4]
  assign RetimeWrapper_144_clock = clock; // @[:@63395.4]
  assign RetimeWrapper_144_reset = reset; // @[:@63396.4]
  assign RetimeWrapper_144_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63398.4]
  assign RetimeWrapper_144_io_in = ~ x431; // @[package.scala 94:16:@63397.4]
  assign RetimeWrapper_145_clock = clock; // @[:@63407.4]
  assign RetimeWrapper_145_reset = reset; // @[:@63408.4]
  assign RetimeWrapper_145_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63410.4]
  assign RetimeWrapper_145_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63409.4]
  assign RetimeWrapper_146_clock = clock; // @[:@63428.4]
  assign RetimeWrapper_146_reset = reset; // @[:@63429.4]
  assign RetimeWrapper_146_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63431.4]
  assign RetimeWrapper_146_io_in = x439_1_io_result; // @[package.scala 94:16:@63430.4]
  assign RetimeWrapper_147_clock = clock; // @[:@63437.4]
  assign RetimeWrapper_147_reset = reset; // @[:@63438.4]
  assign RetimeWrapper_147_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63440.4]
  assign RetimeWrapper_147_io_in = ~ x437; // @[package.scala 94:16:@63439.4]
  assign RetimeWrapper_148_clock = clock; // @[:@63446.4]
  assign RetimeWrapper_148_reset = reset; // @[:@63447.4]
  assign RetimeWrapper_148_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63449.4]
  assign RetimeWrapper_148_io_in = x441_sum_1_io_result; // @[package.scala 94:16:@63448.4]
  assign RetimeWrapper_149_clock = clock; // @[:@63458.4]
  assign RetimeWrapper_149_reset = reset; // @[:@63459.4]
  assign RetimeWrapper_149_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63461.4]
  assign RetimeWrapper_149_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63460.4]
  assign RetimeWrapper_150_clock = clock; // @[:@63479.4]
  assign RetimeWrapper_150_reset = reset; // @[:@63480.4]
  assign RetimeWrapper_150_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63482.4]
  assign RetimeWrapper_150_io_in = x461_sum_1_io_result; // @[package.scala 94:16:@63481.4]
  assign RetimeWrapper_151_clock = clock; // @[:@63488.4]
  assign RetimeWrapper_151_reset = reset; // @[:@63489.4]
  assign RetimeWrapper_151_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63491.4]
  assign RetimeWrapper_151_io_in = ~ x456; // @[package.scala 94:16:@63490.4]
  assign RetimeWrapper_152_clock = clock; // @[:@63497.4]
  assign RetimeWrapper_152_reset = reset; // @[:@63498.4]
  assign RetimeWrapper_152_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63500.4]
  assign RetimeWrapper_152_io_in = $unsigned(_T_885); // @[package.scala 94:16:@63499.4]
  assign RetimeWrapper_153_clock = clock; // @[:@63509.4]
  assign RetimeWrapper_153_reset = reset; // @[:@63510.4]
  assign RetimeWrapper_153_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63512.4]
  assign RetimeWrapper_153_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63511.4]
  assign RetimeWrapper_154_clock = clock; // @[:@63530.4]
  assign RetimeWrapper_154_reset = reset; // @[:@63531.4]
  assign RetimeWrapper_154_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63533.4]
  assign RetimeWrapper_154_io_in = x466_sum_1_io_result; // @[package.scala 94:16:@63532.4]
  assign RetimeWrapper_155_clock = clock; // @[:@63539.4]
  assign RetimeWrapper_155_reset = reset; // @[:@63540.4]
  assign RetimeWrapper_155_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63542.4]
  assign RetimeWrapper_155_io_in = ~ x464; // @[package.scala 94:16:@63541.4]
  assign RetimeWrapper_156_clock = clock; // @[:@63551.4]
  assign RetimeWrapper_156_reset = reset; // @[:@63552.4]
  assign RetimeWrapper_156_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63554.4]
  assign RetimeWrapper_156_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63553.4]
  assign RetimeWrapper_157_clock = clock; // @[:@63572.4]
  assign RetimeWrapper_157_reset = reset; // @[:@63573.4]
  assign RetimeWrapper_157_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63575.4]
  assign RetimeWrapper_157_io_in = x471_sum_1_io_result; // @[package.scala 94:16:@63574.4]
  assign RetimeWrapper_158_clock = clock; // @[:@63581.4]
  assign RetimeWrapper_158_reset = reset; // @[:@63582.4]
  assign RetimeWrapper_158_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63584.4]
  assign RetimeWrapper_158_io_in = ~ x469; // @[package.scala 94:16:@63583.4]
  assign RetimeWrapper_159_clock = clock; // @[:@63593.4]
  assign RetimeWrapper_159_reset = reset; // @[:@63594.4]
  assign RetimeWrapper_159_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63596.4]
  assign RetimeWrapper_159_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63595.4]
  assign RetimeWrapper_160_clock = clock; // @[:@63614.4]
  assign RetimeWrapper_160_reset = reset; // @[:@63615.4]
  assign RetimeWrapper_160_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63617.4]
  assign RetimeWrapper_160_io_in = ~ x474; // @[package.scala 94:16:@63616.4]
  assign RetimeWrapper_161_clock = clock; // @[:@63623.4]
  assign RetimeWrapper_161_reset = reset; // @[:@63624.4]
  assign RetimeWrapper_161_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63626.4]
  assign RetimeWrapper_161_io_in = x476_sum_1_io_result; // @[package.scala 94:16:@63625.4]
  assign RetimeWrapper_162_clock = clock; // @[:@63635.4]
  assign RetimeWrapper_162_reset = reset; // @[:@63636.4]
  assign RetimeWrapper_162_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63638.4]
  assign RetimeWrapper_162_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63637.4]
  assign RetimeWrapper_163_clock = clock; // @[:@63656.4]
  assign RetimeWrapper_163_reset = reset; // @[:@63657.4]
  assign RetimeWrapper_163_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63659.4]
  assign RetimeWrapper_163_io_in = x481_sum_1_io_result; // @[package.scala 94:16:@63658.4]
  assign RetimeWrapper_164_clock = clock; // @[:@63665.4]
  assign RetimeWrapper_164_reset = reset; // @[:@63666.4]
  assign RetimeWrapper_164_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63668.4]
  assign RetimeWrapper_164_io_in = ~ x479; // @[package.scala 94:16:@63667.4]
  assign RetimeWrapper_165_clock = clock; // @[:@63677.4]
  assign RetimeWrapper_165_reset = reset; // @[:@63678.4]
  assign RetimeWrapper_165_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@63680.4]
  assign RetimeWrapper_165_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@63679.4]
  assign x625_1_clock = clock; // @[:@63702.4]
  assign x625_1_io_a = x384_lb2_0_io_rPort_3_output_0; // @[Math.scala 263:17:@63704.4]
  assign x625_1_io_b = 32'h1; // @[Math.scala 264:17:@63705.4]
  assign x625_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63706.4]
  assign x626_1_clock = clock; // @[:@63714.4]
  assign x626_1_io_a = x384_lb2_0_io_rPort_9_output_0; // @[Math.scala 263:17:@63716.4]
  assign x626_1_io_b = 32'h2; // @[Math.scala 264:17:@63717.4]
  assign x626_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63718.4]
  assign x627_1_clock = clock; // @[:@63726.4]
  assign x627_1_io_a = x384_lb2_0_io_rPort_2_output_0; // @[Math.scala 263:17:@63728.4]
  assign x627_1_io_b = 32'h4; // @[Math.scala 264:17:@63729.4]
  assign x627_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63730.4]
  assign x628_1_clock = clock; // @[:@63738.4]
  assign x628_1_io_a = x384_lb2_0_io_rPort_7_output_0; // @[Math.scala 263:17:@63740.4]
  assign x628_1_io_b = 32'h1; // @[Math.scala 264:17:@63741.4]
  assign x628_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63742.4]
  assign x629_x9_1_clock = clock; // @[:@63748.4]
  assign x629_x9_1_reset = reset; // @[:@63749.4]
  assign x629_x9_1_io_a = x625_1_io_result; // @[Math.scala 151:17:@63750.4]
  assign x629_x9_1_io_b = x626_1_io_result; // @[Math.scala 152:17:@63751.4]
  assign x629_x9_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63752.4]
  assign x630_x10_1_clock = clock; // @[:@63758.4]
  assign x630_x10_1_reset = reset; // @[:@63759.4]
  assign x630_x10_1_io_a = x627_1_io_result; // @[Math.scala 151:17:@63760.4]
  assign x630_x10_1_io_b = x628_1_io_result; // @[Math.scala 152:17:@63761.4]
  assign x630_x10_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63762.4]
  assign x631_sum_1_clock = clock; // @[:@63768.4]
  assign x631_sum_1_reset = reset; // @[:@63769.4]
  assign x631_sum_1_io_a = x629_x9_1_io_result; // @[Math.scala 151:17:@63770.4]
  assign x631_sum_1_io_b = x630_x10_1_io_result; // @[Math.scala 152:17:@63771.4]
  assign x631_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63772.4]
  assign x632_1_io_b = x631_sum_1_io_result; // @[Math.scala 721:17:@63780.4]
  assign x633_mul_1_clock = clock; // @[:@63789.4]
  assign x633_mul_1_io_a = x632_1_io_result; // @[Math.scala 263:17:@63791.4]
  assign x633_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@63792.4]
  assign x633_mul_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63793.4]
  assign x634_1_io_b = x633_mul_1_io_result; // @[Math.scala 721:17:@63801.4]
  assign x635_1_clock = clock; // @[:@63810.4]
  assign x635_1_io_a = x384_lb2_0_io_rPort_9_output_0; // @[Math.scala 263:17:@63812.4]
  assign x635_1_io_b = 32'h1; // @[Math.scala 264:17:@63813.4]
  assign x635_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63814.4]
  assign x636_1_clock = clock; // @[:@63822.4]
  assign x636_1_io_a = x384_lb2_0_io_rPort_5_output_0; // @[Math.scala 263:17:@63824.4]
  assign x636_1_io_b = 32'h2; // @[Math.scala 264:17:@63825.4]
  assign x636_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63826.4]
  assign x637_1_clock = clock; // @[:@63834.4]
  assign x637_1_io_a = x384_lb2_0_io_rPort_7_output_0; // @[Math.scala 263:17:@63836.4]
  assign x637_1_io_b = 32'h4; // @[Math.scala 264:17:@63837.4]
  assign x637_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63838.4]
  assign x638_1_clock = clock; // @[:@63846.4]
  assign x638_1_io_a = x384_lb2_0_io_rPort_0_output_0; // @[Math.scala 263:17:@63848.4]
  assign x638_1_io_b = 32'h1; // @[Math.scala 264:17:@63849.4]
  assign x638_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63850.4]
  assign x639_x9_1_clock = clock; // @[:@63856.4]
  assign x639_x9_1_reset = reset; // @[:@63857.4]
  assign x639_x9_1_io_a = x635_1_io_result; // @[Math.scala 151:17:@63858.4]
  assign x639_x9_1_io_b = x636_1_io_result; // @[Math.scala 152:17:@63859.4]
  assign x639_x9_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63860.4]
  assign x640_x10_1_clock = clock; // @[:@63866.4]
  assign x640_x10_1_reset = reset; // @[:@63867.4]
  assign x640_x10_1_io_a = x637_1_io_result; // @[Math.scala 151:17:@63868.4]
  assign x640_x10_1_io_b = x638_1_io_result; // @[Math.scala 152:17:@63869.4]
  assign x640_x10_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63870.4]
  assign x641_sum_1_clock = clock; // @[:@63876.4]
  assign x641_sum_1_reset = reset; // @[:@63877.4]
  assign x641_sum_1_io_a = x639_x9_1_io_result; // @[Math.scala 151:17:@63878.4]
  assign x641_sum_1_io_b = x640_x10_1_io_result; // @[Math.scala 152:17:@63879.4]
  assign x641_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63880.4]
  assign x642_1_io_b = x641_sum_1_io_result; // @[Math.scala 721:17:@63888.4]
  assign x643_mul_1_clock = clock; // @[:@63897.4]
  assign x643_mul_1_io_a = x642_1_io_result; // @[Math.scala 263:17:@63899.4]
  assign x643_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@63900.4]
  assign x643_mul_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63901.4]
  assign x644_1_io_b = x643_mul_1_io_result; // @[Math.scala 721:17:@63909.4]
  assign x645_1_clock = clock; // @[:@63918.4]
  assign x645_1_io_a = x384_lb2_0_io_rPort_5_output_0; // @[Math.scala 263:17:@63920.4]
  assign x645_1_io_b = 32'h1; // @[Math.scala 264:17:@63921.4]
  assign x645_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63922.4]
  assign x646_1_clock = clock; // @[:@63930.4]
  assign x646_1_io_a = x384_lb2_0_io_rPort_4_output_0; // @[Math.scala 263:17:@63932.4]
  assign x646_1_io_b = 32'h2; // @[Math.scala 264:17:@63933.4]
  assign x646_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63934.4]
  assign x647_1_clock = clock; // @[:@63942.4]
  assign x647_1_io_a = x384_lb2_0_io_rPort_0_output_0; // @[Math.scala 263:17:@63944.4]
  assign x647_1_io_b = 32'h4; // @[Math.scala 264:17:@63945.4]
  assign x647_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63946.4]
  assign x648_1_clock = clock; // @[:@63954.4]
  assign x648_1_io_a = x384_lb2_0_io_rPort_6_output_0; // @[Math.scala 263:17:@63956.4]
  assign x648_1_io_b = 32'h1; // @[Math.scala 264:17:@63957.4]
  assign x648_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@63958.4]
  assign x649_x9_1_clock = clock; // @[:@63964.4]
  assign x649_x9_1_reset = reset; // @[:@63965.4]
  assign x649_x9_1_io_a = x645_1_io_result; // @[Math.scala 151:17:@63966.4]
  assign x649_x9_1_io_b = x646_1_io_result; // @[Math.scala 152:17:@63967.4]
  assign x649_x9_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63968.4]
  assign x650_x10_1_clock = clock; // @[:@63976.4]
  assign x650_x10_1_reset = reset; // @[:@63977.4]
  assign x650_x10_1_io_a = x647_1_io_result; // @[Math.scala 151:17:@63978.4]
  assign x650_x10_1_io_b = x648_1_io_result; // @[Math.scala 152:17:@63979.4]
  assign x650_x10_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63980.4]
  assign x651_sum_1_clock = clock; // @[:@63986.4]
  assign x651_sum_1_reset = reset; // @[:@63987.4]
  assign x651_sum_1_io_a = x649_x9_1_io_result; // @[Math.scala 151:17:@63988.4]
  assign x651_sum_1_io_b = x650_x10_1_io_result; // @[Math.scala 152:17:@63989.4]
  assign x651_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@63990.4]
  assign x652_1_io_b = x651_sum_1_io_result; // @[Math.scala 721:17:@63998.4]
  assign x653_mul_1_clock = clock; // @[:@64007.4]
  assign x653_mul_1_io_a = x652_1_io_result; // @[Math.scala 263:17:@64009.4]
  assign x653_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@64010.4]
  assign x653_mul_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@64011.4]
  assign x654_1_io_b = x653_mul_1_io_result; // @[Math.scala 721:17:@64019.4]
  assign x655_1_clock = clock; // @[:@64028.4]
  assign x655_1_io_a = x384_lb2_0_io_rPort_4_output_0; // @[Math.scala 263:17:@64030.4]
  assign x655_1_io_b = 32'h1; // @[Math.scala 264:17:@64031.4]
  assign x655_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@64032.4]
  assign x656_1_clock = clock; // @[:@64040.4]
  assign x656_1_io_a = x384_lb2_0_io_rPort_8_output_0; // @[Math.scala 263:17:@64042.4]
  assign x656_1_io_b = 32'h2; // @[Math.scala 264:17:@64043.4]
  assign x656_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@64044.4]
  assign x657_1_clock = clock; // @[:@64052.4]
  assign x657_1_io_a = x384_lb2_0_io_rPort_6_output_0; // @[Math.scala 263:17:@64054.4]
  assign x657_1_io_b = 32'h4; // @[Math.scala 264:17:@64055.4]
  assign x657_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@64056.4]
  assign x658_1_clock = clock; // @[:@64064.4]
  assign x658_1_io_a = x384_lb2_0_io_rPort_1_output_0; // @[Math.scala 263:17:@64066.4]
  assign x658_1_io_b = 32'h1; // @[Math.scala 264:17:@64067.4]
  assign x658_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@64068.4]
  assign x659_x9_1_clock = clock; // @[:@64074.4]
  assign x659_x9_1_reset = reset; // @[:@64075.4]
  assign x659_x9_1_io_a = x655_1_io_result; // @[Math.scala 151:17:@64076.4]
  assign x659_x9_1_io_b = x656_1_io_result; // @[Math.scala 152:17:@64077.4]
  assign x659_x9_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@64078.4]
  assign x660_x10_1_clock = clock; // @[:@64084.4]
  assign x660_x10_1_reset = reset; // @[:@64085.4]
  assign x660_x10_1_io_a = x657_1_io_result; // @[Math.scala 151:17:@64086.4]
  assign x660_x10_1_io_b = x658_1_io_result; // @[Math.scala 152:17:@64087.4]
  assign x660_x10_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@64088.4]
  assign x661_sum_1_clock = clock; // @[:@64094.4]
  assign x661_sum_1_reset = reset; // @[:@64095.4]
  assign x661_sum_1_io_a = x659_x9_1_io_result; // @[Math.scala 151:17:@64096.4]
  assign x661_sum_1_io_b = x660_x10_1_io_result; // @[Math.scala 152:17:@64097.4]
  assign x661_sum_1_io_flow = io_in_x343_TREADY; // @[Math.scala 153:20:@64098.4]
  assign x662_1_io_b = x661_sum_1_io_result; // @[Math.scala 721:17:@64106.4]
  assign x663_mul_1_clock = clock; // @[:@64115.4]
  assign x663_mul_1_io_a = x662_1_io_result; // @[Math.scala 263:17:@64117.4]
  assign x663_mul_1_io_b = 32'h10; // @[Math.scala 264:17:@64118.4]
  assign x663_mul_1_io_flow = io_in_x343_TREADY; // @[Math.scala 265:20:@64119.4]
  assign x664_1_io_b = x663_mul_1_io_result; // @[Math.scala 721:17:@64127.4]
  assign RetimeWrapper_166_clock = clock; // @[:@64144.4]
  assign RetimeWrapper_166_reset = reset; // @[:@64145.4]
  assign RetimeWrapper_166_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@64147.4]
  assign RetimeWrapper_166_io_in = {_T_2361,_T_2360}; // @[package.scala 94:16:@64146.4]
  assign RetimeWrapper_167_clock = clock; // @[:@64153.4]
  assign RetimeWrapper_167_reset = reset; // @[:@64154.4]
  assign RetimeWrapper_167_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@64156.4]
  assign RetimeWrapper_167_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@64155.4]
  assign RetimeWrapper_168_clock = clock; // @[:@64162.4]
  assign RetimeWrapper_168_reset = reset; // @[:@64163.4]
  assign RetimeWrapper_168_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@64165.4]
  assign RetimeWrapper_168_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@64164.4]
  assign RetimeWrapper_169_clock = clock; // @[:@64171.4]
  assign RetimeWrapper_169_reset = reset; // @[:@64172.4]
  assign RetimeWrapper_169_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@64174.4]
  assign RetimeWrapper_169_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@64173.4]
endmodule
module x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1( // @[:@64192.2]
  input          clock, // @[:@64193.4]
  input          reset, // @[:@64194.4]
  output         io_in_x343_TVALID, // @[:@64195.4]
  input          io_in_x343_TREADY, // @[:@64195.4]
  output [255:0] io_in_x343_TDATA, // @[:@64195.4]
  input          io_in_x342_TVALID, // @[:@64195.4]
  output         io_in_x342_TREADY, // @[:@64195.4]
  input  [255:0] io_in_x342_TDATA, // @[:@64195.4]
  input  [7:0]   io_in_x342_TID, // @[:@64195.4]
  input  [7:0]   io_in_x342_TDEST, // @[:@64195.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@64195.4]
  input          io_sigsIn_smChildAcks_0, // @[:@64195.4]
  output         io_sigsOut_smDoneIn_0, // @[:@64195.4]
  input          io_rr // @[:@64195.4]
);
  wire  x376_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire  x376_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire  x376_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire  x376_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire [12:0] x376_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire [12:0] x376_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire  x376_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire  x376_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire  x376_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@64229.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@64317.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@64317.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@64317.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@64317.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@64317.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@64359.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@64359.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@64359.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@64359.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@64359.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@64367.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@64367.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@64367.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@64367.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@64367.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TVALID; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TREADY; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire [255:0] x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TDATA; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TREADY; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire [255:0] x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TDATA; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire [7:0] x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TID; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire [7:0] x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TDEST; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire [31:0] x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire [31:0] x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
  wire  _T_240; // @[package.scala 96:25:@64322.4 package.scala 96:25:@64323.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x670_outr_UnitPipe.scala 69:66:@64328.4]
  wire  _T_253; // @[package.scala 96:25:@64364.4 package.scala 96:25:@64365.4]
  wire  _T_259; // @[package.scala 96:25:@64372.4 package.scala 96:25:@64373.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@64375.4]
  wire  x669_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@64376.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@64384.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@64385.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@64397.4]
  x350_ctrchain x376_ctrchain ( // @[SpatialBlocks.scala 37:22:@64229.4]
    .clock(x376_ctrchain_clock),
    .reset(x376_ctrchain_reset),
    .io_input_reset(x376_ctrchain_io_input_reset),
    .io_input_enable(x376_ctrchain_io_input_enable),
    .io_output_counts_1(x376_ctrchain_io_output_counts_1),
    .io_output_counts_0(x376_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x376_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x376_ctrchain_io_output_oobs_1),
    .io_output_done(x376_ctrchain_io_output_done)
  );
  x669_inr_Foreach_SAMPLER_BOX_sm x669_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 32:18:@64289.4]
    .clock(x669_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x669_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x669_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x669_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x669_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x669_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x669_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x669_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x669_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@64317.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@64359.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@64367.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1 x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1073:24:@64401.4]
    .clock(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x343_TVALID(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TVALID),
    .io_in_x343_TREADY(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TREADY),
    .io_in_x343_TDATA(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TDATA),
    .io_in_x342_TREADY(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TREADY),
    .io_in_x342_TDATA(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TDATA),
    .io_in_x342_TID(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TID),
    .io_in_x342_TDEST(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TDEST),
    .io_sigsIn_backpressure(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@64322.4 package.scala 96:25:@64323.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x342_TVALID | x669_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x670_outr_UnitPipe.scala 69:66:@64328.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@64364.4 package.scala 96:25:@64365.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@64372.4 package.scala 96:25:@64373.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@64375.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@64376.4]
  assign _T_264 = x669_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@64384.4]
  assign _T_265 = ~ x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@64385.4]
  assign _T_272 = x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@64397.4]
  assign io_in_x343_TVALID = x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TVALID; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 48:23:@64460.4]
  assign io_in_x343_TDATA = x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TDATA; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 48:23:@64458.4]
  assign io_in_x342_TREADY = x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TREADY; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 49:23:@64468.4]
  assign io_sigsOut_smDoneIn_0 = x669_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@64382.4]
  assign x376_ctrchain_clock = clock; // @[:@64230.4]
  assign x376_ctrchain_reset = reset; // @[:@64231.4]
  assign x376_ctrchain_io_input_reset = x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@64400.4]
  assign x376_ctrchain_io_input_enable = _T_272 & x669_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@64352.4 SpatialBlocks.scala 159:42:@64399.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@64290.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@64291.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sm_io_enable = x669_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x669_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@64379.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x670_outr_UnitPipe.scala 67:50:@64325.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@64381.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x343_TREADY | x669_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@64353.4]
  assign x669_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x670_outr_UnitPipe.scala 71:48:@64331.4]
  assign RetimeWrapper_clock = clock; // @[:@64318.4]
  assign RetimeWrapper_reset = reset; // @[:@64319.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@64321.4]
  assign RetimeWrapper_io_in = x376_ctrchain_io_output_done; // @[package.scala 94:16:@64320.4]
  assign RetimeWrapper_1_clock = clock; // @[:@64360.4]
  assign RetimeWrapper_1_reset = reset; // @[:@64361.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@64363.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@64362.4]
  assign RetimeWrapper_2_clock = clock; // @[:@64368.4]
  assign RetimeWrapper_2_reset = reset; // @[:@64369.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@64371.4]
  assign RetimeWrapper_2_io_in = x669_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@64370.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@64402.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@64403.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x343_TREADY = io_in_x343_TREADY; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 48:23:@64459.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TDATA = io_in_x342_TDATA; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 49:23:@64467.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TID = io_in_x342_TID; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 49:23:@64463.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x342_TDEST = io_in_x342_TDEST; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 49:23:@64462.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x343_TREADY | x669_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1078:22:@64486.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1078:22:@64484.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x669_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1078:22:@64482.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x376_ctrchain_io_output_counts_1[12]}},x376_ctrchain_io_output_counts_1}; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1078:22:@64477.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x376_ctrchain_io_output_counts_0[12]}},x376_ctrchain_io_output_counts_0}; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1078:22:@64476.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x376_ctrchain_io_output_oobs_0; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1078:22:@64474.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x376_ctrchain_io_output_oobs_1; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1078:22:@64475.4]
  assign x669_inr_Foreach_SAMPLER_BOX_kernelx669_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x669_inr_Foreach_SAMPLER_BOX.scala 1077:18:@64470.4]
endmodule
module x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1( // @[:@64500.2]
  input          clock, // @[:@64501.4]
  input          reset, // @[:@64502.4]
  output         io_in_x343_TVALID, // @[:@64503.4]
  input          io_in_x343_TREADY, // @[:@64503.4]
  output [255:0] io_in_x343_TDATA, // @[:@64503.4]
  input          io_in_x342_TVALID, // @[:@64503.4]
  output         io_in_x342_TREADY, // @[:@64503.4]
  input  [255:0] io_in_x342_TDATA, // @[:@64503.4]
  input  [7:0]   io_in_x342_TID, // @[:@64503.4]
  input  [7:0]   io_in_x342_TDEST, // @[:@64503.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@64503.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@64503.4]
  input          io_sigsIn_smChildAcks_0, // @[:@64503.4]
  input          io_sigsIn_smChildAcks_1, // @[:@64503.4]
  output         io_sigsOut_smDoneIn_0, // @[:@64503.4]
  output         io_sigsOut_smDoneIn_1, // @[:@64503.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@64503.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@64503.4]
  input          io_rr // @[:@64503.4]
);
  wire  x345_fifoinraw_0_clock; // @[m_x345_fifoinraw_0.scala 27:17:@64517.4]
  wire  x345_fifoinraw_0_reset; // @[m_x345_fifoinraw_0.scala 27:17:@64517.4]
  wire  x346_fifoinpacked_0_clock; // @[m_x346_fifoinpacked_0.scala 27:17:@64541.4]
  wire  x346_fifoinpacked_0_reset; // @[m_x346_fifoinpacked_0.scala 27:17:@64541.4]
  wire  x346_fifoinpacked_0_io_wPort_0_en_0; // @[m_x346_fifoinpacked_0.scala 27:17:@64541.4]
  wire  x346_fifoinpacked_0_io_full; // @[m_x346_fifoinpacked_0.scala 27:17:@64541.4]
  wire  x346_fifoinpacked_0_io_active_0_in; // @[m_x346_fifoinpacked_0.scala 27:17:@64541.4]
  wire  x346_fifoinpacked_0_io_active_0_out; // @[m_x346_fifoinpacked_0.scala 27:17:@64541.4]
  wire  x347_fifooutraw_0_clock; // @[m_x347_fifooutraw_0.scala 27:17:@64565.4]
  wire  x347_fifooutraw_0_reset; // @[m_x347_fifooutraw_0.scala 27:17:@64565.4]
  wire  x350_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire  x350_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire  x350_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire  x350_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire [12:0] x350_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire [12:0] x350_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire  x350_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire  x350_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire  x350_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@64589.4]
  wire  x372_inr_Foreach_sm_clock; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_reset; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_enable; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_done; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_doneLatch; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_ctrDone; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_datapathEn; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_ctrInc; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_ctrRst; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_parentAck; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_backpressure; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  x372_inr_Foreach_sm_io_break; // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@64677.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@64677.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@64677.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@64677.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@64677.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@64723.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@64723.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@64723.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@64723.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@64723.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@64731.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@64731.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@64731.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@64731.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@64731.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_clock; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_reset; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_wPort_0_en_0; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_full; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_active_0_in; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_active_0_out; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire [31:0] x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire [31:0] x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_rr; // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
  wire  x670_outr_UnitPipe_sm_clock; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_reset; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_enable; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_done; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_rst; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_ctrDone; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_ctrInc; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_parentAck; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  x670_outr_UnitPipe_sm_io_childAck_0; // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@64955.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@64955.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@64955.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@64955.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@64955.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@64963.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@64963.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@64963.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@64963.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@64963.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_clock; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_reset; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TVALID; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TREADY; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire [255:0] x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TDATA; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TVALID; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TREADY; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire [255:0] x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TDATA; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire [7:0] x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TID; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire [7:0] x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TDEST; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_rr; // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
  wire  _T_254; // @[package.scala 96:25:@64682.4 package.scala 96:25:@64683.4]
  wire  _T_260; // @[implicits.scala 47:10:@64686.4]
  wire  _T_261; // @[sm_x671_outr_UnitPipe.scala 70:41:@64687.4]
  wire  _T_262; // @[sm_x671_outr_UnitPipe.scala 70:78:@64688.4]
  wire  _T_263; // @[sm_x671_outr_UnitPipe.scala 70:76:@64689.4]
  wire  _T_275; // @[package.scala 96:25:@64728.4 package.scala 96:25:@64729.4]
  wire  _T_281; // @[package.scala 96:25:@64736.4 package.scala 96:25:@64737.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@64739.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@64748.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@64749.4]
  wire  _T_354; // @[package.scala 100:49:@64926.4]
  reg  _T_357; // @[package.scala 48:56:@64927.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@64960.4 package.scala 96:25:@64961.4]
  wire  _T_377; // @[package.scala 96:25:@64968.4 package.scala 96:25:@64969.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@64971.4]
  x345_fifoinraw_0 x345_fifoinraw_0 ( // @[m_x345_fifoinraw_0.scala 27:17:@64517.4]
    .clock(x345_fifoinraw_0_clock),
    .reset(x345_fifoinraw_0_reset)
  );
  x346_fifoinpacked_0 x346_fifoinpacked_0 ( // @[m_x346_fifoinpacked_0.scala 27:17:@64541.4]
    .clock(x346_fifoinpacked_0_clock),
    .reset(x346_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x346_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x346_fifoinpacked_0_io_full),
    .io_active_0_in(x346_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x346_fifoinpacked_0_io_active_0_out)
  );
  x345_fifoinraw_0 x347_fifooutraw_0 ( // @[m_x347_fifooutraw_0.scala 27:17:@64565.4]
    .clock(x347_fifooutraw_0_clock),
    .reset(x347_fifooutraw_0_reset)
  );
  x350_ctrchain x350_ctrchain ( // @[SpatialBlocks.scala 37:22:@64589.4]
    .clock(x350_ctrchain_clock),
    .reset(x350_ctrchain_reset),
    .io_input_reset(x350_ctrchain_io_input_reset),
    .io_input_enable(x350_ctrchain_io_input_enable),
    .io_output_counts_1(x350_ctrchain_io_output_counts_1),
    .io_output_counts_0(x350_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x350_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x350_ctrchain_io_output_oobs_1),
    .io_output_done(x350_ctrchain_io_output_done)
  );
  x372_inr_Foreach_sm x372_inr_Foreach_sm ( // @[sm_x372_inr_Foreach.scala 32:18:@64649.4]
    .clock(x372_inr_Foreach_sm_clock),
    .reset(x372_inr_Foreach_sm_reset),
    .io_enable(x372_inr_Foreach_sm_io_enable),
    .io_done(x372_inr_Foreach_sm_io_done),
    .io_doneLatch(x372_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x372_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x372_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x372_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x372_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x372_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x372_inr_Foreach_sm_io_backpressure),
    .io_break(x372_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@64677.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@64723.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@64731.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x372_inr_Foreach_kernelx372_inr_Foreach_concrete1 x372_inr_Foreach_kernelx372_inr_Foreach_concrete1 ( // @[sm_x372_inr_Foreach.scala 110:24:@64766.4]
    .clock(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_clock),
    .reset(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_reset),
    .io_in_x346_fifoinpacked_0_wPort_0_en_0(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_wPort_0_en_0),
    .io_in_x346_fifoinpacked_0_full(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_full),
    .io_in_x346_fifoinpacked_0_active_0_in(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_active_0_in),
    .io_in_x346_fifoinpacked_0_active_0_out(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x670_outr_UnitPipe_sm ( // @[sm_x670_outr_UnitPipe.scala 32:18:@64898.4]
    .clock(x670_outr_UnitPipe_sm_clock),
    .reset(x670_outr_UnitPipe_sm_reset),
    .io_enable(x670_outr_UnitPipe_sm_io_enable),
    .io_done(x670_outr_UnitPipe_sm_io_done),
    .io_rst(x670_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x670_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x670_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x670_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x670_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x670_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x670_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@64955.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@64963.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1 x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1 ( // @[sm_x670_outr_UnitPipe.scala 76:24:@64993.4]
    .clock(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_clock),
    .reset(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_reset),
    .io_in_x343_TVALID(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TVALID),
    .io_in_x343_TREADY(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TREADY),
    .io_in_x343_TDATA(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TDATA),
    .io_in_x342_TVALID(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TVALID),
    .io_in_x342_TREADY(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TREADY),
    .io_in_x342_TDATA(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TDATA),
    .io_in_x342_TID(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TID),
    .io_in_x342_TDEST(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TDEST),
    .io_sigsIn_smEnableOuts_0(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@64682.4 package.scala 96:25:@64683.4]
  assign _T_260 = x346_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@64686.4]
  assign _T_261 = ~ _T_260; // @[sm_x671_outr_UnitPipe.scala 70:41:@64687.4]
  assign _T_262 = ~ x346_fifoinpacked_0_io_active_0_out; // @[sm_x671_outr_UnitPipe.scala 70:78:@64688.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x671_outr_UnitPipe.scala 70:76:@64689.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@64728.4 package.scala 96:25:@64729.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@64736.4 package.scala 96:25:@64737.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@64739.4]
  assign _T_286 = x372_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@64748.4]
  assign _T_287 = ~ x372_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@64749.4]
  assign _T_354 = x670_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@64926.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@64960.4 package.scala 96:25:@64961.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@64968.4 package.scala 96:25:@64969.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@64971.4]
  assign io_in_x343_TVALID = x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TVALID; // @[sm_x670_outr_UnitPipe.scala 48:23:@65050.4]
  assign io_in_x343_TDATA = x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TDATA; // @[sm_x670_outr_UnitPipe.scala 48:23:@65048.4]
  assign io_in_x342_TREADY = x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TREADY; // @[sm_x670_outr_UnitPipe.scala 49:23:@65058.4]
  assign io_sigsOut_smDoneIn_0 = x372_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@64746.4]
  assign io_sigsOut_smDoneIn_1 = x670_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@64978.4]
  assign io_sigsOut_smCtrCopyDone_0 = x372_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@64765.4]
  assign io_sigsOut_smCtrCopyDone_1 = x670_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@64992.4]
  assign x345_fifoinraw_0_clock = clock; // @[:@64518.4]
  assign x345_fifoinraw_0_reset = reset; // @[:@64519.4]
  assign x346_fifoinpacked_0_clock = clock; // @[:@64542.4]
  assign x346_fifoinpacked_0_reset = reset; // @[:@64543.4]
  assign x346_fifoinpacked_0_io_wPort_0_en_0 = x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@64826.4]
  assign x346_fifoinpacked_0_io_active_0_in = x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@64825.4]
  assign x347_fifooutraw_0_clock = clock; // @[:@64566.4]
  assign x347_fifooutraw_0_reset = reset; // @[:@64567.4]
  assign x350_ctrchain_clock = clock; // @[:@64590.4]
  assign x350_ctrchain_reset = reset; // @[:@64591.4]
  assign x350_ctrchain_io_input_reset = x372_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@64764.4]
  assign x350_ctrchain_io_input_enable = x372_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@64716.4 SpatialBlocks.scala 159:42:@64763.4]
  assign x372_inr_Foreach_sm_clock = clock; // @[:@64650.4]
  assign x372_inr_Foreach_sm_reset = reset; // @[:@64651.4]
  assign x372_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@64743.4]
  assign x372_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x671_outr_UnitPipe.scala 69:38:@64685.4]
  assign x372_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@64745.4]
  assign x372_inr_Foreach_sm_io_backpressure = _T_263 | x372_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@64717.4]
  assign x372_inr_Foreach_sm_io_break = 1'h0; // @[sm_x671_outr_UnitPipe.scala 73:36:@64695.4]
  assign RetimeWrapper_clock = clock; // @[:@64678.4]
  assign RetimeWrapper_reset = reset; // @[:@64679.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@64681.4]
  assign RetimeWrapper_io_in = x350_ctrchain_io_output_done; // @[package.scala 94:16:@64680.4]
  assign RetimeWrapper_1_clock = clock; // @[:@64724.4]
  assign RetimeWrapper_1_reset = reset; // @[:@64725.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@64727.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@64726.4]
  assign RetimeWrapper_2_clock = clock; // @[:@64732.4]
  assign RetimeWrapper_2_reset = reset; // @[:@64733.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@64735.4]
  assign RetimeWrapper_2_io_in = x372_inr_Foreach_sm_io_done; // @[package.scala 94:16:@64734.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_clock = clock; // @[:@64767.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_reset = reset; // @[:@64768.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_full = x346_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@64820.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_in_x346_fifoinpacked_0_active_0_out = x346_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@64819.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x372_inr_Foreach_sm_io_doneLatch; // @[sm_x372_inr_Foreach.scala 115:22:@64849.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x372_inr_Foreach.scala 115:22:@64847.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_break = x372_inr_Foreach_sm_io_break; // @[sm_x372_inr_Foreach.scala 115:22:@64845.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x350_ctrchain_io_output_counts_1[12]}},x350_ctrchain_io_output_counts_1}; // @[sm_x372_inr_Foreach.scala 115:22:@64840.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x350_ctrchain_io_output_counts_0[12]}},x350_ctrchain_io_output_counts_0}; // @[sm_x372_inr_Foreach.scala 115:22:@64839.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x350_ctrchain_io_output_oobs_0; // @[sm_x372_inr_Foreach.scala 115:22:@64837.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x350_ctrchain_io_output_oobs_1; // @[sm_x372_inr_Foreach.scala 115:22:@64838.4]
  assign x372_inr_Foreach_kernelx372_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x372_inr_Foreach.scala 114:18:@64833.4]
  assign x670_outr_UnitPipe_sm_clock = clock; // @[:@64899.4]
  assign x670_outr_UnitPipe_sm_reset = reset; // @[:@64900.4]
  assign x670_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@64975.4]
  assign x670_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@64950.4]
  assign x670_outr_UnitPipe_sm_io_ctrDone = x670_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x671_outr_UnitPipe.scala 78:40:@64930.4]
  assign x670_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@64977.4]
  assign x670_outr_UnitPipe_sm_io_doneIn_0 = x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@64947.4]
  assign RetimeWrapper_3_clock = clock; // @[:@64956.4]
  assign RetimeWrapper_3_reset = reset; // @[:@64957.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@64959.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@64958.4]
  assign RetimeWrapper_4_clock = clock; // @[:@64964.4]
  assign RetimeWrapper_4_reset = reset; // @[:@64965.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@64967.4]
  assign RetimeWrapper_4_io_in = x670_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@64966.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_clock = clock; // @[:@64994.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_reset = reset; // @[:@64995.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x343_TREADY = io_in_x343_TREADY; // @[sm_x670_outr_UnitPipe.scala 48:23:@65049.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TVALID = io_in_x342_TVALID; // @[sm_x670_outr_UnitPipe.scala 49:23:@65059.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TDATA = io_in_x342_TDATA; // @[sm_x670_outr_UnitPipe.scala 49:23:@65057.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TID = io_in_x342_TID; // @[sm_x670_outr_UnitPipe.scala 49:23:@65053.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_in_x342_TDEST = io_in_x342_TDEST; // @[sm_x670_outr_UnitPipe.scala 49:23:@65052.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x670_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x670_outr_UnitPipe.scala 81:22:@65068.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x670_outr_UnitPipe_sm_io_childAck_0; // @[sm_x670_outr_UnitPipe.scala 81:22:@65066.4]
  assign x670_outr_UnitPipe_kernelx670_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x670_outr_UnitPipe.scala 80:18:@65060.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x693_outr_UnitPipe_sm( // @[:@65557.2]
  input   clock, // @[:@65558.4]
  input   reset, // @[:@65559.4]
  input   io_enable, // @[:@65560.4]
  output  io_done, // @[:@65560.4]
  input   io_parentAck, // @[:@65560.4]
  input   io_doneIn_0, // @[:@65560.4]
  input   io_doneIn_1, // @[:@65560.4]
  input   io_doneIn_2, // @[:@65560.4]
  output  io_enableOut_0, // @[:@65560.4]
  output  io_enableOut_1, // @[:@65560.4]
  output  io_enableOut_2, // @[:@65560.4]
  output  io_childAck_0, // @[:@65560.4]
  output  io_childAck_1, // @[:@65560.4]
  output  io_childAck_2, // @[:@65560.4]
  input   io_ctrCopyDone_0, // @[:@65560.4]
  input   io_ctrCopyDone_1, // @[:@65560.4]
  input   io_ctrCopyDone_2 // @[:@65560.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@65563.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@65563.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@65563.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@65563.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@65563.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@65563.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@65566.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@65566.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@65566.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@65566.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@65566.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@65566.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@65569.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@65569.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@65569.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@65569.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@65569.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@65569.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@65572.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@65572.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@65572.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@65572.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@65572.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@65572.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@65575.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@65575.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@65575.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@65575.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@65575.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@65575.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@65578.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@65578.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@65578.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@65578.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@65578.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@65578.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@65619.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@65619.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@65619.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@65619.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@65619.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@65619.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@65622.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@65622.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@65622.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@65622.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@65622.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@65622.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@65625.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@65625.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@65625.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@65625.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@65625.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@65625.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@65676.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@65676.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@65676.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@65676.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@65676.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@65690.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@65690.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@65690.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@65690.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@65690.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@65708.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@65708.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@65708.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@65708.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@65708.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@65745.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@65745.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@65745.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@65745.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@65745.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@65759.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@65759.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@65759.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@65759.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@65759.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@65777.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@65777.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@65777.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@65777.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@65777.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@65814.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@65814.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@65814.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@65814.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@65814.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@65828.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@65828.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@65828.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@65828.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@65828.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@65846.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@65846.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@65846.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@65846.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@65846.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@65903.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@65903.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@65903.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@65903.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@65903.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@65920.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@65920.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@65920.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@65920.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@65920.4]
  wire  _T_77; // @[Controllers.scala 80:47:@65581.4]
  wire  allDone; // @[Controllers.scala 80:47:@65582.4]
  wire  _T_151; // @[Controllers.scala 165:35:@65660.4]
  wire  _T_153; // @[Controllers.scala 165:60:@65661.4]
  wire  _T_154; // @[Controllers.scala 165:58:@65662.4]
  wire  _T_156; // @[Controllers.scala 165:76:@65663.4]
  wire  _T_157; // @[Controllers.scala 165:74:@65664.4]
  wire  _T_161; // @[Controllers.scala 165:109:@65667.4]
  wire  _T_164; // @[Controllers.scala 165:141:@65669.4]
  wire  _T_172; // @[package.scala 96:25:@65681.4 package.scala 96:25:@65682.4]
  wire  _T_176; // @[Controllers.scala 167:54:@65684.4]
  wire  _T_177; // @[Controllers.scala 167:52:@65685.4]
  wire  _T_184; // @[package.scala 96:25:@65695.4 package.scala 96:25:@65696.4]
  wire  _T_202; // @[package.scala 96:25:@65713.4 package.scala 96:25:@65714.4]
  wire  _T_206; // @[Controllers.scala 169:67:@65716.4]
  wire  _T_207; // @[Controllers.scala 169:86:@65717.4]
  wire  _T_219; // @[Controllers.scala 165:35:@65729.4]
  wire  _T_221; // @[Controllers.scala 165:60:@65730.4]
  wire  _T_222; // @[Controllers.scala 165:58:@65731.4]
  wire  _T_224; // @[Controllers.scala 165:76:@65732.4]
  wire  _T_225; // @[Controllers.scala 165:74:@65733.4]
  wire  _T_229; // @[Controllers.scala 165:109:@65736.4]
  wire  _T_232; // @[Controllers.scala 165:141:@65738.4]
  wire  _T_240; // @[package.scala 96:25:@65750.4 package.scala 96:25:@65751.4]
  wire  _T_244; // @[Controllers.scala 167:54:@65753.4]
  wire  _T_245; // @[Controllers.scala 167:52:@65754.4]
  wire  _T_252; // @[package.scala 96:25:@65764.4 package.scala 96:25:@65765.4]
  wire  _T_270; // @[package.scala 96:25:@65782.4 package.scala 96:25:@65783.4]
  wire  _T_274; // @[Controllers.scala 169:67:@65785.4]
  wire  _T_275; // @[Controllers.scala 169:86:@65786.4]
  wire  _T_287; // @[Controllers.scala 165:35:@65798.4]
  wire  _T_289; // @[Controllers.scala 165:60:@65799.4]
  wire  _T_290; // @[Controllers.scala 165:58:@65800.4]
  wire  _T_292; // @[Controllers.scala 165:76:@65801.4]
  wire  _T_293; // @[Controllers.scala 165:74:@65802.4]
  wire  _T_297; // @[Controllers.scala 165:109:@65805.4]
  wire  _T_300; // @[Controllers.scala 165:141:@65807.4]
  wire  _T_308; // @[package.scala 96:25:@65819.4 package.scala 96:25:@65820.4]
  wire  _T_312; // @[Controllers.scala 167:54:@65822.4]
  wire  _T_313; // @[Controllers.scala 167:52:@65823.4]
  wire  _T_320; // @[package.scala 96:25:@65833.4 package.scala 96:25:@65834.4]
  wire  _T_338; // @[package.scala 96:25:@65851.4 package.scala 96:25:@65852.4]
  wire  _T_342; // @[Controllers.scala 169:67:@65854.4]
  wire  _T_343; // @[Controllers.scala 169:86:@65855.4]
  wire  _T_358; // @[Controllers.scala 213:68:@65873.4]
  wire  _T_360; // @[Controllers.scala 213:90:@65875.4]
  wire  _T_362; // @[Controllers.scala 213:132:@65877.4]
  wire  _T_366; // @[Controllers.scala 213:68:@65882.4]
  wire  _T_368; // @[Controllers.scala 213:90:@65884.4]
  wire  _T_374; // @[Controllers.scala 213:68:@65890.4]
  wire  _T_376; // @[Controllers.scala 213:90:@65892.4]
  wire  _T_383; // @[package.scala 100:49:@65898.4]
  reg  _T_386; // @[package.scala 48:56:@65899.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@65901.4]
  reg  _T_400; // @[package.scala 48:56:@65917.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@65563.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@65566.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@65569.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@65572.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@65575.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@65578.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@65619.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@65622.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@65625.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@65676.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@65690.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@65708.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@65745.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@65759.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@65777.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@65814.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@65828.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@65846.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@65903.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@65920.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@65581.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@65582.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@65660.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@65661.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@65662.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@65663.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@65664.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@65667.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@65669.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@65681.4 package.scala 96:25:@65682.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@65684.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@65685.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@65695.4 package.scala 96:25:@65696.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@65713.4 package.scala 96:25:@65714.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@65716.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@65717.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@65729.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@65730.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@65731.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@65732.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@65733.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@65736.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@65738.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@65750.4 package.scala 96:25:@65751.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@65753.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@65754.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@65764.4 package.scala 96:25:@65765.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@65782.4 package.scala 96:25:@65783.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@65785.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@65786.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@65798.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@65799.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@65800.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@65801.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@65802.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@65805.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@65807.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@65819.4 package.scala 96:25:@65820.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@65822.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@65823.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@65833.4 package.scala 96:25:@65834.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@65851.4 package.scala 96:25:@65852.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@65854.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@65855.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@65873.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@65875.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@65877.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@65882.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@65884.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@65890.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@65892.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@65898.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@65901.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@65927.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@65881.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@65889.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@65897.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@65868.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@65870.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@65872.4]
  assign active_0_clock = clock; // @[:@65564.4]
  assign active_0_reset = reset; // @[:@65565.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@65671.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@65675.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@65585.4]
  assign active_1_clock = clock; // @[:@65567.4]
  assign active_1_reset = reset; // @[:@65568.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@65740.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@65744.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@65586.4]
  assign active_2_clock = clock; // @[:@65570.4]
  assign active_2_reset = reset; // @[:@65571.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@65809.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@65813.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@65587.4]
  assign done_0_clock = clock; // @[:@65573.4]
  assign done_0_reset = reset; // @[:@65574.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@65721.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@65599.4 Controllers.scala 170:32:@65728.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@65588.4]
  assign done_1_clock = clock; // @[:@65576.4]
  assign done_1_reset = reset; // @[:@65577.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@65790.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@65608.4 Controllers.scala 170:32:@65797.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@65589.4]
  assign done_2_clock = clock; // @[:@65579.4]
  assign done_2_reset = reset; // @[:@65580.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@65859.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@65617.4 Controllers.scala 170:32:@65866.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@65590.4]
  assign iterDone_0_clock = clock; // @[:@65620.4]
  assign iterDone_0_reset = reset; // @[:@65621.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@65689.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@65639.4 Controllers.scala 168:36:@65705.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@65628.4]
  assign iterDone_1_clock = clock; // @[:@65623.4]
  assign iterDone_1_reset = reset; // @[:@65624.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@65758.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@65648.4 Controllers.scala 168:36:@65774.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@65629.4]
  assign iterDone_2_clock = clock; // @[:@65626.4]
  assign iterDone_2_reset = reset; // @[:@65627.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@65827.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@65657.4 Controllers.scala 168:36:@65843.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@65630.4]
  assign RetimeWrapper_clock = clock; // @[:@65677.4]
  assign RetimeWrapper_reset = reset; // @[:@65678.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@65680.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@65679.4]
  assign RetimeWrapper_1_clock = clock; // @[:@65691.4]
  assign RetimeWrapper_1_reset = reset; // @[:@65692.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@65694.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@65693.4]
  assign RetimeWrapper_2_clock = clock; // @[:@65709.4]
  assign RetimeWrapper_2_reset = reset; // @[:@65710.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@65712.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@65711.4]
  assign RetimeWrapper_3_clock = clock; // @[:@65746.4]
  assign RetimeWrapper_3_reset = reset; // @[:@65747.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@65749.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@65748.4]
  assign RetimeWrapper_4_clock = clock; // @[:@65760.4]
  assign RetimeWrapper_4_reset = reset; // @[:@65761.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@65763.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@65762.4]
  assign RetimeWrapper_5_clock = clock; // @[:@65778.4]
  assign RetimeWrapper_5_reset = reset; // @[:@65779.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@65781.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@65780.4]
  assign RetimeWrapper_6_clock = clock; // @[:@65815.4]
  assign RetimeWrapper_6_reset = reset; // @[:@65816.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@65818.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@65817.4]
  assign RetimeWrapper_7_clock = clock; // @[:@65829.4]
  assign RetimeWrapper_7_reset = reset; // @[:@65830.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@65832.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@65831.4]
  assign RetimeWrapper_8_clock = clock; // @[:@65847.4]
  assign RetimeWrapper_8_reset = reset; // @[:@65848.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@65850.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@65849.4]
  assign RetimeWrapper_9_clock = clock; // @[:@65904.4]
  assign RetimeWrapper_9_reset = reset; // @[:@65905.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@65907.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@65906.4]
  assign RetimeWrapper_10_clock = clock; // @[:@65921.4]
  assign RetimeWrapper_10_reset = reset; // @[:@65922.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@65924.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@65923.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x679_inr_UnitPipe_sm( // @[:@66100.2]
  input   clock, // @[:@66101.4]
  input   reset, // @[:@66102.4]
  input   io_enable, // @[:@66103.4]
  output  io_done, // @[:@66103.4]
  output  io_doneLatch, // @[:@66103.4]
  input   io_ctrDone, // @[:@66103.4]
  output  io_datapathEn, // @[:@66103.4]
  output  io_ctrInc, // @[:@66103.4]
  input   io_parentAck, // @[:@66103.4]
  input   io_backpressure // @[:@66103.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@66105.4]
  wire  active_reset; // @[Controllers.scala 261:22:@66105.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@66105.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@66105.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@66105.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@66105.4]
  wire  done_clock; // @[Controllers.scala 262:20:@66108.4]
  wire  done_reset; // @[Controllers.scala 262:20:@66108.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@66108.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@66108.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@66108.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@66108.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@66162.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@66162.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@66162.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@66162.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@66162.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@66170.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@66170.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@66170.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@66170.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@66170.4]
  wire  _T_80; // @[Controllers.scala 264:48:@66113.4]
  wire  _T_81; // @[Controllers.scala 264:46:@66114.4]
  wire  _T_82; // @[Controllers.scala 264:62:@66115.4]
  wire  _T_83; // @[Controllers.scala 264:60:@66116.4]
  wire  _T_100; // @[package.scala 100:49:@66133.4]
  reg  _T_103; // @[package.scala 48:56:@66134.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@66142.4]
  wire  _T_116; // @[Controllers.scala 283:41:@66150.4]
  wire  _T_117; // @[Controllers.scala 283:59:@66151.4]
  wire  _T_119; // @[Controllers.scala 284:37:@66154.4]
  reg  _T_125; // @[package.scala 48:56:@66158.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@66180.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@66183.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@66185.4]
  wire  _T_152; // @[Controllers.scala 292:61:@66186.4]
  wire  _T_153; // @[Controllers.scala 292:24:@66187.4]
  SRFF active ( // @[Controllers.scala 261:22:@66105.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@66108.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@66162.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@66170.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@66113.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@66114.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@66115.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@66116.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@66133.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@66142.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@66150.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@66151.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@66154.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@66185.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@66186.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@66187.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@66161.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@66189.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@66153.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@66156.4]
  assign active_clock = clock; // @[:@66106.4]
  assign active_reset = reset; // @[:@66107.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@66118.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@66122.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@66123.4]
  assign done_clock = clock; // @[:@66109.4]
  assign done_reset = reset; // @[:@66110.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@66138.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@66131.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@66132.4]
  assign RetimeWrapper_clock = clock; // @[:@66163.4]
  assign RetimeWrapper_reset = reset; // @[:@66164.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@66166.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@66165.4]
  assign RetimeWrapper_1_clock = clock; // @[:@66171.4]
  assign RetimeWrapper_1_reset = reset; // @[:@66172.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@66174.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@66173.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1( // @[:@66264.2]
  input  [63:0] io_in_x340_outdram_number, // @[:@66267.4]
  output        io_in_x672_valid, // @[:@66267.4]
  output [63:0] io_in_x672_bits_addr, // @[:@66267.4]
  output [31:0] io_in_x672_bits_size, // @[:@66267.4]
  input         io_sigsIn_backpressure, // @[:@66267.4]
  input         io_sigsIn_datapathEn, // @[:@66267.4]
  input         io_rr // @[:@66267.4]
);
  wire [96:0] x676_tuple; // @[Cat.scala 30:58:@66281.4]
  wire  _T_135; // @[implicits.scala 55:10:@66284.4]
  assign x676_tuple = {33'h7e9000,io_in_x340_outdram_number}; // @[Cat.scala 30:58:@66281.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@66284.4]
  assign io_in_x672_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x679_inr_UnitPipe.scala 65:18:@66287.4]
  assign io_in_x672_bits_addr = x676_tuple[63:0]; // @[sm_x679_inr_UnitPipe.scala 66:22:@66289.4]
  assign io_in_x672_bits_size = x676_tuple[95:64]; // @[sm_x679_inr_UnitPipe.scala 67:22:@66291.4]
endmodule
module FF_13( // @[:@66293.2]
  input         clock, // @[:@66294.4]
  input         reset, // @[:@66295.4]
  output [22:0] io_rPort_0_output_0, // @[:@66296.4]
  input  [22:0] io_wPort_0_data_0, // @[:@66296.4]
  input         io_wPort_0_reset, // @[:@66296.4]
  input         io_wPort_0_en_0 // @[:@66296.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@66311.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@66313.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@66314.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@66313.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@66314.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@66316.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@66331.2]
  input         clock, // @[:@66332.4]
  input         reset, // @[:@66333.4]
  input         io_input_reset, // @[:@66334.4]
  input         io_input_enable, // @[:@66334.4]
  output [22:0] io_output_count_0, // @[:@66334.4]
  output        io_output_oobs_0, // @[:@66334.4]
  output        io_output_done // @[:@66334.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@66347.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@66347.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@66347.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@66347.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@66347.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@66347.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@66363.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@66363.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@66363.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@66363.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@66363.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@66363.4]
  wire  _T_36; // @[Counter.scala 264:45:@66366.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@66391.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@66392.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@66393.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@66394.4]
  wire  _T_57; // @[Counter.scala 293:18:@66396.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@66404.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@66407.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@66408.4]
  wire  _T_75; // @[Counter.scala 322:102:@66412.4]
  wire  _T_77; // @[Counter.scala 322:130:@66413.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@66347.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@66363.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@66366.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@66391.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@66392.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@66393.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@66394.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@66396.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@66404.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@66407.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@66408.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@66412.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@66413.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@66411.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@66415.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@66417.4]
  assign bases_0_clock = clock; // @[:@66348.4]
  assign bases_0_reset = reset; // @[:@66349.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@66410.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@66389.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@66390.4]
  assign SRFF_clock = clock; // @[:@66364.4]
  assign SRFF_reset = reset; // @[:@66365.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@66368.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@66370.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@66371.4]
endmodule
module x681_ctrchain( // @[:@66422.2]
  input         clock, // @[:@66423.4]
  input         reset, // @[:@66424.4]
  input         io_input_reset, // @[:@66425.4]
  input         io_input_enable, // @[:@66425.4]
  output [22:0] io_output_counts_0, // @[:@66425.4]
  output        io_output_oobs_0, // @[:@66425.4]
  output        io_output_done // @[:@66425.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@66427.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@66427.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@66427.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@66427.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@66427.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@66427.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@66427.4]
  reg  wasDone; // @[Counter.scala 542:24:@66436.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@66442.4]
  wire  _T_47; // @[Counter.scala 546:80:@66443.4]
  reg  doneLatch; // @[Counter.scala 550:26:@66448.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@66449.4]
  wire  _T_55; // @[Counter.scala 551:19:@66450.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@66427.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@66442.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@66443.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@66449.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@66450.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@66452.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@66454.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@66445.4]
  assign ctrs_0_clock = clock; // @[:@66428.4]
  assign ctrs_0_reset = reset; // @[:@66429.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@66433.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@66434.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x688_inr_Foreach_sm( // @[:@66642.2]
  input   clock, // @[:@66643.4]
  input   reset, // @[:@66644.4]
  input   io_enable, // @[:@66645.4]
  output  io_done, // @[:@66645.4]
  output  io_doneLatch, // @[:@66645.4]
  input   io_ctrDone, // @[:@66645.4]
  output  io_datapathEn, // @[:@66645.4]
  output  io_ctrInc, // @[:@66645.4]
  output  io_ctrRst, // @[:@66645.4]
  input   io_parentAck, // @[:@66645.4]
  input   io_backpressure, // @[:@66645.4]
  input   io_break // @[:@66645.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@66647.4]
  wire  active_reset; // @[Controllers.scala 261:22:@66647.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@66647.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@66647.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@66647.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@66647.4]
  wire  done_clock; // @[Controllers.scala 262:20:@66650.4]
  wire  done_reset; // @[Controllers.scala 262:20:@66650.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@66650.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@66650.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@66650.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@66650.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@66684.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@66684.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@66684.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@66684.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@66684.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@66706.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@66706.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@66706.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@66706.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@66706.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@66718.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@66718.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@66718.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@66718.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@66718.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@66726.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@66726.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@66726.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@66726.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@66726.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@66742.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@66742.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@66742.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@66742.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@66742.4]
  wire  _T_80; // @[Controllers.scala 264:48:@66655.4]
  wire  _T_81; // @[Controllers.scala 264:46:@66656.4]
  wire  _T_82; // @[Controllers.scala 264:62:@66657.4]
  wire  _T_83; // @[Controllers.scala 264:60:@66658.4]
  wire  _T_100; // @[package.scala 100:49:@66675.4]
  reg  _T_103; // @[package.scala 48:56:@66676.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@66689.4 package.scala 96:25:@66690.4]
  wire  _T_110; // @[package.scala 100:49:@66691.4]
  reg  _T_113; // @[package.scala 48:56:@66692.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@66694.4]
  wire  _T_118; // @[Controllers.scala 283:41:@66699.4]
  wire  _T_119; // @[Controllers.scala 283:59:@66700.4]
  wire  _T_121; // @[Controllers.scala 284:37:@66703.4]
  wire  _T_124; // @[package.scala 96:25:@66711.4 package.scala 96:25:@66712.4]
  wire  _T_126; // @[package.scala 100:49:@66713.4]
  reg  _T_129; // @[package.scala 48:56:@66714.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@66736.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@66738.4]
  reg  _T_153; // @[package.scala 48:56:@66739.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@66747.4 package.scala 96:25:@66748.4]
  wire  _T_158; // @[Controllers.scala 292:61:@66749.4]
  wire  _T_159; // @[Controllers.scala 292:24:@66750.4]
  SRFF active ( // @[Controllers.scala 261:22:@66647.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@66650.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@66684.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@66706.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@66718.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@66726.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@66742.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@66655.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@66656.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@66657.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@66658.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@66675.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@66689.4 package.scala 96:25:@66690.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@66691.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@66694.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@66699.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@66700.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@66703.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@66711.4 package.scala 96:25:@66712.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@66713.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@66738.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@66747.4 package.scala 96:25:@66748.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@66749.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@66750.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@66717.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@66752.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@66702.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@66705.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@66697.4]
  assign active_clock = clock; // @[:@66648.4]
  assign active_reset = reset; // @[:@66649.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@66660.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@66664.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@66665.4]
  assign done_clock = clock; // @[:@66651.4]
  assign done_reset = reset; // @[:@66652.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@66680.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@66673.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@66674.4]
  assign RetimeWrapper_clock = clock; // @[:@66685.4]
  assign RetimeWrapper_reset = reset; // @[:@66686.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@66688.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@66687.4]
  assign RetimeWrapper_1_clock = clock; // @[:@66707.4]
  assign RetimeWrapper_1_reset = reset; // @[:@66708.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@66710.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@66709.4]
  assign RetimeWrapper_2_clock = clock; // @[:@66719.4]
  assign RetimeWrapper_2_reset = reset; // @[:@66720.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@66722.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@66721.4]
  assign RetimeWrapper_3_clock = clock; // @[:@66727.4]
  assign RetimeWrapper_3_reset = reset; // @[:@66728.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@66730.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@66729.4]
  assign RetimeWrapper_4_clock = clock; // @[:@66743.4]
  assign RetimeWrapper_4_reset = reset; // @[:@66744.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@66746.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@66745.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x688_inr_Foreach_kernelx688_inr_Foreach_concrete1( // @[:@66959.2]
  input         clock, // @[:@66960.4]
  input         reset, // @[:@66961.4]
  output [20:0] io_in_x344_outbuf_0_rPort_0_ofs_0, // @[:@66962.4]
  output        io_in_x344_outbuf_0_rPort_0_en_0, // @[:@66962.4]
  output        io_in_x344_outbuf_0_rPort_0_backpressure, // @[:@66962.4]
  input  [31:0] io_in_x344_outbuf_0_rPort_0_output_0, // @[:@66962.4]
  output        io_in_x673_valid, // @[:@66962.4]
  output [31:0] io_in_x673_bits_wdata_0, // @[:@66962.4]
  output        io_in_x673_bits_wstrb, // @[:@66962.4]
  input         io_sigsIn_backpressure, // @[:@66962.4]
  input         io_sigsIn_datapathEn, // @[:@66962.4]
  input         io_sigsIn_break, // @[:@66962.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@66962.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@66962.4]
  input         io_rr // @[:@66962.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@66989.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@66989.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@67018.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@67018.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@67018.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@67018.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@67018.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@67027.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@67027.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@67027.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@67027.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@67027.4]
  wire  b683; // @[sm_x688_inr_Foreach.scala 62:18:@66997.4]
  wire  _T_274; // @[sm_x688_inr_Foreach.scala 67:129:@67001.4]
  wire  _T_278; // @[implicits.scala 55:10:@67004.4]
  wire  _T_279; // @[sm_x688_inr_Foreach.scala 67:146:@67005.4]
  wire [32:0] x686_tuple; // @[Cat.scala 30:58:@67015.4]
  wire  _T_290; // @[package.scala 96:25:@67032.4 package.scala 96:25:@67033.4]
  wire  _T_292; // @[implicits.scala 55:10:@67034.4]
  wire  x864_b683_D2; // @[package.scala 96:25:@67023.4 package.scala 96:25:@67024.4]
  wire  _T_293; // @[sm_x688_inr_Foreach.scala 74:112:@67035.4]
  wire [31:0] b682_number; // @[Math.scala 723:22:@66994.4 Math.scala 724:14:@66995.4]
  _ _ ( // @[Math.scala 720:24:@66989.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@67018.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@67027.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b683 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x688_inr_Foreach.scala 62:18:@66997.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x688_inr_Foreach.scala 67:129:@67001.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@67004.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x688_inr_Foreach.scala 67:146:@67005.4]
  assign x686_tuple = {1'h1,io_in_x344_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@67015.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@67032.4 package.scala 96:25:@67033.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@67034.4]
  assign x864_b683_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@67023.4 package.scala 96:25:@67024.4]
  assign _T_293 = _T_292 & x864_b683_D2; // @[sm_x688_inr_Foreach.scala 74:112:@67035.4]
  assign b682_number = __io_result; // @[Math.scala 723:22:@66994.4 Math.scala 724:14:@66995.4]
  assign io_in_x344_outbuf_0_rPort_0_ofs_0 = b682_number[20:0]; // @[MemInterfaceType.scala 107:54:@67008.4]
  assign io_in_x344_outbuf_0_rPort_0_en_0 = _T_279 & b683; // @[MemInterfaceType.scala 110:79:@67010.4]
  assign io_in_x344_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@67009.4]
  assign io_in_x673_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x688_inr_Foreach.scala 74:18:@67037.4]
  assign io_in_x673_bits_wdata_0 = x686_tuple[31:0]; // @[sm_x688_inr_Foreach.scala 75:26:@67039.4]
  assign io_in_x673_bits_wstrb = x686_tuple[32]; // @[sm_x688_inr_Foreach.scala 76:23:@67041.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@66992.4]
  assign RetimeWrapper_clock = clock; // @[:@67019.4]
  assign RetimeWrapper_reset = reset; // @[:@67020.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@67022.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@67021.4]
  assign RetimeWrapper_1_clock = clock; // @[:@67028.4]
  assign RetimeWrapper_1_reset = reset; // @[:@67029.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@67031.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@67030.4]
endmodule
module x692_inr_UnitPipe_sm( // @[:@67197.2]
  input   clock, // @[:@67198.4]
  input   reset, // @[:@67199.4]
  input   io_enable, // @[:@67200.4]
  output  io_done, // @[:@67200.4]
  output  io_doneLatch, // @[:@67200.4]
  input   io_ctrDone, // @[:@67200.4]
  output  io_datapathEn, // @[:@67200.4]
  output  io_ctrInc, // @[:@67200.4]
  input   io_parentAck // @[:@67200.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@67202.4]
  wire  active_reset; // @[Controllers.scala 261:22:@67202.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@67202.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@67202.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@67202.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@67202.4]
  wire  done_clock; // @[Controllers.scala 262:20:@67205.4]
  wire  done_reset; // @[Controllers.scala 262:20:@67205.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@67205.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@67205.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@67205.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@67205.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@67239.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@67239.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@67239.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@67239.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@67239.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@67261.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@67261.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@67261.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@67261.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@67261.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@67273.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@67273.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@67273.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@67273.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@67273.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@67281.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@67281.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@67281.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@67281.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@67281.4]
  wire  _T_80; // @[Controllers.scala 264:48:@67210.4]
  wire  _T_81; // @[Controllers.scala 264:46:@67211.4]
  wire  _T_82; // @[Controllers.scala 264:62:@67212.4]
  wire  _T_100; // @[package.scala 100:49:@67230.4]
  reg  _T_103; // @[package.scala 48:56:@67231.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@67254.4]
  wire  _T_124; // @[package.scala 96:25:@67266.4 package.scala 96:25:@67267.4]
  wire  _T_126; // @[package.scala 100:49:@67268.4]
  reg  _T_129; // @[package.scala 48:56:@67269.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@67291.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@67293.4]
  reg  _T_153; // @[package.scala 48:56:@67294.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@67296.4]
  wire  _T_156; // @[Controllers.scala 292:61:@67297.4]
  wire  _T_157; // @[Controllers.scala 292:24:@67298.4]
  SRFF active ( // @[Controllers.scala 261:22:@67202.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@67205.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@67239.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@67261.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@67273.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@67281.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@67210.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@67211.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@67212.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@67230.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@67254.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@67266.4 package.scala 96:25:@67267.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@67268.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@67293.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@67296.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@67297.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@67298.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@67272.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@67300.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@67257.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@67260.4]
  assign active_clock = clock; // @[:@67203.4]
  assign active_reset = reset; // @[:@67204.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@67215.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@67219.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@67220.4]
  assign done_clock = clock; // @[:@67206.4]
  assign done_reset = reset; // @[:@67207.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@67235.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@67228.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@67229.4]
  assign RetimeWrapper_clock = clock; // @[:@67240.4]
  assign RetimeWrapper_reset = reset; // @[:@67241.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@67243.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@67242.4]
  assign RetimeWrapper_1_clock = clock; // @[:@67262.4]
  assign RetimeWrapper_1_reset = reset; // @[:@67263.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@67265.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@67264.4]
  assign RetimeWrapper_2_clock = clock; // @[:@67274.4]
  assign RetimeWrapper_2_reset = reset; // @[:@67275.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@67277.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@67276.4]
  assign RetimeWrapper_3_clock = clock; // @[:@67282.4]
  assign RetimeWrapper_3_reset = reset; // @[:@67283.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@67285.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@67284.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1( // @[:@67375.2]
  output  io_in_x674_ready, // @[:@67378.4]
  input   io_sigsIn_datapathEn // @[:@67378.4]
);
  assign io_in_x674_ready = io_sigsIn_datapathEn; // @[sm_x692_inr_UnitPipe.scala 57:18:@67390.4]
endmodule
module x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1( // @[:@67393.2]
  input         clock, // @[:@67394.4]
  input         reset, // @[:@67395.4]
  input  [63:0] io_in_x340_outdram_number, // @[:@67396.4]
  output [20:0] io_in_x344_outbuf_0_rPort_0_ofs_0, // @[:@67396.4]
  output        io_in_x344_outbuf_0_rPort_0_en_0, // @[:@67396.4]
  output        io_in_x344_outbuf_0_rPort_0_backpressure, // @[:@67396.4]
  input  [31:0] io_in_x344_outbuf_0_rPort_0_output_0, // @[:@67396.4]
  output        io_in_x674_ready, // @[:@67396.4]
  input         io_in_x674_valid, // @[:@67396.4]
  input         io_in_x672_ready, // @[:@67396.4]
  output        io_in_x672_valid, // @[:@67396.4]
  output [63:0] io_in_x672_bits_addr, // @[:@67396.4]
  output [31:0] io_in_x672_bits_size, // @[:@67396.4]
  input         io_in_x673_ready, // @[:@67396.4]
  output        io_in_x673_valid, // @[:@67396.4]
  output [31:0] io_in_x673_bits_wdata_0, // @[:@67396.4]
  output        io_in_x673_bits_wstrb, // @[:@67396.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@67396.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@67396.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@67396.4]
  input         io_sigsIn_smChildAcks_0, // @[:@67396.4]
  input         io_sigsIn_smChildAcks_1, // @[:@67396.4]
  input         io_sigsIn_smChildAcks_2, // @[:@67396.4]
  output        io_sigsOut_smDoneIn_0, // @[:@67396.4]
  output        io_sigsOut_smDoneIn_1, // @[:@67396.4]
  output        io_sigsOut_smDoneIn_2, // @[:@67396.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@67396.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@67396.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@67396.4]
  input         io_rr // @[:@67396.4]
);
  wire  x679_inr_UnitPipe_sm_clock; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_reset; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_io_enable; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_io_done; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_io_doneLatch; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_io_ctrDone; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_io_datapathEn; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_io_ctrInc; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_io_parentAck; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  x679_inr_UnitPipe_sm_io_backpressure; // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@67520.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@67520.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@67520.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@67520.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@67520.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@67528.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@67528.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@67528.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@67528.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@67528.4]
  wire [63:0] x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x340_outdram_number; // @[sm_x679_inr_UnitPipe.scala 69:24:@67558.4]
  wire  x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_valid; // @[sm_x679_inr_UnitPipe.scala 69:24:@67558.4]
  wire [63:0] x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_bits_addr; // @[sm_x679_inr_UnitPipe.scala 69:24:@67558.4]
  wire [31:0] x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_bits_size; // @[sm_x679_inr_UnitPipe.scala 69:24:@67558.4]
  wire  x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x679_inr_UnitPipe.scala 69:24:@67558.4]
  wire  x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x679_inr_UnitPipe.scala 69:24:@67558.4]
  wire  x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_rr; // @[sm_x679_inr_UnitPipe.scala 69:24:@67558.4]
  wire  x681_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@67626.4]
  wire  x681_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@67626.4]
  wire  x681_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@67626.4]
  wire  x681_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@67626.4]
  wire [22:0] x681_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@67626.4]
  wire  x681_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@67626.4]
  wire  x681_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@67626.4]
  wire  x688_inr_Foreach_sm_clock; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_reset; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_enable; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_done; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_doneLatch; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_ctrDone; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_datapathEn; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_ctrInc; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_ctrRst; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_parentAck; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_backpressure; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  x688_inr_Foreach_sm_io_break; // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@67707.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@67707.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@67707.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@67707.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@67707.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@67747.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@67747.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@67747.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@67747.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@67747.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@67755.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@67755.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@67755.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@67755.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@67755.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_clock; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_reset; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire [20:0] x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_en_0; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire [31:0] x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_output_0; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_valid; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire [31:0] x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_bits_wdata_0; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_bits_wstrb; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire [31:0] x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_rr; // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
  wire  x692_inr_UnitPipe_sm_clock; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  x692_inr_UnitPipe_sm_reset; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  x692_inr_UnitPipe_sm_io_enable; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  x692_inr_UnitPipe_sm_io_done; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  x692_inr_UnitPipe_sm_io_doneLatch; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  x692_inr_UnitPipe_sm_io_ctrDone; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  x692_inr_UnitPipe_sm_io_datapathEn; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  x692_inr_UnitPipe_sm_io_ctrInc; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  x692_inr_UnitPipe_sm_io_parentAck; // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@67967.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@67967.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@67967.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@67967.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@67967.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@67975.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@67975.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@67975.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@67975.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@67975.4]
  wire  x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1_io_in_x674_ready; // @[sm_x692_inr_UnitPipe.scala 60:24:@68005.4]
  wire  x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x692_inr_UnitPipe.scala 60:24:@68005.4]
  wire  _T_359; // @[package.scala 100:49:@67491.4]
  reg  _T_362; // @[package.scala 48:56:@67492.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@67525.4 package.scala 96:25:@67526.4]
  wire  _T_381; // @[package.scala 96:25:@67533.4 package.scala 96:25:@67534.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@67536.4]
  wire  _T_454; // @[package.scala 96:25:@67712.4 package.scala 96:25:@67713.4]
  wire  _T_468; // @[package.scala 96:25:@67752.4 package.scala 96:25:@67753.4]
  wire  _T_474; // @[package.scala 96:25:@67760.4 package.scala 96:25:@67761.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@67763.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@67772.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@67773.4]
  wire  _T_547; // @[package.scala 100:49:@67938.4]
  reg  _T_550; // @[package.scala 48:56:@67939.4]
  reg [31:0] _RAND_1;
  wire  x692_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x693_outr_UnitPipe.scala 101:55:@67945.4]
  wire  _T_563; // @[package.scala 96:25:@67972.4 package.scala 96:25:@67973.4]
  wire  _T_569; // @[package.scala 96:25:@67980.4 package.scala 96:25:@67981.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@67983.4]
  wire  x692_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@67984.4]
  x679_inr_UnitPipe_sm x679_inr_UnitPipe_sm ( // @[sm_x679_inr_UnitPipe.scala 33:18:@67463.4]
    .clock(x679_inr_UnitPipe_sm_clock),
    .reset(x679_inr_UnitPipe_sm_reset),
    .io_enable(x679_inr_UnitPipe_sm_io_enable),
    .io_done(x679_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x679_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x679_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x679_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x679_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x679_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x679_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@67520.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@67528.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1 x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1 ( // @[sm_x679_inr_UnitPipe.scala 69:24:@67558.4]
    .io_in_x340_outdram_number(x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x340_outdram_number),
    .io_in_x672_valid(x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_valid),
    .io_in_x672_bits_addr(x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_bits_addr),
    .io_in_x672_bits_size(x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_bits_size),
    .io_sigsIn_backpressure(x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_rr)
  );
  x681_ctrchain x681_ctrchain ( // @[SpatialBlocks.scala 37:22:@67626.4]
    .clock(x681_ctrchain_clock),
    .reset(x681_ctrchain_reset),
    .io_input_reset(x681_ctrchain_io_input_reset),
    .io_input_enable(x681_ctrchain_io_input_enable),
    .io_output_counts_0(x681_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x681_ctrchain_io_output_oobs_0),
    .io_output_done(x681_ctrchain_io_output_done)
  );
  x688_inr_Foreach_sm x688_inr_Foreach_sm ( // @[sm_x688_inr_Foreach.scala 33:18:@67679.4]
    .clock(x688_inr_Foreach_sm_clock),
    .reset(x688_inr_Foreach_sm_reset),
    .io_enable(x688_inr_Foreach_sm_io_enable),
    .io_done(x688_inr_Foreach_sm_io_done),
    .io_doneLatch(x688_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x688_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x688_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x688_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x688_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x688_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x688_inr_Foreach_sm_io_backpressure),
    .io_break(x688_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@67707.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@67747.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@67755.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x688_inr_Foreach_kernelx688_inr_Foreach_concrete1 x688_inr_Foreach_kernelx688_inr_Foreach_concrete1 ( // @[sm_x688_inr_Foreach.scala 78:24:@67790.4]
    .clock(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_clock),
    .reset(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_reset),
    .io_in_x344_outbuf_0_rPort_0_ofs_0(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0),
    .io_in_x344_outbuf_0_rPort_0_en_0(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_en_0),
    .io_in_x344_outbuf_0_rPort_0_backpressure(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure),
    .io_in_x344_outbuf_0_rPort_0_output_0(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_output_0),
    .io_in_x673_valid(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_valid),
    .io_in_x673_bits_wdata_0(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_bits_wdata_0),
    .io_in_x673_bits_wstrb(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_bits_wstrb),
    .io_sigsIn_backpressure(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_rr)
  );
  x692_inr_UnitPipe_sm x692_inr_UnitPipe_sm ( // @[sm_x692_inr_UnitPipe.scala 32:18:@67910.4]
    .clock(x692_inr_UnitPipe_sm_clock),
    .reset(x692_inr_UnitPipe_sm_reset),
    .io_enable(x692_inr_UnitPipe_sm_io_enable),
    .io_done(x692_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x692_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x692_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x692_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x692_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x692_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@67967.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@67975.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1 x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1 ( // @[sm_x692_inr_UnitPipe.scala 60:24:@68005.4]
    .io_in_x674_ready(x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1_io_in_x674_ready),
    .io_sigsIn_datapathEn(x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x679_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@67491.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@67525.4 package.scala 96:25:@67526.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@67533.4 package.scala 96:25:@67534.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@67536.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@67712.4 package.scala 96:25:@67713.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@67752.4 package.scala 96:25:@67753.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@67760.4 package.scala 96:25:@67761.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@67763.4]
  assign _T_479 = x688_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@67772.4]
  assign _T_480 = ~ x688_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@67773.4]
  assign _T_547 = x692_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@67938.4]
  assign x692_inr_UnitPipe_sigsIn_forwardpressure = io_in_x674_valid | x692_inr_UnitPipe_sm_io_doneLatch; // @[sm_x693_outr_UnitPipe.scala 101:55:@67945.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@67972.4 package.scala 96:25:@67973.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@67980.4 package.scala 96:25:@67981.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@67983.4]
  assign x692_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@67984.4]
  assign io_in_x344_outbuf_0_rPort_0_ofs_0 = x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@67841.4]
  assign io_in_x344_outbuf_0_rPort_0_en_0 = x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@67840.4]
  assign io_in_x344_outbuf_0_rPort_0_backpressure = x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@67839.4]
  assign io_in_x674_ready = x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1_io_in_x674_ready; // @[sm_x692_inr_UnitPipe.scala 46:23:@68041.4]
  assign io_in_x672_valid = x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_valid; // @[sm_x679_inr_UnitPipe.scala 50:23:@67597.4]
  assign io_in_x672_bits_addr = x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_bits_addr; // @[sm_x679_inr_UnitPipe.scala 50:23:@67596.4]
  assign io_in_x672_bits_size = x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x672_bits_size; // @[sm_x679_inr_UnitPipe.scala 50:23:@67595.4]
  assign io_in_x673_valid = x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_valid; // @[sm_x688_inr_Foreach.scala 50:23:@67845.4]
  assign io_in_x673_bits_wdata_0 = x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_bits_wdata_0; // @[sm_x688_inr_Foreach.scala 50:23:@67844.4]
  assign io_in_x673_bits_wstrb = x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x673_bits_wstrb; // @[sm_x688_inr_Foreach.scala 50:23:@67843.4]
  assign io_sigsOut_smDoneIn_0 = x679_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@67543.4]
  assign io_sigsOut_smDoneIn_1 = x688_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@67770.4]
  assign io_sigsOut_smDoneIn_2 = x692_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@67990.4]
  assign io_sigsOut_smCtrCopyDone_0 = x679_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@67557.4]
  assign io_sigsOut_smCtrCopyDone_1 = x688_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@67789.4]
  assign io_sigsOut_smCtrCopyDone_2 = x692_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@68004.4]
  assign x679_inr_UnitPipe_sm_clock = clock; // @[:@67464.4]
  assign x679_inr_UnitPipe_sm_reset = reset; // @[:@67465.4]
  assign x679_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@67540.4]
  assign x679_inr_UnitPipe_sm_io_ctrDone = x679_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x693_outr_UnitPipe.scala 77:39:@67495.4]
  assign x679_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@67542.4]
  assign x679_inr_UnitPipe_sm_io_backpressure = io_in_x672_ready | x679_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@67514.4]
  assign RetimeWrapper_clock = clock; // @[:@67521.4]
  assign RetimeWrapper_reset = reset; // @[:@67522.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@67524.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@67523.4]
  assign RetimeWrapper_1_clock = clock; // @[:@67529.4]
  assign RetimeWrapper_1_reset = reset; // @[:@67530.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@67532.4]
  assign RetimeWrapper_1_io_in = x679_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@67531.4]
  assign x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_in_x340_outdram_number = io_in_x340_outdram_number; // @[sm_x679_inr_UnitPipe.scala 49:31:@67594.4]
  assign x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x672_ready | x679_inr_UnitPipe_sm_io_doneLatch; // @[sm_x679_inr_UnitPipe.scala 74:22:@67613.4]
  assign x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x679_inr_UnitPipe_sm_io_datapathEn; // @[sm_x679_inr_UnitPipe.scala 74:22:@67611.4]
  assign x679_inr_UnitPipe_kernelx679_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x679_inr_UnitPipe.scala 73:18:@67599.4]
  assign x681_ctrchain_clock = clock; // @[:@67627.4]
  assign x681_ctrchain_reset = reset; // @[:@67628.4]
  assign x681_ctrchain_io_input_reset = x688_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@67788.4]
  assign x681_ctrchain_io_input_enable = x688_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@67740.4 SpatialBlocks.scala 159:42:@67787.4]
  assign x688_inr_Foreach_sm_clock = clock; // @[:@67680.4]
  assign x688_inr_Foreach_sm_reset = reset; // @[:@67681.4]
  assign x688_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@67767.4]
  assign x688_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x693_outr_UnitPipe.scala 90:38:@67715.4]
  assign x688_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@67769.4]
  assign x688_inr_Foreach_sm_io_backpressure = io_in_x673_ready | x688_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@67741.4]
  assign x688_inr_Foreach_sm_io_break = 1'h0; // @[sm_x693_outr_UnitPipe.scala 94:36:@67721.4]
  assign RetimeWrapper_2_clock = clock; // @[:@67708.4]
  assign RetimeWrapper_2_reset = reset; // @[:@67709.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@67711.4]
  assign RetimeWrapper_2_io_in = x681_ctrchain_io_output_done; // @[package.scala 94:16:@67710.4]
  assign RetimeWrapper_3_clock = clock; // @[:@67748.4]
  assign RetimeWrapper_3_reset = reset; // @[:@67749.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@67751.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@67750.4]
  assign RetimeWrapper_4_clock = clock; // @[:@67756.4]
  assign RetimeWrapper_4_reset = reset; // @[:@67757.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@67759.4]
  assign RetimeWrapper_4_io_in = x688_inr_Foreach_sm_io_done; // @[package.scala 94:16:@67758.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_clock = clock; // @[:@67791.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_reset = reset; // @[:@67792.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_in_x344_outbuf_0_rPort_0_output_0 = io_in_x344_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@67838.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x673_ready | x688_inr_Foreach_sm_io_doneLatch; // @[sm_x688_inr_Foreach.scala 83:22:@67861.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x688_inr_Foreach.scala 83:22:@67859.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_break = x688_inr_Foreach_sm_io_break; // @[sm_x688_inr_Foreach.scala 83:22:@67857.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x681_ctrchain_io_output_counts_0[22]}},x681_ctrchain_io_output_counts_0}; // @[sm_x688_inr_Foreach.scala 83:22:@67852.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x681_ctrchain_io_output_oobs_0; // @[sm_x688_inr_Foreach.scala 83:22:@67851.4]
  assign x688_inr_Foreach_kernelx688_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x688_inr_Foreach.scala 82:18:@67847.4]
  assign x692_inr_UnitPipe_sm_clock = clock; // @[:@67911.4]
  assign x692_inr_UnitPipe_sm_reset = reset; // @[:@67912.4]
  assign x692_inr_UnitPipe_sm_io_enable = x692_inr_UnitPipe_sigsIn_baseEn & x692_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@67987.4]
  assign x692_inr_UnitPipe_sm_io_ctrDone = x692_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x693_outr_UnitPipe.scala 99:39:@67942.4]
  assign x692_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@67989.4]
  assign RetimeWrapper_5_clock = clock; // @[:@67968.4]
  assign RetimeWrapper_5_reset = reset; // @[:@67969.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@67971.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@67970.4]
  assign RetimeWrapper_6_clock = clock; // @[:@67976.4]
  assign RetimeWrapper_6_reset = reset; // @[:@67977.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@67979.4]
  assign RetimeWrapper_6_io_in = x692_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@67978.4]
  assign x692_inr_UnitPipe_kernelx692_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x692_inr_UnitPipe_sm_io_datapathEn; // @[sm_x692_inr_UnitPipe.scala 65:22:@68054.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x740_kernelx740_concrete1( // @[:@68070.2]
  input          clock, // @[:@68071.4]
  input          reset, // @[:@68072.4]
  input  [63:0]  io_in_x340_outdram_number, // @[:@68073.4]
  output [20:0]  io_in_x344_outbuf_0_rPort_0_ofs_0, // @[:@68073.4]
  output         io_in_x344_outbuf_0_rPort_0_en_0, // @[:@68073.4]
  output         io_in_x344_outbuf_0_rPort_0_backpressure, // @[:@68073.4]
  input  [31:0]  io_in_x344_outbuf_0_rPort_0_output_0, // @[:@68073.4]
  output         io_in_x343_TVALID, // @[:@68073.4]
  input          io_in_x343_TREADY, // @[:@68073.4]
  output [255:0] io_in_x343_TDATA, // @[:@68073.4]
  output         io_in_x674_ready, // @[:@68073.4]
  input          io_in_x674_valid, // @[:@68073.4]
  input          io_in_x672_ready, // @[:@68073.4]
  output         io_in_x672_valid, // @[:@68073.4]
  output [63:0]  io_in_x672_bits_addr, // @[:@68073.4]
  output [31:0]  io_in_x672_bits_size, // @[:@68073.4]
  input          io_in_x342_TVALID, // @[:@68073.4]
  output         io_in_x342_TREADY, // @[:@68073.4]
  input  [255:0] io_in_x342_TDATA, // @[:@68073.4]
  input  [7:0]   io_in_x342_TID, // @[:@68073.4]
  input  [7:0]   io_in_x342_TDEST, // @[:@68073.4]
  input          io_in_x673_ready, // @[:@68073.4]
  output         io_in_x673_valid, // @[:@68073.4]
  output [31:0]  io_in_x673_bits_wdata_0, // @[:@68073.4]
  output         io_in_x673_bits_wstrb, // @[:@68073.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@68073.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@68073.4]
  input          io_sigsIn_smChildAcks_0, // @[:@68073.4]
  input          io_sigsIn_smChildAcks_1, // @[:@68073.4]
  output         io_sigsOut_smDoneIn_0, // @[:@68073.4]
  output         io_sigsOut_smDoneIn_1, // @[:@68073.4]
  input          io_rr // @[:@68073.4]
);
  wire  x671_outr_UnitPipe_sm_clock; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_reset; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_enable; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_done; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_parentAck; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_childAck_0; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_childAck_1; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  x671_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@68208.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@68208.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@68208.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@68208.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@68208.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@68216.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@68216.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_clock; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_reset; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TVALID; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TREADY; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire [255:0] x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TDATA; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TVALID; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TREADY; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire [255:0] x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TDATA; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire [7:0] x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TID; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire [7:0] x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TDEST; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_rr; // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
  wire  x693_outr_UnitPipe_sm_clock; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_reset; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_enable; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_done; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_parentAck; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_childAck_0; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_childAck_1; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_childAck_2; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  x693_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@68497.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@68497.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@68497.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@68497.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@68497.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@68505.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@68505.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@68505.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@68505.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@68505.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_clock; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_reset; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire [63:0] x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x340_outdram_number; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire [20:0] x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_en_0; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire [31:0] x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_output_0; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x674_ready; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x674_valid; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_ready; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_valid; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire [63:0] x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_bits_addr; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire [31:0] x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_bits_size; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_ready; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_valid; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire [31:0] x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_bits_wdata_0; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_bits_wstrb; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_rr; // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
  wire  _T_408; // @[package.scala 96:25:@68213.4 package.scala 96:25:@68214.4]
  wire  _T_414; // @[package.scala 96:25:@68221.4 package.scala 96:25:@68222.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@68224.4]
  wire  _T_508; // @[package.scala 96:25:@68502.4 package.scala 96:25:@68503.4]
  wire  _T_514; // @[package.scala 96:25:@68510.4 package.scala 96:25:@68511.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@68513.4]
  x671_outr_UnitPipe_sm x671_outr_UnitPipe_sm ( // @[sm_x671_outr_UnitPipe.scala 32:18:@68146.4]
    .clock(x671_outr_UnitPipe_sm_clock),
    .reset(x671_outr_UnitPipe_sm_reset),
    .io_enable(x671_outr_UnitPipe_sm_io_enable),
    .io_done(x671_outr_UnitPipe_sm_io_done),
    .io_parentAck(x671_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x671_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x671_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x671_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x671_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x671_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x671_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x671_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x671_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@68208.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@68216.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1 x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1 ( // @[sm_x671_outr_UnitPipe.scala 87:24:@68247.4]
    .clock(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_clock),
    .reset(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_reset),
    .io_in_x343_TVALID(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TVALID),
    .io_in_x343_TREADY(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TREADY),
    .io_in_x343_TDATA(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TDATA),
    .io_in_x342_TVALID(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TVALID),
    .io_in_x342_TREADY(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TREADY),
    .io_in_x342_TDATA(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TDATA),
    .io_in_x342_TID(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TID),
    .io_in_x342_TDEST(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TDEST),
    .io_sigsIn_smEnableOuts_0(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_rr)
  );
  x693_outr_UnitPipe_sm x693_outr_UnitPipe_sm ( // @[sm_x693_outr_UnitPipe.scala 36:18:@68425.4]
    .clock(x693_outr_UnitPipe_sm_clock),
    .reset(x693_outr_UnitPipe_sm_reset),
    .io_enable(x693_outr_UnitPipe_sm_io_enable),
    .io_done(x693_outr_UnitPipe_sm_io_done),
    .io_parentAck(x693_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x693_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x693_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x693_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x693_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x693_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x693_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x693_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x693_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x693_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x693_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x693_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x693_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@68497.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@68505.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1 x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1 ( // @[sm_x693_outr_UnitPipe.scala 108:24:@68537.4]
    .clock(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_clock),
    .reset(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_reset),
    .io_in_x340_outdram_number(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x340_outdram_number),
    .io_in_x344_outbuf_0_rPort_0_ofs_0(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0),
    .io_in_x344_outbuf_0_rPort_0_en_0(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_en_0),
    .io_in_x344_outbuf_0_rPort_0_backpressure(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure),
    .io_in_x344_outbuf_0_rPort_0_output_0(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_output_0),
    .io_in_x674_ready(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x674_ready),
    .io_in_x674_valid(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x674_valid),
    .io_in_x672_ready(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_ready),
    .io_in_x672_valid(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_valid),
    .io_in_x672_bits_addr(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_bits_addr),
    .io_in_x672_bits_size(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_bits_size),
    .io_in_x673_ready(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_ready),
    .io_in_x673_valid(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_valid),
    .io_in_x673_bits_wdata_0(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_bits_wdata_0),
    .io_in_x673_bits_wstrb(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@68213.4 package.scala 96:25:@68214.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@68221.4 package.scala 96:25:@68222.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@68224.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@68502.4 package.scala 96:25:@68503.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@68510.4 package.scala 96:25:@68511.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@68513.4]
  assign io_in_x344_outbuf_0_rPort_0_ofs_0 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@68621.4]
  assign io_in_x344_outbuf_0_rPort_0_en_0 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@68620.4]
  assign io_in_x344_outbuf_0_rPort_0_backpressure = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@68619.4]
  assign io_in_x343_TVALID = x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TVALID; // @[sm_x671_outr_UnitPipe.scala 48:23:@68316.4]
  assign io_in_x343_TDATA = x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TDATA; // @[sm_x671_outr_UnitPipe.scala 48:23:@68314.4]
  assign io_in_x674_ready = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x674_ready; // @[sm_x693_outr_UnitPipe.scala 60:23:@68625.4]
  assign io_in_x672_valid = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_valid; // @[sm_x693_outr_UnitPipe.scala 61:23:@68628.4]
  assign io_in_x672_bits_addr = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_bits_addr; // @[sm_x693_outr_UnitPipe.scala 61:23:@68627.4]
  assign io_in_x672_bits_size = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_bits_size; // @[sm_x693_outr_UnitPipe.scala 61:23:@68626.4]
  assign io_in_x342_TREADY = x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TREADY; // @[sm_x671_outr_UnitPipe.scala 49:23:@68324.4]
  assign io_in_x673_valid = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_valid; // @[sm_x693_outr_UnitPipe.scala 62:23:@68632.4]
  assign io_in_x673_bits_wdata_0 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_bits_wdata_0; // @[sm_x693_outr_UnitPipe.scala 62:23:@68631.4]
  assign io_in_x673_bits_wstrb = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_bits_wstrb; // @[sm_x693_outr_UnitPipe.scala 62:23:@68630.4]
  assign io_sigsOut_smDoneIn_0 = x671_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@68231.4]
  assign io_sigsOut_smDoneIn_1 = x693_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@68520.4]
  assign x671_outr_UnitPipe_sm_clock = clock; // @[:@68147.4]
  assign x671_outr_UnitPipe_sm_reset = reset; // @[:@68148.4]
  assign x671_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@68228.4]
  assign x671_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@68230.4]
  assign x671_outr_UnitPipe_sm_io_doneIn_0 = x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@68198.4]
  assign x671_outr_UnitPipe_sm_io_doneIn_1 = x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@68199.4]
  assign x671_outr_UnitPipe_sm_io_ctrCopyDone_0 = x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@68245.4]
  assign x671_outr_UnitPipe_sm_io_ctrCopyDone_1 = x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@68246.4]
  assign RetimeWrapper_clock = clock; // @[:@68209.4]
  assign RetimeWrapper_reset = reset; // @[:@68210.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@68212.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@68211.4]
  assign RetimeWrapper_1_clock = clock; // @[:@68217.4]
  assign RetimeWrapper_1_reset = reset; // @[:@68218.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@68220.4]
  assign RetimeWrapper_1_io_in = x671_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@68219.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_clock = clock; // @[:@68248.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_reset = reset; // @[:@68249.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x343_TREADY = io_in_x343_TREADY; // @[sm_x671_outr_UnitPipe.scala 48:23:@68315.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TVALID = io_in_x342_TVALID; // @[sm_x671_outr_UnitPipe.scala 49:23:@68325.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TDATA = io_in_x342_TDATA; // @[sm_x671_outr_UnitPipe.scala 49:23:@68323.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TID = io_in_x342_TID; // @[sm_x671_outr_UnitPipe.scala 49:23:@68319.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_in_x342_TDEST = io_in_x342_TDEST; // @[sm_x671_outr_UnitPipe.scala 49:23:@68318.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x671_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x671_outr_UnitPipe.scala 92:22:@68341.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x671_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x671_outr_UnitPipe.scala 92:22:@68342.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x671_outr_UnitPipe_sm_io_childAck_0; // @[sm_x671_outr_UnitPipe.scala 92:22:@68337.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x671_outr_UnitPipe_sm_io_childAck_1; // @[sm_x671_outr_UnitPipe.scala 92:22:@68338.4]
  assign x671_outr_UnitPipe_kernelx671_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x671_outr_UnitPipe.scala 91:18:@68326.4]
  assign x693_outr_UnitPipe_sm_clock = clock; // @[:@68426.4]
  assign x693_outr_UnitPipe_sm_reset = reset; // @[:@68427.4]
  assign x693_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@68517.4]
  assign x693_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@68519.4]
  assign x693_outr_UnitPipe_sm_io_doneIn_0 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@68485.4]
  assign x693_outr_UnitPipe_sm_io_doneIn_1 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@68486.4]
  assign x693_outr_UnitPipe_sm_io_doneIn_2 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@68487.4]
  assign x693_outr_UnitPipe_sm_io_ctrCopyDone_0 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@68534.4]
  assign x693_outr_UnitPipe_sm_io_ctrCopyDone_1 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@68535.4]
  assign x693_outr_UnitPipe_sm_io_ctrCopyDone_2 = x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@68536.4]
  assign RetimeWrapper_2_clock = clock; // @[:@68498.4]
  assign RetimeWrapper_2_reset = reset; // @[:@68499.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@68501.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@68500.4]
  assign RetimeWrapper_3_clock = clock; // @[:@68506.4]
  assign RetimeWrapper_3_reset = reset; // @[:@68507.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@68509.4]
  assign RetimeWrapper_3_io_in = x693_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@68508.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_clock = clock; // @[:@68538.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_reset = reset; // @[:@68539.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x340_outdram_number = io_in_x340_outdram_number; // @[sm_x693_outr_UnitPipe.scala 58:31:@68617.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x344_outbuf_0_rPort_0_output_0 = io_in_x344_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@68618.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x674_valid = io_in_x674_valid; // @[sm_x693_outr_UnitPipe.scala 60:23:@68624.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x672_ready = io_in_x672_ready; // @[sm_x693_outr_UnitPipe.scala 61:23:@68629.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_in_x673_ready = io_in_x673_ready; // @[sm_x693_outr_UnitPipe.scala 62:23:@68633.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x693_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x693_outr_UnitPipe.scala 113:22:@68656.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x693_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x693_outr_UnitPipe.scala 113:22:@68657.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x693_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x693_outr_UnitPipe.scala 113:22:@68658.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x693_outr_UnitPipe_sm_io_childAck_0; // @[sm_x693_outr_UnitPipe.scala 113:22:@68650.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x693_outr_UnitPipe_sm_io_childAck_1; // @[sm_x693_outr_UnitPipe.scala 113:22:@68651.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x693_outr_UnitPipe_sm_io_childAck_2; // @[sm_x693_outr_UnitPipe.scala 113:22:@68652.4]
  assign x693_outr_UnitPipe_kernelx693_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x693_outr_UnitPipe.scala 112:18:@68634.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@68686.2]
  input          clock, // @[:@68687.4]
  input          reset, // @[:@68688.4]
  input  [63:0]  io_in_x340_outdram_number, // @[:@68689.4]
  output         io_in_x343_TVALID, // @[:@68689.4]
  input          io_in_x343_TREADY, // @[:@68689.4]
  output [255:0] io_in_x343_TDATA, // @[:@68689.4]
  output         io_in_x674_ready, // @[:@68689.4]
  input          io_in_x674_valid, // @[:@68689.4]
  input          io_in_x672_ready, // @[:@68689.4]
  output         io_in_x672_valid, // @[:@68689.4]
  output [63:0]  io_in_x672_bits_addr, // @[:@68689.4]
  output [31:0]  io_in_x672_bits_size, // @[:@68689.4]
  input          io_in_x342_TVALID, // @[:@68689.4]
  output         io_in_x342_TREADY, // @[:@68689.4]
  input  [255:0] io_in_x342_TDATA, // @[:@68689.4]
  input  [7:0]   io_in_x342_TID, // @[:@68689.4]
  input  [7:0]   io_in_x342_TDEST, // @[:@68689.4]
  input          io_in_x673_ready, // @[:@68689.4]
  output         io_in_x673_valid, // @[:@68689.4]
  output [31:0]  io_in_x673_bits_wdata_0, // @[:@68689.4]
  output         io_in_x673_bits_wstrb, // @[:@68689.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@68689.4]
  input          io_sigsIn_smChildAcks_0, // @[:@68689.4]
  output         io_sigsOut_smDoneIn_0, // @[:@68689.4]
  input          io_rr // @[:@68689.4]
);
  wire  x344_outbuf_0_clock; // @[m_x344_outbuf_0.scala 27:17:@68699.4]
  wire  x344_outbuf_0_reset; // @[m_x344_outbuf_0.scala 27:17:@68699.4]
  wire [20:0] x344_outbuf_0_io_rPort_0_ofs_0; // @[m_x344_outbuf_0.scala 27:17:@68699.4]
  wire  x344_outbuf_0_io_rPort_0_en_0; // @[m_x344_outbuf_0.scala 27:17:@68699.4]
  wire  x344_outbuf_0_io_rPort_0_backpressure; // @[m_x344_outbuf_0.scala 27:17:@68699.4]
  wire [31:0] x344_outbuf_0_io_rPort_0_output_0; // @[m_x344_outbuf_0.scala 27:17:@68699.4]
  wire  x740_sm_clock; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_reset; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_enable; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_done; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_ctrDone; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_ctrInc; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_parentAck; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_doneIn_0; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_doneIn_1; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_enableOut_0; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_enableOut_1; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_childAck_0; // @[sm_x740.scala 37:18:@68757.4]
  wire  x740_sm_io_childAck_1; // @[sm_x740.scala 37:18:@68757.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@68824.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@68824.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@68824.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@68824.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@68824.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@68832.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@68832.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@68832.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@68832.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@68832.4]
  wire  x740_kernelx740_concrete1_clock; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_reset; // @[sm_x740.scala 102:24:@68861.4]
  wire [63:0] x740_kernelx740_concrete1_io_in_x340_outdram_number; // @[sm_x740.scala 102:24:@68861.4]
  wire [20:0] x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_en_0; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure; // @[sm_x740.scala 102:24:@68861.4]
  wire [31:0] x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_output_0; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x343_TVALID; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x343_TREADY; // @[sm_x740.scala 102:24:@68861.4]
  wire [255:0] x740_kernelx740_concrete1_io_in_x343_TDATA; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x674_ready; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x674_valid; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x672_ready; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x672_valid; // @[sm_x740.scala 102:24:@68861.4]
  wire [63:0] x740_kernelx740_concrete1_io_in_x672_bits_addr; // @[sm_x740.scala 102:24:@68861.4]
  wire [31:0] x740_kernelx740_concrete1_io_in_x672_bits_size; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x342_TVALID; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x342_TREADY; // @[sm_x740.scala 102:24:@68861.4]
  wire [255:0] x740_kernelx740_concrete1_io_in_x342_TDATA; // @[sm_x740.scala 102:24:@68861.4]
  wire [7:0] x740_kernelx740_concrete1_io_in_x342_TID; // @[sm_x740.scala 102:24:@68861.4]
  wire [7:0] x740_kernelx740_concrete1_io_in_x342_TDEST; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x673_ready; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x673_valid; // @[sm_x740.scala 102:24:@68861.4]
  wire [31:0] x740_kernelx740_concrete1_io_in_x673_bits_wdata_0; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_in_x673_bits_wstrb; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x740.scala 102:24:@68861.4]
  wire  x740_kernelx740_concrete1_io_rr; // @[sm_x740.scala 102:24:@68861.4]
  wire  _T_266; // @[package.scala 100:49:@68790.4]
  reg  _T_269; // @[package.scala 48:56:@68791.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@68829.4 package.scala 96:25:@68830.4]
  wire  _T_289; // @[package.scala 96:25:@68837.4 package.scala 96:25:@68838.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@68840.4]
  x344_outbuf_0 x344_outbuf_0 ( // @[m_x344_outbuf_0.scala 27:17:@68699.4]
    .clock(x344_outbuf_0_clock),
    .reset(x344_outbuf_0_reset),
    .io_rPort_0_ofs_0(x344_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x344_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x344_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x344_outbuf_0_io_rPort_0_output_0)
  );
  x740_sm x740_sm ( // @[sm_x740.scala 37:18:@68757.4]
    .clock(x740_sm_clock),
    .reset(x740_sm_reset),
    .io_enable(x740_sm_io_enable),
    .io_done(x740_sm_io_done),
    .io_ctrDone(x740_sm_io_ctrDone),
    .io_ctrInc(x740_sm_io_ctrInc),
    .io_parentAck(x740_sm_io_parentAck),
    .io_doneIn_0(x740_sm_io_doneIn_0),
    .io_doneIn_1(x740_sm_io_doneIn_1),
    .io_enableOut_0(x740_sm_io_enableOut_0),
    .io_enableOut_1(x740_sm_io_enableOut_1),
    .io_childAck_0(x740_sm_io_childAck_0),
    .io_childAck_1(x740_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@68824.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@68832.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x740_kernelx740_concrete1 x740_kernelx740_concrete1 ( // @[sm_x740.scala 102:24:@68861.4]
    .clock(x740_kernelx740_concrete1_clock),
    .reset(x740_kernelx740_concrete1_reset),
    .io_in_x340_outdram_number(x740_kernelx740_concrete1_io_in_x340_outdram_number),
    .io_in_x344_outbuf_0_rPort_0_ofs_0(x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0),
    .io_in_x344_outbuf_0_rPort_0_en_0(x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_en_0),
    .io_in_x344_outbuf_0_rPort_0_backpressure(x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure),
    .io_in_x344_outbuf_0_rPort_0_output_0(x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_output_0),
    .io_in_x343_TVALID(x740_kernelx740_concrete1_io_in_x343_TVALID),
    .io_in_x343_TREADY(x740_kernelx740_concrete1_io_in_x343_TREADY),
    .io_in_x343_TDATA(x740_kernelx740_concrete1_io_in_x343_TDATA),
    .io_in_x674_ready(x740_kernelx740_concrete1_io_in_x674_ready),
    .io_in_x674_valid(x740_kernelx740_concrete1_io_in_x674_valid),
    .io_in_x672_ready(x740_kernelx740_concrete1_io_in_x672_ready),
    .io_in_x672_valid(x740_kernelx740_concrete1_io_in_x672_valid),
    .io_in_x672_bits_addr(x740_kernelx740_concrete1_io_in_x672_bits_addr),
    .io_in_x672_bits_size(x740_kernelx740_concrete1_io_in_x672_bits_size),
    .io_in_x342_TVALID(x740_kernelx740_concrete1_io_in_x342_TVALID),
    .io_in_x342_TREADY(x740_kernelx740_concrete1_io_in_x342_TREADY),
    .io_in_x342_TDATA(x740_kernelx740_concrete1_io_in_x342_TDATA),
    .io_in_x342_TID(x740_kernelx740_concrete1_io_in_x342_TID),
    .io_in_x342_TDEST(x740_kernelx740_concrete1_io_in_x342_TDEST),
    .io_in_x673_ready(x740_kernelx740_concrete1_io_in_x673_ready),
    .io_in_x673_valid(x740_kernelx740_concrete1_io_in_x673_valid),
    .io_in_x673_bits_wdata_0(x740_kernelx740_concrete1_io_in_x673_bits_wdata_0),
    .io_in_x673_bits_wstrb(x740_kernelx740_concrete1_io_in_x673_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(x740_kernelx740_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x740_kernelx740_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x740_kernelx740_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x740_kernelx740_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x740_kernelx740_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x740_kernelx740_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x740_kernelx740_concrete1_io_rr)
  );
  assign _T_266 = x740_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@68790.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@68829.4 package.scala 96:25:@68830.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@68837.4 package.scala 96:25:@68838.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@68840.4]
  assign io_in_x343_TVALID = x740_kernelx740_concrete1_io_in_x343_TVALID; // @[sm_x740.scala 65:23:@68954.4]
  assign io_in_x343_TDATA = x740_kernelx740_concrete1_io_in_x343_TDATA; // @[sm_x740.scala 65:23:@68952.4]
  assign io_in_x674_ready = x740_kernelx740_concrete1_io_in_x674_ready; // @[sm_x740.scala 66:23:@68957.4]
  assign io_in_x672_valid = x740_kernelx740_concrete1_io_in_x672_valid; // @[sm_x740.scala 67:23:@68960.4]
  assign io_in_x672_bits_addr = x740_kernelx740_concrete1_io_in_x672_bits_addr; // @[sm_x740.scala 67:23:@68959.4]
  assign io_in_x672_bits_size = x740_kernelx740_concrete1_io_in_x672_bits_size; // @[sm_x740.scala 67:23:@68958.4]
  assign io_in_x342_TREADY = x740_kernelx740_concrete1_io_in_x342_TREADY; // @[sm_x740.scala 68:23:@68969.4]
  assign io_in_x673_valid = x740_kernelx740_concrete1_io_in_x673_valid; // @[sm_x740.scala 69:23:@68973.4]
  assign io_in_x673_bits_wdata_0 = x740_kernelx740_concrete1_io_in_x673_bits_wdata_0; // @[sm_x740.scala 69:23:@68972.4]
  assign io_in_x673_bits_wstrb = x740_kernelx740_concrete1_io_in_x673_bits_wstrb; // @[sm_x740.scala 69:23:@68971.4]
  assign io_sigsOut_smDoneIn_0 = x740_sm_io_done; // @[SpatialBlocks.scala 156:53:@68847.4]
  assign x344_outbuf_0_clock = clock; // @[:@68700.4]
  assign x344_outbuf_0_reset = reset; // @[:@68701.4]
  assign x344_outbuf_0_io_rPort_0_ofs_0 = x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@68944.4]
  assign x344_outbuf_0_io_rPort_0_en_0 = x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@68943.4]
  assign x344_outbuf_0_io_rPort_0_backpressure = x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@68942.4]
  assign x740_sm_clock = clock; // @[:@68758.4]
  assign x740_sm_reset = reset; // @[:@68759.4]
  assign x740_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@68844.4]
  assign x740_sm_io_ctrDone = x740_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@68794.4]
  assign x740_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@68846.4]
  assign x740_sm_io_doneIn_0 = x740_kernelx740_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@68814.4]
  assign x740_sm_io_doneIn_1 = x740_kernelx740_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@68815.4]
  assign RetimeWrapper_clock = clock; // @[:@68825.4]
  assign RetimeWrapper_reset = reset; // @[:@68826.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@68828.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@68827.4]
  assign RetimeWrapper_1_clock = clock; // @[:@68833.4]
  assign RetimeWrapper_1_reset = reset; // @[:@68834.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@68836.4]
  assign RetimeWrapper_1_io_in = x740_sm_io_done; // @[package.scala 94:16:@68835.4]
  assign x740_kernelx740_concrete1_clock = clock; // @[:@68862.4]
  assign x740_kernelx740_concrete1_reset = reset; // @[:@68863.4]
  assign x740_kernelx740_concrete1_io_in_x340_outdram_number = io_in_x340_outdram_number; // @[sm_x740.scala 63:31:@68940.4]
  assign x740_kernelx740_concrete1_io_in_x344_outbuf_0_rPort_0_output_0 = x344_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@68941.4]
  assign x740_kernelx740_concrete1_io_in_x343_TREADY = io_in_x343_TREADY; // @[sm_x740.scala 65:23:@68953.4]
  assign x740_kernelx740_concrete1_io_in_x674_valid = io_in_x674_valid; // @[sm_x740.scala 66:23:@68956.4]
  assign x740_kernelx740_concrete1_io_in_x672_ready = io_in_x672_ready; // @[sm_x740.scala 67:23:@68961.4]
  assign x740_kernelx740_concrete1_io_in_x342_TVALID = io_in_x342_TVALID; // @[sm_x740.scala 68:23:@68970.4]
  assign x740_kernelx740_concrete1_io_in_x342_TDATA = io_in_x342_TDATA; // @[sm_x740.scala 68:23:@68968.4]
  assign x740_kernelx740_concrete1_io_in_x342_TID = io_in_x342_TID; // @[sm_x740.scala 68:23:@68964.4]
  assign x740_kernelx740_concrete1_io_in_x342_TDEST = io_in_x342_TDEST; // @[sm_x740.scala 68:23:@68963.4]
  assign x740_kernelx740_concrete1_io_in_x673_ready = io_in_x673_ready; // @[sm_x740.scala 69:23:@68974.4]
  assign x740_kernelx740_concrete1_io_sigsIn_smEnableOuts_0 = x740_sm_io_enableOut_0; // @[sm_x740.scala 107:22:@68985.4]
  assign x740_kernelx740_concrete1_io_sigsIn_smEnableOuts_1 = x740_sm_io_enableOut_1; // @[sm_x740.scala 107:22:@68986.4]
  assign x740_kernelx740_concrete1_io_sigsIn_smChildAcks_0 = x740_sm_io_childAck_0; // @[sm_x740.scala 107:22:@68981.4]
  assign x740_kernelx740_concrete1_io_sigsIn_smChildAcks_1 = x740_sm_io_childAck_1; // @[sm_x740.scala 107:22:@68982.4]
  assign x740_kernelx740_concrete1_io_rr = io_rr; // @[sm_x740.scala 106:18:@68975.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@69008.2]
  input          clock, // @[:@69009.4]
  input          reset, // @[:@69010.4]
  input          io_enable, // @[:@69011.4]
  output         io_done, // @[:@69011.4]
  input          io_reset, // @[:@69011.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@69011.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@69011.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@69011.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@69011.4]
  output         io_memStreams_loads_0_data_ready, // @[:@69011.4]
  input          io_memStreams_loads_0_data_valid, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@69011.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@69011.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@69011.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@69011.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@69011.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@69011.4]
  input          io_memStreams_stores_0_data_ready, // @[:@69011.4]
  output         io_memStreams_stores_0_data_valid, // @[:@69011.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@69011.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@69011.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@69011.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@69011.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@69011.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@69011.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@69011.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@69011.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@69011.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@69011.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@69011.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@69011.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@69011.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@69011.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@69011.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@69011.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@69011.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@69011.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@69011.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@69011.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@69011.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@69011.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@69011.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@69011.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@69011.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@69011.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@69011.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@69011.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@69011.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@69011.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@69011.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@69011.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@69011.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@69011.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@69011.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@69011.4]
  output         io_heap_0_req_valid, // @[:@69011.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@69011.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@69011.4]
  input          io_heap_0_resp_valid, // @[:@69011.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@69011.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@69011.4]
  input  [63:0]  io_argIns_0, // @[:@69011.4]
  input  [63:0]  io_argIns_1, // @[:@69011.4]
  input          io_argOuts_0_port_ready, // @[:@69011.4]
  output         io_argOuts_0_port_valid, // @[:@69011.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@69011.4]
  input  [63:0]  io_argOuts_0_echo // @[:@69011.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@69159.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@69159.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@69159.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@69159.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@69177.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@69177.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@69177.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@69177.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@69177.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@69186.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@69186.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@69186.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@69186.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@69186.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@69186.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@69225.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@69257.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@69257.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@69257.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@69257.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@69257.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@69319.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x340_outdram_number; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x343_TVALID; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x343_TREADY; // @[sm_RootController.scala 91:24:@69319.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x343_TDATA; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x674_ready; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x674_valid; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x672_ready; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x672_valid; // @[sm_RootController.scala 91:24:@69319.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x672_bits_addr; // @[sm_RootController.scala 91:24:@69319.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x672_bits_size; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x342_TVALID; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x342_TREADY; // @[sm_RootController.scala 91:24:@69319.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x342_TDATA; // @[sm_RootController.scala 91:24:@69319.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x342_TID; // @[sm_RootController.scala 91:24:@69319.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x342_TDEST; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x673_ready; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x673_valid; // @[sm_RootController.scala 91:24:@69319.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x673_bits_wdata_0; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_in_x673_bits_wstrb; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@69319.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@69319.4]
  wire  _T_599; // @[package.scala 96:25:@69182.4 package.scala 96:25:@69183.4]
  wire  _T_664; // @[Main.scala 46:50:@69253.4]
  wire  _T_665; // @[Main.scala 46:59:@69254.4]
  wire  _T_677; // @[package.scala 100:49:@69274.4]
  reg  _T_680; // @[package.scala 48:56:@69275.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@69159.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@69177.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@69186.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@69225.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@69257.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@69319.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x340_outdram_number(RootController_kernelRootController_concrete1_io_in_x340_outdram_number),
    .io_in_x343_TVALID(RootController_kernelRootController_concrete1_io_in_x343_TVALID),
    .io_in_x343_TREADY(RootController_kernelRootController_concrete1_io_in_x343_TREADY),
    .io_in_x343_TDATA(RootController_kernelRootController_concrete1_io_in_x343_TDATA),
    .io_in_x674_ready(RootController_kernelRootController_concrete1_io_in_x674_ready),
    .io_in_x674_valid(RootController_kernelRootController_concrete1_io_in_x674_valid),
    .io_in_x672_ready(RootController_kernelRootController_concrete1_io_in_x672_ready),
    .io_in_x672_valid(RootController_kernelRootController_concrete1_io_in_x672_valid),
    .io_in_x672_bits_addr(RootController_kernelRootController_concrete1_io_in_x672_bits_addr),
    .io_in_x672_bits_size(RootController_kernelRootController_concrete1_io_in_x672_bits_size),
    .io_in_x342_TVALID(RootController_kernelRootController_concrete1_io_in_x342_TVALID),
    .io_in_x342_TREADY(RootController_kernelRootController_concrete1_io_in_x342_TREADY),
    .io_in_x342_TDATA(RootController_kernelRootController_concrete1_io_in_x342_TDATA),
    .io_in_x342_TID(RootController_kernelRootController_concrete1_io_in_x342_TID),
    .io_in_x342_TDEST(RootController_kernelRootController_concrete1_io_in_x342_TDEST),
    .io_in_x673_ready(RootController_kernelRootController_concrete1_io_in_x673_ready),
    .io_in_x673_valid(RootController_kernelRootController_concrete1_io_in_x673_valid),
    .io_in_x673_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x673_bits_wdata_0),
    .io_in_x673_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x673_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@69182.4 package.scala 96:25:@69183.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@69253.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@69254.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@69274.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@69273.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x672_valid; // @[sm_RootController.scala 63:23:@69395.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x672_bits_addr; // @[sm_RootController.scala 63:23:@69394.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x672_bits_size; // @[sm_RootController.scala 63:23:@69393.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x673_valid; // @[sm_RootController.scala 65:23:@69408.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x673_bits_wdata_0; // @[sm_RootController.scala 65:23:@69407.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x673_bits_wstrb; // @[sm_RootController.scala 65:23:@69406.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x674_ready; // @[sm_RootController.scala 62:23:@69392.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x342_TREADY; // @[sm_RootController.scala 64:23:@69404.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x343_TVALID; // @[sm_RootController.scala 61:23:@69389.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x343_TDATA; // @[sm_RootController.scala 61:23:@69387.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 61:23:@69386.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 61:23:@69385.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 61:23:@69384.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 61:23:@69383.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 61:23:@69382.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 61:23:@69381.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@69160.4]
  assign SingleCounter_reset = reset; // @[:@69161.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@69175.4]
  assign RetimeWrapper_clock = clock; // @[:@69178.4]
  assign RetimeWrapper_reset = reset; // @[:@69179.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@69181.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@69180.4]
  assign SRFF_clock = clock; // @[:@69187.4]
  assign SRFF_reset = reset; // @[:@69188.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@69437.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@69271.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@69272.4]
  assign RootController_sm_clock = clock; // @[:@69226.4]
  assign RootController_sm_reset = reset; // @[:@69227.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@69270.4 SpatialBlocks.scala 140:18:@69304.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@69298.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@69278.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@69266.4 SpatialBlocks.scala 142:21:@69306.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@69295.4]
  assign RetimeWrapper_1_clock = clock; // @[:@69258.4]
  assign RetimeWrapper_1_reset = reset; // @[:@69259.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@69261.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@69260.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@69320.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@69321.4]
  assign RootController_kernelRootController_concrete1_io_in_x340_outdram_number = io_argIns_1; // @[sm_RootController.scala 60:31:@69380.4]
  assign RootController_kernelRootController_concrete1_io_in_x343_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 61:23:@69388.4]
  assign RootController_kernelRootController_concrete1_io_in_x674_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 62:23:@69391.4]
  assign RootController_kernelRootController_concrete1_io_in_x672_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 63:23:@69396.4]
  assign RootController_kernelRootController_concrete1_io_in_x342_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 64:23:@69405.4]
  assign RootController_kernelRootController_concrete1_io_in_x342_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 64:23:@69403.4]
  assign RootController_kernelRootController_concrete1_io_in_x342_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 64:23:@69399.4]
  assign RootController_kernelRootController_concrete1_io_in_x342_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 64:23:@69398.4]
  assign RootController_kernelRootController_concrete1_io_in_x673_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 65:23:@69409.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@69418.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@69416.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@69410.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@69439.2]
  input        clock, // @[:@69440.4]
  input        reset, // @[:@69441.4]
  input        io_enable, // @[:@69442.4]
  output [5:0] io_out, // @[:@69442.4]
  output [5:0] io_next // @[:@69442.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@69444.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@69445.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@69446.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@69451.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@69445.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@69446.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@69451.6]
  assign io_out = count; // @[Counter.scala 25:10:@69454.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@69455.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_49( // @[:@69491.2]
  input         clock, // @[:@69492.4]
  input         reset, // @[:@69493.4]
  input  [5:0]  io_raddr, // @[:@69494.4]
  input         io_wen, // @[:@69494.4]
  input  [5:0]  io_waddr, // @[:@69494.4]
  input  [63:0] io_wdata_addr, // @[:@69494.4]
  input  [31:0] io_wdata_size, // @[:@69494.4]
  output [63:0] io_rdata_addr, // @[:@69494.4]
  output [31:0] io_rdata_size // @[:@69494.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@69496.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@69496.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@69496.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@69496.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@69496.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@69496.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@69496.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@69496.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@69496.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@69510.4]
  wire  _T_20; // @[SRAM.scala 182:49:@69515.4]
  wire  _T_21; // @[SRAM.scala 182:37:@69516.4]
  reg  _T_24; // @[SRAM.scala 182:29:@69517.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@69520.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@69522.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@69496.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@69510.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@69515.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@69516.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@69522.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@69531.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@69530.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@69511.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@69512.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@69508.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@69514.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@69513.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@69509.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@69507.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@69506.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@69533.2]
  input         clock, // @[:@69534.4]
  input         reset, // @[:@69535.4]
  output        io_in_ready, // @[:@69536.4]
  input         io_in_valid, // @[:@69536.4]
  input  [63:0] io_in_bits_addr, // @[:@69536.4]
  input  [31:0] io_in_bits_size, // @[:@69536.4]
  input         io_out_ready, // @[:@69536.4]
  output        io_out_valid, // @[:@69536.4]
  output [63:0] io_out_bits_addr, // @[:@69536.4]
  output [31:0] io_out_bits_size // @[:@69536.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@69932.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@69932.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@69932.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@69932.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@69932.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@69942.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@69942.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@69942.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@69942.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@69942.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@69957.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@69957.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@69957.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@69957.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@69957.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@69957.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@69957.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@69957.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@69957.4]
  wire  writeEn; // @[FIFO.scala 30:29:@69930.4]
  wire  readEn; // @[FIFO.scala 31:29:@69931.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@69952.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@69953.4]
  wire  _T_824; // @[FIFO.scala 45:27:@69954.4]
  wire  empty; // @[FIFO.scala 45:24:@69955.4]
  wire  full; // @[FIFO.scala 46:23:@69956.4]
  wire  _T_827; // @[FIFO.scala 83:17:@69969.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@69970.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@69932.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@69942.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_49 SRAM ( // @[FIFO.scala 73:19:@69957.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@69930.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@69931.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@69953.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@69954.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@69955.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@69956.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@69969.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@69970.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@69976.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@69974.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@69967.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@69966.4]
  assign enqCounter_clock = clock; // @[:@69933.4]
  assign enqCounter_reset = reset; // @[:@69934.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@69940.4]
  assign deqCounter_clock = clock; // @[:@69943.4]
  assign deqCounter_reset = reset; // @[:@69944.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@69950.4]
  assign SRAM_clock = clock; // @[:@69958.4]
  assign SRAM_reset = reset; // @[:@69959.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@69961.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@69962.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@69963.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@69965.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@69964.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@69978.2]
  input        clock, // @[:@69979.4]
  input        reset, // @[:@69980.4]
  input        io_enable, // @[:@69981.4]
  output [3:0] io_out // @[:@69981.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@69983.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@69984.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@69985.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@69990.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@69984.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@69985.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@69990.6]
  assign io_out = count; // @[Counter.scala 25:10:@69993.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@70014.2]
  input        clock, // @[:@70015.4]
  input        reset, // @[:@70016.4]
  input        io_reset, // @[:@70017.4]
  input        io_enable, // @[:@70017.4]
  input  [1:0] io_stride, // @[:@70017.4]
  output [1:0] io_out, // @[:@70017.4]
  output [1:0] io_next // @[:@70017.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@70019.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@70020.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@70021.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@70026.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@70022.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@70020.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@70021.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@70026.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@70022.4]
  assign io_out = count; // @[Counter.scala 25:10:@70029.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@70030.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_50( // @[:@70066.2]
  input         clock, // @[:@70067.4]
  input         reset, // @[:@70068.4]
  input  [1:0]  io_raddr, // @[:@70069.4]
  input         io_wen, // @[:@70069.4]
  input  [1:0]  io_waddr, // @[:@70069.4]
  input  [31:0] io_wdata, // @[:@70069.4]
  output [31:0] io_rdata, // @[:@70069.4]
  input         io_backpressure // @[:@70069.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@70071.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@70071.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@70071.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@70071.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@70071.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@70071.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@70071.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@70071.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@70071.4]
  wire  _T_19; // @[SRAM.scala 182:49:@70089.4]
  wire  _T_20; // @[SRAM.scala 182:37:@70090.4]
  reg  _T_23; // @[SRAM.scala 182:29:@70091.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@70093.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@70071.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@70089.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@70090.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@70098.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@70085.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@70086.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@70083.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@70088.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@70087.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@70084.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@70082.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@70081.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@70100.2]
  input         clock, // @[:@70101.4]
  input         reset, // @[:@70102.4]
  output        io_in_ready, // @[:@70103.4]
  input         io_in_valid, // @[:@70103.4]
  input  [31:0] io_in_bits, // @[:@70103.4]
  input         io_out_ready, // @[:@70103.4]
  output        io_out_valid, // @[:@70103.4]
  output [31:0] io_out_bits // @[:@70103.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@70129.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@70129.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@70129.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@70129.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@70129.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@70129.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@70129.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@70139.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@70139.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@70139.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@70139.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@70139.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@70139.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@70139.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@70154.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@70154.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@70154.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@70154.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@70154.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@70154.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@70154.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@70154.4]
  wire  writeEn; // @[FIFO.scala 30:29:@70127.4]
  wire  readEn; // @[FIFO.scala 31:29:@70128.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@70149.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@70150.4]
  wire  _T_104; // @[FIFO.scala 45:27:@70151.4]
  wire  empty; // @[FIFO.scala 45:24:@70152.4]
  wire  full; // @[FIFO.scala 46:23:@70153.4]
  wire  _T_107; // @[FIFO.scala 83:17:@70164.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@70165.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@70129.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@70139.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_50 SRAM ( // @[FIFO.scala 73:19:@70154.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@70127.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@70128.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@70150.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@70151.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@70152.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@70153.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@70164.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@70165.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@70171.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@70169.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@70162.4]
  assign enqCounter_clock = clock; // @[:@70130.4]
  assign enqCounter_reset = reset; // @[:@70131.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@70137.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@70138.4]
  assign deqCounter_clock = clock; // @[:@70140.4]
  assign deqCounter_reset = reset; // @[:@70141.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@70147.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@70148.4]
  assign SRAM_clock = clock; // @[:@70155.4]
  assign SRAM_reset = reset; // @[:@70156.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@70158.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@70159.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@70160.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@70161.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@70163.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@72558.2]
  input         clock, // @[:@72559.4]
  input         reset, // @[:@72560.4]
  output        io_in_ready, // @[:@72561.4]
  input         io_in_valid, // @[:@72561.4]
  input  [31:0] io_in_bits_0, // @[:@72561.4]
  input         io_out_ready, // @[:@72561.4]
  output        io_out_valid, // @[:@72561.4]
  output [31:0] io_out_bits_0, // @[:@72561.4]
  output [31:0] io_out_bits_1, // @[:@72561.4]
  output [31:0] io_out_bits_2, // @[:@72561.4]
  output [31:0] io_out_bits_3, // @[:@72561.4]
  output [31:0] io_out_bits_4, // @[:@72561.4]
  output [31:0] io_out_bits_5, // @[:@72561.4]
  output [31:0] io_out_bits_6, // @[:@72561.4]
  output [31:0] io_out_bits_7, // @[:@72561.4]
  output [31:0] io_out_bits_8, // @[:@72561.4]
  output [31:0] io_out_bits_9, // @[:@72561.4]
  output [31:0] io_out_bits_10, // @[:@72561.4]
  output [31:0] io_out_bits_11, // @[:@72561.4]
  output [31:0] io_out_bits_12, // @[:@72561.4]
  output [31:0] io_out_bits_13, // @[:@72561.4]
  output [31:0] io_out_bits_14, // @[:@72561.4]
  output [31:0] io_out_bits_15 // @[:@72561.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@72565.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@72565.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@72565.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@72565.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@72576.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@72576.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@72576.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@72576.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@72589.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@72589.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@72589.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@72589.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@72589.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@72589.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@72589.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@72589.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@72624.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@72624.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@72624.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@72624.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@72624.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@72624.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@72624.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@72624.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@72659.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@72659.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@72659.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@72659.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@72659.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@72659.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@72659.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@72659.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@72694.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@72694.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@72694.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@72694.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@72694.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@72694.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@72694.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@72694.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@72729.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@72729.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@72729.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@72729.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@72729.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@72729.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@72729.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@72729.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@72764.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@72764.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@72764.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@72764.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@72764.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@72764.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@72764.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@72764.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@72799.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@72799.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@72799.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@72799.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@72799.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@72799.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@72799.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@72799.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@72834.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@72834.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@72834.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@72834.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@72834.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@72834.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@72834.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@72834.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@72869.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@72869.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@72869.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@72869.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@72869.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@72869.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@72869.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@72869.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@72904.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@72904.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@72904.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@72904.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@72904.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@72904.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@72904.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@72904.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@72939.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@72939.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@72939.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@72939.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@72939.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@72939.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@72939.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@72939.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@72974.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@72974.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@72974.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@72974.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@72974.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@72974.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@72974.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@72974.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@73009.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@73009.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@73009.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@73009.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@73009.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@73009.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@73009.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@73009.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@73044.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@73044.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@73044.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@73044.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@73044.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@73044.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@73044.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@73044.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@73079.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@73079.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@73079.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@73079.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@73079.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@73079.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@73079.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@73079.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@73114.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@73114.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@73114.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@73114.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@73114.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@73114.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@73114.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@73114.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@72564.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@72587.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@72614.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@72649.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@72684.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@72719.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@72754.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@72789.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@72824.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@72859.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@72894.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@72929.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@72964.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@72999.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@73034.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@73069.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@73104.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@73139.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73150.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73151.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73152.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73153.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73154.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73155.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73156.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73157.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73158.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73159.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73160.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73161.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73162.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73163.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73164.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@73181.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73165.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@73200.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@73201.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@73202.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@73203.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@73204.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@73205.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@73206.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@73207.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@73208.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@73209.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@73210.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@73211.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@73212.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@73213.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@72565.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@72576.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@72589.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@72624.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@72659.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@72694.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@72729.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@72764.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@72799.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@72834.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@72869.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@72904.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@72939.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@72974.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@73009.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@73044.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@73079.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@73114.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@72564.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@72587.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@72614.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@72649.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@72684.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@72719.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@72754.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@72789.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@72824.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@72859.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@72894.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@72929.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@72964.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@72999.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@73034.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@73069.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@73104.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@73139.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73150.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73151.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73152.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73153.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73154.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73155.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73156.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73157.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73158.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73159.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73160.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73161.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73162.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73163.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73164.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@73181.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@73149.4 FIFOVec.scala 49:42:@73165.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@73200.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@73201.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@73202.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@73203.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@73204.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@73205.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@73206.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@73207.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@73208.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@73209.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@73210.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@73211.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@73212.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@73213.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@73182.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@73216.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@73524.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@73525.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@73526.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@73527.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@73528.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@73529.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@73530.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@73531.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@73532.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@73533.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@73534.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@73535.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@73536.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@73537.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@73538.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@73539.4]
  assign enqCounter_clock = clock; // @[:@72566.4]
  assign enqCounter_reset = reset; // @[:@72567.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@72574.4]
  assign deqCounter_clock = clock; // @[:@72577.4]
  assign deqCounter_reset = reset; // @[:@72578.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@72585.4]
  assign fifos_0_clock = clock; // @[:@72590.4]
  assign fifos_0_reset = reset; // @[:@72591.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@72617.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72619.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72623.4]
  assign fifos_1_clock = clock; // @[:@72625.4]
  assign fifos_1_reset = reset; // @[:@72626.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@72652.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72654.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72658.4]
  assign fifos_2_clock = clock; // @[:@72660.4]
  assign fifos_2_reset = reset; // @[:@72661.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@72687.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72689.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72693.4]
  assign fifos_3_clock = clock; // @[:@72695.4]
  assign fifos_3_reset = reset; // @[:@72696.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@72722.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72724.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72728.4]
  assign fifos_4_clock = clock; // @[:@72730.4]
  assign fifos_4_reset = reset; // @[:@72731.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@72757.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72759.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72763.4]
  assign fifos_5_clock = clock; // @[:@72765.4]
  assign fifos_5_reset = reset; // @[:@72766.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@72792.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72794.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72798.4]
  assign fifos_6_clock = clock; // @[:@72800.4]
  assign fifos_6_reset = reset; // @[:@72801.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@72827.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72829.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72833.4]
  assign fifos_7_clock = clock; // @[:@72835.4]
  assign fifos_7_reset = reset; // @[:@72836.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@72862.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72864.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72868.4]
  assign fifos_8_clock = clock; // @[:@72870.4]
  assign fifos_8_reset = reset; // @[:@72871.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@72897.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72899.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72903.4]
  assign fifos_9_clock = clock; // @[:@72905.4]
  assign fifos_9_reset = reset; // @[:@72906.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@72932.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72934.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72938.4]
  assign fifos_10_clock = clock; // @[:@72940.4]
  assign fifos_10_reset = reset; // @[:@72941.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@72967.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@72969.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@72973.4]
  assign fifos_11_clock = clock; // @[:@72975.4]
  assign fifos_11_reset = reset; // @[:@72976.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@73002.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@73004.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@73008.4]
  assign fifos_12_clock = clock; // @[:@73010.4]
  assign fifos_12_reset = reset; // @[:@73011.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@73037.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@73039.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@73043.4]
  assign fifos_13_clock = clock; // @[:@73045.4]
  assign fifos_13_reset = reset; // @[:@73046.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@73072.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@73074.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@73078.4]
  assign fifos_14_clock = clock; // @[:@73080.4]
  assign fifos_14_reset = reset; // @[:@73081.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@73107.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@73109.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@73113.4]
  assign fifos_15_clock = clock; // @[:@73115.4]
  assign fifos_15_reset = reset; // @[:@73116.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@73142.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@73144.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@73148.4]
endmodule
module FFRAM( // @[:@73613.2]
  input        clock, // @[:@73614.4]
  input        reset, // @[:@73615.4]
  input  [1:0] io_raddr, // @[:@73616.4]
  input        io_wen, // @[:@73616.4]
  input  [1:0] io_waddr, // @[:@73616.4]
  input        io_wdata, // @[:@73616.4]
  output       io_rdata, // @[:@73616.4]
  input        io_banks_0_wdata_valid, // @[:@73616.4]
  input        io_banks_0_wdata_bits, // @[:@73616.4]
  input        io_banks_1_wdata_valid, // @[:@73616.4]
  input        io_banks_1_wdata_bits, // @[:@73616.4]
  input        io_banks_2_wdata_valid, // @[:@73616.4]
  input        io_banks_2_wdata_bits, // @[:@73616.4]
  input        io_banks_3_wdata_valid, // @[:@73616.4]
  input        io_banks_3_wdata_bits // @[:@73616.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@73620.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@73621.4]
  wire  _T_89; // @[SRAM.scala 148:25:@73622.4]
  wire  _T_90; // @[SRAM.scala 148:15:@73623.4]
  wire  _T_91; // @[SRAM.scala 149:15:@73625.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@73624.4]
  reg  regs_1; // @[SRAM.scala 145:20:@73631.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@73632.4]
  wire  _T_98; // @[SRAM.scala 148:25:@73633.4]
  wire  _T_99; // @[SRAM.scala 148:15:@73634.4]
  wire  _T_100; // @[SRAM.scala 149:15:@73636.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@73635.4]
  reg  regs_2; // @[SRAM.scala 145:20:@73642.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@73643.4]
  wire  _T_107; // @[SRAM.scala 148:25:@73644.4]
  wire  _T_108; // @[SRAM.scala 148:15:@73645.4]
  wire  _T_109; // @[SRAM.scala 149:15:@73647.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@73646.4]
  reg  regs_3; // @[SRAM.scala 145:20:@73653.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@73654.4]
  wire  _T_116; // @[SRAM.scala 148:25:@73655.4]
  wire  _T_117; // @[SRAM.scala 148:15:@73656.4]
  wire  _T_118; // @[SRAM.scala 149:15:@73658.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@73657.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@73667.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@73667.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@73621.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@73622.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@73623.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@73625.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@73624.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@73632.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@73633.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@73634.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@73636.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@73635.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@73643.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@73644.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@73645.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@73647.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@73646.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@73654.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@73655.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@73656.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@73658.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@73657.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@73667.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@73667.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@73667.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@73669.2]
  input   clock, // @[:@73670.4]
  input   reset, // @[:@73671.4]
  output  io_in_ready, // @[:@73672.4]
  input   io_in_valid, // @[:@73672.4]
  input   io_in_bits, // @[:@73672.4]
  input   io_out_ready, // @[:@73672.4]
  output  io_out_valid, // @[:@73672.4]
  output  io_out_bits // @[:@73672.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@73698.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@73698.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@73698.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@73698.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@73698.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@73698.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@73698.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@73708.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@73708.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@73708.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@73708.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@73708.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@73708.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@73708.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@73723.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@73723.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@73723.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@73723.4]
  wire  writeEn; // @[FIFO.scala 30:29:@73696.4]
  wire  readEn; // @[FIFO.scala 31:29:@73697.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@73718.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@73719.4]
  wire  _T_104; // @[FIFO.scala 45:27:@73720.4]
  wire  empty; // @[FIFO.scala 45:24:@73721.4]
  wire  full; // @[FIFO.scala 46:23:@73722.4]
  wire  _T_157; // @[FIFO.scala 83:17:@73809.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@73810.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@73698.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@73708.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@73723.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@73696.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@73697.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@73719.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@73720.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@73721.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@73722.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@73809.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@73810.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@73816.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@73814.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@73748.4]
  assign enqCounter_clock = clock; // @[:@73699.4]
  assign enqCounter_reset = reset; // @[:@73700.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@73706.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@73707.4]
  assign deqCounter_clock = clock; // @[:@73709.4]
  assign deqCounter_reset = reset; // @[:@73710.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@73716.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@73717.4]
  assign FFRAM_clock = clock; // @[:@73724.4]
  assign FFRAM_reset = reset; // @[:@73725.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@73744.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@73745.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@73746.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@73747.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@73750.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@73749.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@73753.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@73752.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@73756.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@73755.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@73759.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@73758.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@77433.2]
  input   clock, // @[:@77434.4]
  input   reset, // @[:@77435.4]
  output  io_in_ready, // @[:@77436.4]
  input   io_in_valid, // @[:@77436.4]
  input   io_in_bits_0, // @[:@77436.4]
  input   io_out_ready, // @[:@77436.4]
  output  io_out_valid, // @[:@77436.4]
  output  io_out_bits_0, // @[:@77436.4]
  output  io_out_bits_1, // @[:@77436.4]
  output  io_out_bits_2, // @[:@77436.4]
  output  io_out_bits_3, // @[:@77436.4]
  output  io_out_bits_4, // @[:@77436.4]
  output  io_out_bits_5, // @[:@77436.4]
  output  io_out_bits_6, // @[:@77436.4]
  output  io_out_bits_7, // @[:@77436.4]
  output  io_out_bits_8, // @[:@77436.4]
  output  io_out_bits_9, // @[:@77436.4]
  output  io_out_bits_10, // @[:@77436.4]
  output  io_out_bits_11, // @[:@77436.4]
  output  io_out_bits_12, // @[:@77436.4]
  output  io_out_bits_13, // @[:@77436.4]
  output  io_out_bits_14, // @[:@77436.4]
  output  io_out_bits_15 // @[:@77436.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@77440.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@77440.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@77440.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@77440.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@77451.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@77451.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@77451.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@77451.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@77464.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@77464.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@77464.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@77464.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@77464.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@77464.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@77464.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@77464.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@77499.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@77499.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@77499.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@77499.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@77499.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@77499.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@77499.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@77499.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@77534.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@77534.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@77534.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@77534.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@77534.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@77534.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@77534.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@77534.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@77569.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@77569.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@77569.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@77569.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@77569.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@77569.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@77569.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@77569.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@77604.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@77604.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@77604.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@77604.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@77604.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@77604.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@77604.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@77604.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@77639.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@77639.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@77639.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@77639.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@77639.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@77639.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@77639.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@77639.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@77674.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@77674.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@77674.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@77674.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@77674.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@77674.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@77674.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@77674.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@77709.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@77709.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@77709.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@77709.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@77709.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@77709.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@77709.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@77709.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@77744.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@77744.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@77744.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@77744.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@77744.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@77744.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@77744.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@77744.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@77779.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@77779.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@77779.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@77779.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@77779.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@77779.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@77779.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@77779.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@77814.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@77814.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@77814.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@77814.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@77814.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@77814.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@77814.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@77814.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@77849.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@77849.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@77849.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@77849.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@77849.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@77849.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@77849.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@77849.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@77884.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@77884.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@77884.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@77884.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@77884.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@77884.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@77884.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@77884.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@77919.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@77919.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@77919.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@77919.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@77919.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@77919.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@77919.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@77919.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@77954.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@77954.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@77954.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@77954.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@77954.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@77954.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@77954.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@77954.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@77989.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@77989.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@77989.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@77989.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@77989.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@77989.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@77989.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@77989.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@77439.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@77462.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@77489.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@77524.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@77559.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@77594.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@77629.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@77664.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@77699.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@77734.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@77769.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@77804.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@77839.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@77874.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@77909.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@77944.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@77979.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@78014.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78025.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78026.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78027.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78028.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78029.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78030.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78031.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78032.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78033.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78034.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78035.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78036.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78037.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78038.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78039.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@78056.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78040.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@78075.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@78076.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@78077.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@78078.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@78079.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@78080.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@78081.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@78082.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@78083.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@78084.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@78085.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@78086.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@78087.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@78088.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@77440.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@77451.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@77464.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@77499.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@77534.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@77569.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@77604.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@77639.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@77674.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@77709.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@77744.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@77779.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@77814.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@77849.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@77884.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@77919.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@77954.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@77989.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@77439.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@77462.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@77489.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@77524.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@77559.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@77594.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@77629.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@77664.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@77699.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@77734.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@77769.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@77804.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@77839.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@77874.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@77909.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@77944.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@77979.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@78014.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78025.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78026.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78027.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78028.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78029.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78030.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78031.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78032.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78033.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78034.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78035.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78036.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78037.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78038.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78039.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@78056.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@78024.4 FIFOVec.scala 49:42:@78040.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@78075.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@78076.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@78077.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@78078.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@78079.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@78080.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@78081.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@78082.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@78083.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@78084.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@78085.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@78086.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@78087.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@78088.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@78057.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@78091.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@78399.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@78400.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@78401.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@78402.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@78403.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@78404.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@78405.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@78406.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@78407.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@78408.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@78409.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@78410.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@78411.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@78412.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@78413.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@78414.4]
  assign enqCounter_clock = clock; // @[:@77441.4]
  assign enqCounter_reset = reset; // @[:@77442.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@77449.4]
  assign deqCounter_clock = clock; // @[:@77452.4]
  assign deqCounter_reset = reset; // @[:@77453.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@77460.4]
  assign fifos_0_clock = clock; // @[:@77465.4]
  assign fifos_0_reset = reset; // @[:@77466.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@77492.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77494.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77498.4]
  assign fifos_1_clock = clock; // @[:@77500.4]
  assign fifos_1_reset = reset; // @[:@77501.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@77527.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77529.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77533.4]
  assign fifos_2_clock = clock; // @[:@77535.4]
  assign fifos_2_reset = reset; // @[:@77536.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@77562.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77564.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77568.4]
  assign fifos_3_clock = clock; // @[:@77570.4]
  assign fifos_3_reset = reset; // @[:@77571.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@77597.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77599.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77603.4]
  assign fifos_4_clock = clock; // @[:@77605.4]
  assign fifos_4_reset = reset; // @[:@77606.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@77632.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77634.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77638.4]
  assign fifos_5_clock = clock; // @[:@77640.4]
  assign fifos_5_reset = reset; // @[:@77641.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@77667.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77669.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77673.4]
  assign fifos_6_clock = clock; // @[:@77675.4]
  assign fifos_6_reset = reset; // @[:@77676.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@77702.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77704.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77708.4]
  assign fifos_7_clock = clock; // @[:@77710.4]
  assign fifos_7_reset = reset; // @[:@77711.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@77737.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77739.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77743.4]
  assign fifos_8_clock = clock; // @[:@77745.4]
  assign fifos_8_reset = reset; // @[:@77746.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@77772.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77774.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77778.4]
  assign fifos_9_clock = clock; // @[:@77780.4]
  assign fifos_9_reset = reset; // @[:@77781.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@77807.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77809.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77813.4]
  assign fifos_10_clock = clock; // @[:@77815.4]
  assign fifos_10_reset = reset; // @[:@77816.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@77842.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77844.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77848.4]
  assign fifos_11_clock = clock; // @[:@77850.4]
  assign fifos_11_reset = reset; // @[:@77851.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@77877.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77879.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77883.4]
  assign fifos_12_clock = clock; // @[:@77885.4]
  assign fifos_12_reset = reset; // @[:@77886.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@77912.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77914.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77918.4]
  assign fifos_13_clock = clock; // @[:@77920.4]
  assign fifos_13_reset = reset; // @[:@77921.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@77947.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77949.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77953.4]
  assign fifos_14_clock = clock; // @[:@77955.4]
  assign fifos_14_reset = reset; // @[:@77956.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@77982.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@77984.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@77988.4]
  assign fifos_15_clock = clock; // @[:@77990.4]
  assign fifos_15_reset = reset; // @[:@77991.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@78017.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@78019.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@78023.4]
endmodule
module FIFOWidthConvert( // @[:@78416.2]
  input         clock, // @[:@78417.4]
  input         reset, // @[:@78418.4]
  output        io_in_ready, // @[:@78419.4]
  input         io_in_valid, // @[:@78419.4]
  input  [31:0] io_in_bits_data_0, // @[:@78419.4]
  input         io_in_bits_strobe, // @[:@78419.4]
  input         io_out_ready, // @[:@78419.4]
  output        io_out_valid, // @[:@78419.4]
  output [31:0] io_out_bits_data_0, // @[:@78419.4]
  output [31:0] io_out_bits_data_1, // @[:@78419.4]
  output [31:0] io_out_bits_data_2, // @[:@78419.4]
  output [31:0] io_out_bits_data_3, // @[:@78419.4]
  output [31:0] io_out_bits_data_4, // @[:@78419.4]
  output [31:0] io_out_bits_data_5, // @[:@78419.4]
  output [31:0] io_out_bits_data_6, // @[:@78419.4]
  output [31:0] io_out_bits_data_7, // @[:@78419.4]
  output [31:0] io_out_bits_data_8, // @[:@78419.4]
  output [31:0] io_out_bits_data_9, // @[:@78419.4]
  output [31:0] io_out_bits_data_10, // @[:@78419.4]
  output [31:0] io_out_bits_data_11, // @[:@78419.4]
  output [31:0] io_out_bits_data_12, // @[:@78419.4]
  output [31:0] io_out_bits_data_13, // @[:@78419.4]
  output [31:0] io_out_bits_data_14, // @[:@78419.4]
  output [31:0] io_out_bits_data_15, // @[:@78419.4]
  output [63:0] io_out_bits_strobe // @[:@78419.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@78421.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@78462.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@78521.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@78527.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@78585.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@78591.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@78592.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@78596.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@78600.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@78604.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@78608.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@78612.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@78616.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@78620.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@78624.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@78628.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@78632.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@78636.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@78640.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@78644.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@78648.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@78652.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@78729.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@78738.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@78747.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@78756.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@78765.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@78774.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@78782.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@78421.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@78462.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@78521.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@78527.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@78585.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@78591.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@78592.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@78596.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@78600.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@78604.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@78608.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@78612.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@78616.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@78620.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@78624.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@78628.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@78632.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@78636.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@78640.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@78644.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@78648.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@78652.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@78729.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@78738.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@78747.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@78756.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@78765.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@78774.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@78782.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@78511.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@78512.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@78561.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@78562.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@78563.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@78564.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@78565.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@78566.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@78567.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@78568.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@78569.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@78570.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@78571.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@78572.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@78573.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@78574.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@78575.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@78576.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@78784.4]
  assign FIFOVec_clock = clock; // @[:@78422.4]
  assign FIFOVec_reset = reset; // @[:@78423.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@78508.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@78507.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@78785.4]
  assign FIFOVec_1_clock = clock; // @[:@78463.4]
  assign FIFOVec_1_reset = reset; // @[:@78464.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@78510.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@78509.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@78786.4]
endmodule
module FFRAM_16( // @[:@78824.2]
  input        clock, // @[:@78825.4]
  input        reset, // @[:@78826.4]
  input  [5:0] io_raddr, // @[:@78827.4]
  input        io_wen, // @[:@78827.4]
  input  [5:0] io_waddr, // @[:@78827.4]
  input        io_wdata, // @[:@78827.4]
  output       io_rdata, // @[:@78827.4]
  input        io_banks_0_wdata_valid, // @[:@78827.4]
  input        io_banks_0_wdata_bits, // @[:@78827.4]
  input        io_banks_1_wdata_valid, // @[:@78827.4]
  input        io_banks_1_wdata_bits, // @[:@78827.4]
  input        io_banks_2_wdata_valid, // @[:@78827.4]
  input        io_banks_2_wdata_bits, // @[:@78827.4]
  input        io_banks_3_wdata_valid, // @[:@78827.4]
  input        io_banks_3_wdata_bits, // @[:@78827.4]
  input        io_banks_4_wdata_valid, // @[:@78827.4]
  input        io_banks_4_wdata_bits, // @[:@78827.4]
  input        io_banks_5_wdata_valid, // @[:@78827.4]
  input        io_banks_5_wdata_bits, // @[:@78827.4]
  input        io_banks_6_wdata_valid, // @[:@78827.4]
  input        io_banks_6_wdata_bits, // @[:@78827.4]
  input        io_banks_7_wdata_valid, // @[:@78827.4]
  input        io_banks_7_wdata_bits, // @[:@78827.4]
  input        io_banks_8_wdata_valid, // @[:@78827.4]
  input        io_banks_8_wdata_bits, // @[:@78827.4]
  input        io_banks_9_wdata_valid, // @[:@78827.4]
  input        io_banks_9_wdata_bits, // @[:@78827.4]
  input        io_banks_10_wdata_valid, // @[:@78827.4]
  input        io_banks_10_wdata_bits, // @[:@78827.4]
  input        io_banks_11_wdata_valid, // @[:@78827.4]
  input        io_banks_11_wdata_bits, // @[:@78827.4]
  input        io_banks_12_wdata_valid, // @[:@78827.4]
  input        io_banks_12_wdata_bits, // @[:@78827.4]
  input        io_banks_13_wdata_valid, // @[:@78827.4]
  input        io_banks_13_wdata_bits, // @[:@78827.4]
  input        io_banks_14_wdata_valid, // @[:@78827.4]
  input        io_banks_14_wdata_bits, // @[:@78827.4]
  input        io_banks_15_wdata_valid, // @[:@78827.4]
  input        io_banks_15_wdata_bits, // @[:@78827.4]
  input        io_banks_16_wdata_valid, // @[:@78827.4]
  input        io_banks_16_wdata_bits, // @[:@78827.4]
  input        io_banks_17_wdata_valid, // @[:@78827.4]
  input        io_banks_17_wdata_bits, // @[:@78827.4]
  input        io_banks_18_wdata_valid, // @[:@78827.4]
  input        io_banks_18_wdata_bits, // @[:@78827.4]
  input        io_banks_19_wdata_valid, // @[:@78827.4]
  input        io_banks_19_wdata_bits, // @[:@78827.4]
  input        io_banks_20_wdata_valid, // @[:@78827.4]
  input        io_banks_20_wdata_bits, // @[:@78827.4]
  input        io_banks_21_wdata_valid, // @[:@78827.4]
  input        io_banks_21_wdata_bits, // @[:@78827.4]
  input        io_banks_22_wdata_valid, // @[:@78827.4]
  input        io_banks_22_wdata_bits, // @[:@78827.4]
  input        io_banks_23_wdata_valid, // @[:@78827.4]
  input        io_banks_23_wdata_bits, // @[:@78827.4]
  input        io_banks_24_wdata_valid, // @[:@78827.4]
  input        io_banks_24_wdata_bits, // @[:@78827.4]
  input        io_banks_25_wdata_valid, // @[:@78827.4]
  input        io_banks_25_wdata_bits, // @[:@78827.4]
  input        io_banks_26_wdata_valid, // @[:@78827.4]
  input        io_banks_26_wdata_bits, // @[:@78827.4]
  input        io_banks_27_wdata_valid, // @[:@78827.4]
  input        io_banks_27_wdata_bits, // @[:@78827.4]
  input        io_banks_28_wdata_valid, // @[:@78827.4]
  input        io_banks_28_wdata_bits, // @[:@78827.4]
  input        io_banks_29_wdata_valid, // @[:@78827.4]
  input        io_banks_29_wdata_bits, // @[:@78827.4]
  input        io_banks_30_wdata_valid, // @[:@78827.4]
  input        io_banks_30_wdata_bits, // @[:@78827.4]
  input        io_banks_31_wdata_valid, // @[:@78827.4]
  input        io_banks_31_wdata_bits, // @[:@78827.4]
  input        io_banks_32_wdata_valid, // @[:@78827.4]
  input        io_banks_32_wdata_bits, // @[:@78827.4]
  input        io_banks_33_wdata_valid, // @[:@78827.4]
  input        io_banks_33_wdata_bits, // @[:@78827.4]
  input        io_banks_34_wdata_valid, // @[:@78827.4]
  input        io_banks_34_wdata_bits, // @[:@78827.4]
  input        io_banks_35_wdata_valid, // @[:@78827.4]
  input        io_banks_35_wdata_bits, // @[:@78827.4]
  input        io_banks_36_wdata_valid, // @[:@78827.4]
  input        io_banks_36_wdata_bits, // @[:@78827.4]
  input        io_banks_37_wdata_valid, // @[:@78827.4]
  input        io_banks_37_wdata_bits, // @[:@78827.4]
  input        io_banks_38_wdata_valid, // @[:@78827.4]
  input        io_banks_38_wdata_bits, // @[:@78827.4]
  input        io_banks_39_wdata_valid, // @[:@78827.4]
  input        io_banks_39_wdata_bits, // @[:@78827.4]
  input        io_banks_40_wdata_valid, // @[:@78827.4]
  input        io_banks_40_wdata_bits, // @[:@78827.4]
  input        io_banks_41_wdata_valid, // @[:@78827.4]
  input        io_banks_41_wdata_bits, // @[:@78827.4]
  input        io_banks_42_wdata_valid, // @[:@78827.4]
  input        io_banks_42_wdata_bits, // @[:@78827.4]
  input        io_banks_43_wdata_valid, // @[:@78827.4]
  input        io_banks_43_wdata_bits, // @[:@78827.4]
  input        io_banks_44_wdata_valid, // @[:@78827.4]
  input        io_banks_44_wdata_bits, // @[:@78827.4]
  input        io_banks_45_wdata_valid, // @[:@78827.4]
  input        io_banks_45_wdata_bits, // @[:@78827.4]
  input        io_banks_46_wdata_valid, // @[:@78827.4]
  input        io_banks_46_wdata_bits, // @[:@78827.4]
  input        io_banks_47_wdata_valid, // @[:@78827.4]
  input        io_banks_47_wdata_bits, // @[:@78827.4]
  input        io_banks_48_wdata_valid, // @[:@78827.4]
  input        io_banks_48_wdata_bits, // @[:@78827.4]
  input        io_banks_49_wdata_valid, // @[:@78827.4]
  input        io_banks_49_wdata_bits, // @[:@78827.4]
  input        io_banks_50_wdata_valid, // @[:@78827.4]
  input        io_banks_50_wdata_bits, // @[:@78827.4]
  input        io_banks_51_wdata_valid, // @[:@78827.4]
  input        io_banks_51_wdata_bits, // @[:@78827.4]
  input        io_banks_52_wdata_valid, // @[:@78827.4]
  input        io_banks_52_wdata_bits, // @[:@78827.4]
  input        io_banks_53_wdata_valid, // @[:@78827.4]
  input        io_banks_53_wdata_bits, // @[:@78827.4]
  input        io_banks_54_wdata_valid, // @[:@78827.4]
  input        io_banks_54_wdata_bits, // @[:@78827.4]
  input        io_banks_55_wdata_valid, // @[:@78827.4]
  input        io_banks_55_wdata_bits, // @[:@78827.4]
  input        io_banks_56_wdata_valid, // @[:@78827.4]
  input        io_banks_56_wdata_bits, // @[:@78827.4]
  input        io_banks_57_wdata_valid, // @[:@78827.4]
  input        io_banks_57_wdata_bits, // @[:@78827.4]
  input        io_banks_58_wdata_valid, // @[:@78827.4]
  input        io_banks_58_wdata_bits, // @[:@78827.4]
  input        io_banks_59_wdata_valid, // @[:@78827.4]
  input        io_banks_59_wdata_bits, // @[:@78827.4]
  input        io_banks_60_wdata_valid, // @[:@78827.4]
  input        io_banks_60_wdata_bits, // @[:@78827.4]
  input        io_banks_61_wdata_valid, // @[:@78827.4]
  input        io_banks_61_wdata_bits, // @[:@78827.4]
  input        io_banks_62_wdata_valid, // @[:@78827.4]
  input        io_banks_62_wdata_bits, // @[:@78827.4]
  input        io_banks_63_wdata_valid, // @[:@78827.4]
  input        io_banks_63_wdata_bits // @[:@78827.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@78831.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@78832.4]
  wire  _T_689; // @[SRAM.scala 148:25:@78833.4]
  wire  _T_690; // @[SRAM.scala 148:15:@78834.4]
  wire  _T_691; // @[SRAM.scala 149:15:@78836.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@78835.4]
  reg  regs_1; // @[SRAM.scala 145:20:@78842.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@78843.4]
  wire  _T_698; // @[SRAM.scala 148:25:@78844.4]
  wire  _T_699; // @[SRAM.scala 148:15:@78845.4]
  wire  _T_700; // @[SRAM.scala 149:15:@78847.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@78846.4]
  reg  regs_2; // @[SRAM.scala 145:20:@78853.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@78854.4]
  wire  _T_707; // @[SRAM.scala 148:25:@78855.4]
  wire  _T_708; // @[SRAM.scala 148:15:@78856.4]
  wire  _T_709; // @[SRAM.scala 149:15:@78858.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@78857.4]
  reg  regs_3; // @[SRAM.scala 145:20:@78864.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@78865.4]
  wire  _T_716; // @[SRAM.scala 148:25:@78866.4]
  wire  _T_717; // @[SRAM.scala 148:15:@78867.4]
  wire  _T_718; // @[SRAM.scala 149:15:@78869.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@78868.4]
  reg  regs_4; // @[SRAM.scala 145:20:@78875.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@78876.4]
  wire  _T_725; // @[SRAM.scala 148:25:@78877.4]
  wire  _T_726; // @[SRAM.scala 148:15:@78878.4]
  wire  _T_727; // @[SRAM.scala 149:15:@78880.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@78879.4]
  reg  regs_5; // @[SRAM.scala 145:20:@78886.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@78887.4]
  wire  _T_734; // @[SRAM.scala 148:25:@78888.4]
  wire  _T_735; // @[SRAM.scala 148:15:@78889.4]
  wire  _T_736; // @[SRAM.scala 149:15:@78891.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@78890.4]
  reg  regs_6; // @[SRAM.scala 145:20:@78897.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@78898.4]
  wire  _T_743; // @[SRAM.scala 148:25:@78899.4]
  wire  _T_744; // @[SRAM.scala 148:15:@78900.4]
  wire  _T_745; // @[SRAM.scala 149:15:@78902.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@78901.4]
  reg  regs_7; // @[SRAM.scala 145:20:@78908.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@78909.4]
  wire  _T_752; // @[SRAM.scala 148:25:@78910.4]
  wire  _T_753; // @[SRAM.scala 148:15:@78911.4]
  wire  _T_754; // @[SRAM.scala 149:15:@78913.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@78912.4]
  reg  regs_8; // @[SRAM.scala 145:20:@78919.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@78920.4]
  wire  _T_761; // @[SRAM.scala 148:25:@78921.4]
  wire  _T_762; // @[SRAM.scala 148:15:@78922.4]
  wire  _T_763; // @[SRAM.scala 149:15:@78924.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@78923.4]
  reg  regs_9; // @[SRAM.scala 145:20:@78930.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@78931.4]
  wire  _T_770; // @[SRAM.scala 148:25:@78932.4]
  wire  _T_771; // @[SRAM.scala 148:15:@78933.4]
  wire  _T_772; // @[SRAM.scala 149:15:@78935.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@78934.4]
  reg  regs_10; // @[SRAM.scala 145:20:@78941.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@78942.4]
  wire  _T_779; // @[SRAM.scala 148:25:@78943.4]
  wire  _T_780; // @[SRAM.scala 148:15:@78944.4]
  wire  _T_781; // @[SRAM.scala 149:15:@78946.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@78945.4]
  reg  regs_11; // @[SRAM.scala 145:20:@78952.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@78953.4]
  wire  _T_788; // @[SRAM.scala 148:25:@78954.4]
  wire  _T_789; // @[SRAM.scala 148:15:@78955.4]
  wire  _T_790; // @[SRAM.scala 149:15:@78957.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@78956.4]
  reg  regs_12; // @[SRAM.scala 145:20:@78963.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@78964.4]
  wire  _T_797; // @[SRAM.scala 148:25:@78965.4]
  wire  _T_798; // @[SRAM.scala 148:15:@78966.4]
  wire  _T_799; // @[SRAM.scala 149:15:@78968.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@78967.4]
  reg  regs_13; // @[SRAM.scala 145:20:@78974.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@78975.4]
  wire  _T_806; // @[SRAM.scala 148:25:@78976.4]
  wire  _T_807; // @[SRAM.scala 148:15:@78977.4]
  wire  _T_808; // @[SRAM.scala 149:15:@78979.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@78978.4]
  reg  regs_14; // @[SRAM.scala 145:20:@78985.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@78986.4]
  wire  _T_815; // @[SRAM.scala 148:25:@78987.4]
  wire  _T_816; // @[SRAM.scala 148:15:@78988.4]
  wire  _T_817; // @[SRAM.scala 149:15:@78990.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@78989.4]
  reg  regs_15; // @[SRAM.scala 145:20:@78996.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@78997.4]
  wire  _T_824; // @[SRAM.scala 148:25:@78998.4]
  wire  _T_825; // @[SRAM.scala 148:15:@78999.4]
  wire  _T_826; // @[SRAM.scala 149:15:@79001.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@79000.4]
  reg  regs_16; // @[SRAM.scala 145:20:@79007.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@79008.4]
  wire  _T_833; // @[SRAM.scala 148:25:@79009.4]
  wire  _T_834; // @[SRAM.scala 148:15:@79010.4]
  wire  _T_835; // @[SRAM.scala 149:15:@79012.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@79011.4]
  reg  regs_17; // @[SRAM.scala 145:20:@79018.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@79019.4]
  wire  _T_842; // @[SRAM.scala 148:25:@79020.4]
  wire  _T_843; // @[SRAM.scala 148:15:@79021.4]
  wire  _T_844; // @[SRAM.scala 149:15:@79023.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@79022.4]
  reg  regs_18; // @[SRAM.scala 145:20:@79029.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@79030.4]
  wire  _T_851; // @[SRAM.scala 148:25:@79031.4]
  wire  _T_852; // @[SRAM.scala 148:15:@79032.4]
  wire  _T_853; // @[SRAM.scala 149:15:@79034.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@79033.4]
  reg  regs_19; // @[SRAM.scala 145:20:@79040.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@79041.4]
  wire  _T_860; // @[SRAM.scala 148:25:@79042.4]
  wire  _T_861; // @[SRAM.scala 148:15:@79043.4]
  wire  _T_862; // @[SRAM.scala 149:15:@79045.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@79044.4]
  reg  regs_20; // @[SRAM.scala 145:20:@79051.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@79052.4]
  wire  _T_869; // @[SRAM.scala 148:25:@79053.4]
  wire  _T_870; // @[SRAM.scala 148:15:@79054.4]
  wire  _T_871; // @[SRAM.scala 149:15:@79056.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@79055.4]
  reg  regs_21; // @[SRAM.scala 145:20:@79062.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@79063.4]
  wire  _T_878; // @[SRAM.scala 148:25:@79064.4]
  wire  _T_879; // @[SRAM.scala 148:15:@79065.4]
  wire  _T_880; // @[SRAM.scala 149:15:@79067.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@79066.4]
  reg  regs_22; // @[SRAM.scala 145:20:@79073.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@79074.4]
  wire  _T_887; // @[SRAM.scala 148:25:@79075.4]
  wire  _T_888; // @[SRAM.scala 148:15:@79076.4]
  wire  _T_889; // @[SRAM.scala 149:15:@79078.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@79077.4]
  reg  regs_23; // @[SRAM.scala 145:20:@79084.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@79085.4]
  wire  _T_896; // @[SRAM.scala 148:25:@79086.4]
  wire  _T_897; // @[SRAM.scala 148:15:@79087.4]
  wire  _T_898; // @[SRAM.scala 149:15:@79089.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@79088.4]
  reg  regs_24; // @[SRAM.scala 145:20:@79095.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@79096.4]
  wire  _T_905; // @[SRAM.scala 148:25:@79097.4]
  wire  _T_906; // @[SRAM.scala 148:15:@79098.4]
  wire  _T_907; // @[SRAM.scala 149:15:@79100.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@79099.4]
  reg  regs_25; // @[SRAM.scala 145:20:@79106.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@79107.4]
  wire  _T_914; // @[SRAM.scala 148:25:@79108.4]
  wire  _T_915; // @[SRAM.scala 148:15:@79109.4]
  wire  _T_916; // @[SRAM.scala 149:15:@79111.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@79110.4]
  reg  regs_26; // @[SRAM.scala 145:20:@79117.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@79118.4]
  wire  _T_923; // @[SRAM.scala 148:25:@79119.4]
  wire  _T_924; // @[SRAM.scala 148:15:@79120.4]
  wire  _T_925; // @[SRAM.scala 149:15:@79122.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@79121.4]
  reg  regs_27; // @[SRAM.scala 145:20:@79128.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@79129.4]
  wire  _T_932; // @[SRAM.scala 148:25:@79130.4]
  wire  _T_933; // @[SRAM.scala 148:15:@79131.4]
  wire  _T_934; // @[SRAM.scala 149:15:@79133.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@79132.4]
  reg  regs_28; // @[SRAM.scala 145:20:@79139.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@79140.4]
  wire  _T_941; // @[SRAM.scala 148:25:@79141.4]
  wire  _T_942; // @[SRAM.scala 148:15:@79142.4]
  wire  _T_943; // @[SRAM.scala 149:15:@79144.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@79143.4]
  reg  regs_29; // @[SRAM.scala 145:20:@79150.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@79151.4]
  wire  _T_950; // @[SRAM.scala 148:25:@79152.4]
  wire  _T_951; // @[SRAM.scala 148:15:@79153.4]
  wire  _T_952; // @[SRAM.scala 149:15:@79155.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@79154.4]
  reg  regs_30; // @[SRAM.scala 145:20:@79161.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@79162.4]
  wire  _T_959; // @[SRAM.scala 148:25:@79163.4]
  wire  _T_960; // @[SRAM.scala 148:15:@79164.4]
  wire  _T_961; // @[SRAM.scala 149:15:@79166.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@79165.4]
  reg  regs_31; // @[SRAM.scala 145:20:@79172.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@79173.4]
  wire  _T_968; // @[SRAM.scala 148:25:@79174.4]
  wire  _T_969; // @[SRAM.scala 148:15:@79175.4]
  wire  _T_970; // @[SRAM.scala 149:15:@79177.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@79176.4]
  reg  regs_32; // @[SRAM.scala 145:20:@79183.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@79184.4]
  wire  _T_977; // @[SRAM.scala 148:25:@79185.4]
  wire  _T_978; // @[SRAM.scala 148:15:@79186.4]
  wire  _T_979; // @[SRAM.scala 149:15:@79188.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@79187.4]
  reg  regs_33; // @[SRAM.scala 145:20:@79194.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@79195.4]
  wire  _T_986; // @[SRAM.scala 148:25:@79196.4]
  wire  _T_987; // @[SRAM.scala 148:15:@79197.4]
  wire  _T_988; // @[SRAM.scala 149:15:@79199.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@79198.4]
  reg  regs_34; // @[SRAM.scala 145:20:@79205.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@79206.4]
  wire  _T_995; // @[SRAM.scala 148:25:@79207.4]
  wire  _T_996; // @[SRAM.scala 148:15:@79208.4]
  wire  _T_997; // @[SRAM.scala 149:15:@79210.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@79209.4]
  reg  regs_35; // @[SRAM.scala 145:20:@79216.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@79217.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@79218.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@79219.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@79221.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@79220.4]
  reg  regs_36; // @[SRAM.scala 145:20:@79227.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@79228.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@79229.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@79230.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@79232.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@79231.4]
  reg  regs_37; // @[SRAM.scala 145:20:@79238.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@79239.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@79240.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@79241.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@79243.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@79242.4]
  reg  regs_38; // @[SRAM.scala 145:20:@79249.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@79250.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@79251.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@79252.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@79254.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@79253.4]
  reg  regs_39; // @[SRAM.scala 145:20:@79260.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@79261.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@79262.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@79263.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@79265.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@79264.4]
  reg  regs_40; // @[SRAM.scala 145:20:@79271.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@79272.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@79273.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@79274.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@79276.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@79275.4]
  reg  regs_41; // @[SRAM.scala 145:20:@79282.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@79283.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@79284.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@79285.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@79287.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@79286.4]
  reg  regs_42; // @[SRAM.scala 145:20:@79293.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@79294.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@79295.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@79296.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@79298.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@79297.4]
  reg  regs_43; // @[SRAM.scala 145:20:@79304.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@79305.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@79306.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@79307.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@79309.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@79308.4]
  reg  regs_44; // @[SRAM.scala 145:20:@79315.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@79316.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@79317.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@79318.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@79320.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@79319.4]
  reg  regs_45; // @[SRAM.scala 145:20:@79326.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@79327.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@79328.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@79329.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@79331.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@79330.4]
  reg  regs_46; // @[SRAM.scala 145:20:@79337.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@79338.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@79339.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@79340.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@79342.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@79341.4]
  reg  regs_47; // @[SRAM.scala 145:20:@79348.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@79349.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@79350.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@79351.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@79353.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@79352.4]
  reg  regs_48; // @[SRAM.scala 145:20:@79359.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@79360.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@79361.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@79362.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@79364.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@79363.4]
  reg  regs_49; // @[SRAM.scala 145:20:@79370.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@79371.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@79372.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@79373.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@79375.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@79374.4]
  reg  regs_50; // @[SRAM.scala 145:20:@79381.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@79382.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@79383.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@79384.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@79386.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@79385.4]
  reg  regs_51; // @[SRAM.scala 145:20:@79392.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@79393.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@79394.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@79395.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@79397.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@79396.4]
  reg  regs_52; // @[SRAM.scala 145:20:@79403.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@79404.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@79405.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@79406.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@79408.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@79407.4]
  reg  regs_53; // @[SRAM.scala 145:20:@79414.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@79415.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@79416.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@79417.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@79419.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@79418.4]
  reg  regs_54; // @[SRAM.scala 145:20:@79425.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@79426.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@79427.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@79428.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@79430.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@79429.4]
  reg  regs_55; // @[SRAM.scala 145:20:@79436.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@79437.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@79438.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@79439.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@79441.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@79440.4]
  reg  regs_56; // @[SRAM.scala 145:20:@79447.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@79448.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@79449.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@79450.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@79452.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@79451.4]
  reg  regs_57; // @[SRAM.scala 145:20:@79458.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@79459.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@79460.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@79461.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@79463.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@79462.4]
  reg  regs_58; // @[SRAM.scala 145:20:@79469.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@79470.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@79471.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@79472.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@79474.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@79473.4]
  reg  regs_59; // @[SRAM.scala 145:20:@79480.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@79481.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@79482.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@79483.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@79485.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@79484.4]
  reg  regs_60; // @[SRAM.scala 145:20:@79491.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@79492.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@79493.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@79494.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@79496.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@79495.4]
  reg  regs_61; // @[SRAM.scala 145:20:@79502.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@79503.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@79504.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@79505.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@79507.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@79506.4]
  reg  regs_62; // @[SRAM.scala 145:20:@79513.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@79514.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@79515.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@79516.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@79518.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@79517.4]
  reg  regs_63; // @[SRAM.scala 145:20:@79524.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@79525.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@79526.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@79527.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@79529.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@79528.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@79598.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@79598.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@78832.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@78833.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@78834.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78836.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@78835.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@78843.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@78844.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@78845.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78847.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@78846.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@78854.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@78855.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@78856.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78858.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@78857.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@78865.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@78866.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@78867.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78869.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@78868.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@78876.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@78877.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@78878.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78880.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@78879.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@78887.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@78888.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@78889.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78891.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@78890.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@78898.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@78899.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@78900.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78902.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@78901.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@78909.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@78910.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@78911.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78913.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@78912.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@78920.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@78921.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@78922.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78924.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@78923.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@78931.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@78932.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@78933.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78935.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@78934.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@78942.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@78943.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@78944.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78946.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@78945.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@78953.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@78954.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@78955.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78957.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@78956.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@78964.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@78965.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@78966.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78968.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@78967.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@78975.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@78976.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@78977.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78979.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@78978.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@78986.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@78987.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@78988.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@78990.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@78989.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@78997.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@78998.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@78999.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79001.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@79000.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@79008.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@79009.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@79010.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79012.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@79011.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@79019.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@79020.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@79021.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79023.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@79022.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@79030.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@79031.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@79032.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79034.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@79033.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@79041.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@79042.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@79043.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79045.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@79044.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@79052.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@79053.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@79054.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79056.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@79055.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@79063.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@79064.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@79065.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79067.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@79066.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@79074.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@79075.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@79076.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79078.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@79077.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@79085.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@79086.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@79087.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79089.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@79088.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@79096.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@79097.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@79098.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79100.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@79099.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@79107.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@79108.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@79109.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79111.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@79110.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@79118.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@79119.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@79120.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79122.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@79121.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@79129.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@79130.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@79131.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79133.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@79132.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@79140.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@79141.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@79142.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79144.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@79143.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@79151.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@79152.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@79153.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79155.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@79154.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@79162.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@79163.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@79164.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79166.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@79165.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@79173.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@79174.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@79175.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79177.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@79176.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@79184.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@79185.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@79186.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79188.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@79187.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@79195.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@79196.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@79197.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79199.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@79198.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@79206.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@79207.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@79208.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79210.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@79209.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@79217.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@79218.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@79219.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79221.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@79220.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@79228.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@79229.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@79230.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79232.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@79231.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@79239.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@79240.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@79241.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79243.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@79242.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@79250.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@79251.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@79252.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79254.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@79253.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@79261.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@79262.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@79263.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79265.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@79264.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@79272.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@79273.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@79274.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79276.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@79275.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@79283.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@79284.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@79285.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79287.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@79286.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@79294.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@79295.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@79296.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79298.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@79297.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@79305.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@79306.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@79307.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79309.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@79308.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@79316.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@79317.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@79318.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79320.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@79319.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@79327.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@79328.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@79329.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79331.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@79330.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@79338.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@79339.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@79340.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79342.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@79341.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@79349.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@79350.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@79351.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79353.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@79352.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@79360.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@79361.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@79362.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79364.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@79363.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@79371.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@79372.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@79373.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79375.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@79374.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@79382.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@79383.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@79384.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79386.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@79385.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@79393.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@79394.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@79395.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79397.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@79396.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@79404.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@79405.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@79406.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79408.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@79407.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@79415.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@79416.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@79417.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79419.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@79418.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@79426.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@79427.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@79428.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79430.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@79429.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@79437.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@79438.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@79439.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79441.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@79440.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@79448.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@79449.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@79450.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79452.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@79451.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@79459.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@79460.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@79461.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79463.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@79462.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@79470.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@79471.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@79472.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79474.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@79473.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@79481.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@79482.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@79483.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79485.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@79484.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@79492.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@79493.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@79494.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79496.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@79495.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@79503.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@79504.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@79505.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79507.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@79506.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@79514.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@79515.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@79516.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79518.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@79517.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@79525.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@79526.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@79527.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@79529.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@79528.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@79598.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@79598.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@79598.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@79600.2]
  input   clock, // @[:@79601.4]
  input   reset, // @[:@79602.4]
  output  io_in_ready, // @[:@79603.4]
  input   io_in_valid, // @[:@79603.4]
  input   io_in_bits, // @[:@79603.4]
  input   io_out_ready, // @[:@79603.4]
  output  io_out_valid, // @[:@79603.4]
  output  io_out_bits, // @[:@79603.4]
  input   io_banks_0_wdata_valid, // @[:@79603.4]
  input   io_banks_0_wdata_bits, // @[:@79603.4]
  input   io_banks_1_wdata_valid, // @[:@79603.4]
  input   io_banks_1_wdata_bits, // @[:@79603.4]
  input   io_banks_2_wdata_valid, // @[:@79603.4]
  input   io_banks_2_wdata_bits, // @[:@79603.4]
  input   io_banks_3_wdata_valid, // @[:@79603.4]
  input   io_banks_3_wdata_bits, // @[:@79603.4]
  input   io_banks_4_wdata_valid, // @[:@79603.4]
  input   io_banks_4_wdata_bits, // @[:@79603.4]
  input   io_banks_5_wdata_valid, // @[:@79603.4]
  input   io_banks_5_wdata_bits, // @[:@79603.4]
  input   io_banks_6_wdata_valid, // @[:@79603.4]
  input   io_banks_6_wdata_bits, // @[:@79603.4]
  input   io_banks_7_wdata_valid, // @[:@79603.4]
  input   io_banks_7_wdata_bits, // @[:@79603.4]
  input   io_banks_8_wdata_valid, // @[:@79603.4]
  input   io_banks_8_wdata_bits, // @[:@79603.4]
  input   io_banks_9_wdata_valid, // @[:@79603.4]
  input   io_banks_9_wdata_bits, // @[:@79603.4]
  input   io_banks_10_wdata_valid, // @[:@79603.4]
  input   io_banks_10_wdata_bits, // @[:@79603.4]
  input   io_banks_11_wdata_valid, // @[:@79603.4]
  input   io_banks_11_wdata_bits, // @[:@79603.4]
  input   io_banks_12_wdata_valid, // @[:@79603.4]
  input   io_banks_12_wdata_bits, // @[:@79603.4]
  input   io_banks_13_wdata_valid, // @[:@79603.4]
  input   io_banks_13_wdata_bits, // @[:@79603.4]
  input   io_banks_14_wdata_valid, // @[:@79603.4]
  input   io_banks_14_wdata_bits, // @[:@79603.4]
  input   io_banks_15_wdata_valid, // @[:@79603.4]
  input   io_banks_15_wdata_bits, // @[:@79603.4]
  input   io_banks_16_wdata_valid, // @[:@79603.4]
  input   io_banks_16_wdata_bits, // @[:@79603.4]
  input   io_banks_17_wdata_valid, // @[:@79603.4]
  input   io_banks_17_wdata_bits, // @[:@79603.4]
  input   io_banks_18_wdata_valid, // @[:@79603.4]
  input   io_banks_18_wdata_bits, // @[:@79603.4]
  input   io_banks_19_wdata_valid, // @[:@79603.4]
  input   io_banks_19_wdata_bits, // @[:@79603.4]
  input   io_banks_20_wdata_valid, // @[:@79603.4]
  input   io_banks_20_wdata_bits, // @[:@79603.4]
  input   io_banks_21_wdata_valid, // @[:@79603.4]
  input   io_banks_21_wdata_bits, // @[:@79603.4]
  input   io_banks_22_wdata_valid, // @[:@79603.4]
  input   io_banks_22_wdata_bits, // @[:@79603.4]
  input   io_banks_23_wdata_valid, // @[:@79603.4]
  input   io_banks_23_wdata_bits, // @[:@79603.4]
  input   io_banks_24_wdata_valid, // @[:@79603.4]
  input   io_banks_24_wdata_bits, // @[:@79603.4]
  input   io_banks_25_wdata_valid, // @[:@79603.4]
  input   io_banks_25_wdata_bits, // @[:@79603.4]
  input   io_banks_26_wdata_valid, // @[:@79603.4]
  input   io_banks_26_wdata_bits, // @[:@79603.4]
  input   io_banks_27_wdata_valid, // @[:@79603.4]
  input   io_banks_27_wdata_bits, // @[:@79603.4]
  input   io_banks_28_wdata_valid, // @[:@79603.4]
  input   io_banks_28_wdata_bits, // @[:@79603.4]
  input   io_banks_29_wdata_valid, // @[:@79603.4]
  input   io_banks_29_wdata_bits, // @[:@79603.4]
  input   io_banks_30_wdata_valid, // @[:@79603.4]
  input   io_banks_30_wdata_bits, // @[:@79603.4]
  input   io_banks_31_wdata_valid, // @[:@79603.4]
  input   io_banks_31_wdata_bits, // @[:@79603.4]
  input   io_banks_32_wdata_valid, // @[:@79603.4]
  input   io_banks_32_wdata_bits, // @[:@79603.4]
  input   io_banks_33_wdata_valid, // @[:@79603.4]
  input   io_banks_33_wdata_bits, // @[:@79603.4]
  input   io_banks_34_wdata_valid, // @[:@79603.4]
  input   io_banks_34_wdata_bits, // @[:@79603.4]
  input   io_banks_35_wdata_valid, // @[:@79603.4]
  input   io_banks_35_wdata_bits, // @[:@79603.4]
  input   io_banks_36_wdata_valid, // @[:@79603.4]
  input   io_banks_36_wdata_bits, // @[:@79603.4]
  input   io_banks_37_wdata_valid, // @[:@79603.4]
  input   io_banks_37_wdata_bits, // @[:@79603.4]
  input   io_banks_38_wdata_valid, // @[:@79603.4]
  input   io_banks_38_wdata_bits, // @[:@79603.4]
  input   io_banks_39_wdata_valid, // @[:@79603.4]
  input   io_banks_39_wdata_bits, // @[:@79603.4]
  input   io_banks_40_wdata_valid, // @[:@79603.4]
  input   io_banks_40_wdata_bits, // @[:@79603.4]
  input   io_banks_41_wdata_valid, // @[:@79603.4]
  input   io_banks_41_wdata_bits, // @[:@79603.4]
  input   io_banks_42_wdata_valid, // @[:@79603.4]
  input   io_banks_42_wdata_bits, // @[:@79603.4]
  input   io_banks_43_wdata_valid, // @[:@79603.4]
  input   io_banks_43_wdata_bits, // @[:@79603.4]
  input   io_banks_44_wdata_valid, // @[:@79603.4]
  input   io_banks_44_wdata_bits, // @[:@79603.4]
  input   io_banks_45_wdata_valid, // @[:@79603.4]
  input   io_banks_45_wdata_bits, // @[:@79603.4]
  input   io_banks_46_wdata_valid, // @[:@79603.4]
  input   io_banks_46_wdata_bits, // @[:@79603.4]
  input   io_banks_47_wdata_valid, // @[:@79603.4]
  input   io_banks_47_wdata_bits, // @[:@79603.4]
  input   io_banks_48_wdata_valid, // @[:@79603.4]
  input   io_banks_48_wdata_bits, // @[:@79603.4]
  input   io_banks_49_wdata_valid, // @[:@79603.4]
  input   io_banks_49_wdata_bits, // @[:@79603.4]
  input   io_banks_50_wdata_valid, // @[:@79603.4]
  input   io_banks_50_wdata_bits, // @[:@79603.4]
  input   io_banks_51_wdata_valid, // @[:@79603.4]
  input   io_banks_51_wdata_bits, // @[:@79603.4]
  input   io_banks_52_wdata_valid, // @[:@79603.4]
  input   io_banks_52_wdata_bits, // @[:@79603.4]
  input   io_banks_53_wdata_valid, // @[:@79603.4]
  input   io_banks_53_wdata_bits, // @[:@79603.4]
  input   io_banks_54_wdata_valid, // @[:@79603.4]
  input   io_banks_54_wdata_bits, // @[:@79603.4]
  input   io_banks_55_wdata_valid, // @[:@79603.4]
  input   io_banks_55_wdata_bits, // @[:@79603.4]
  input   io_banks_56_wdata_valid, // @[:@79603.4]
  input   io_banks_56_wdata_bits, // @[:@79603.4]
  input   io_banks_57_wdata_valid, // @[:@79603.4]
  input   io_banks_57_wdata_bits, // @[:@79603.4]
  input   io_banks_58_wdata_valid, // @[:@79603.4]
  input   io_banks_58_wdata_bits, // @[:@79603.4]
  input   io_banks_59_wdata_valid, // @[:@79603.4]
  input   io_banks_59_wdata_bits, // @[:@79603.4]
  input   io_banks_60_wdata_valid, // @[:@79603.4]
  input   io_banks_60_wdata_bits, // @[:@79603.4]
  input   io_banks_61_wdata_valid, // @[:@79603.4]
  input   io_banks_61_wdata_bits, // @[:@79603.4]
  input   io_banks_62_wdata_valid, // @[:@79603.4]
  input   io_banks_62_wdata_bits, // @[:@79603.4]
  input   io_banks_63_wdata_valid, // @[:@79603.4]
  input   io_banks_63_wdata_bits // @[:@79603.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@79869.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@79869.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@79869.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@79869.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@79869.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@79879.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@79879.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@79879.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@79879.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@79879.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@79894.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@79894.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@79894.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@79894.4]
  wire  writeEn; // @[FIFO.scala 30:29:@79867.4]
  wire  readEn; // @[FIFO.scala 31:29:@79868.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@79889.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@79890.4]
  wire  _T_824; // @[FIFO.scala 45:27:@79891.4]
  wire  empty; // @[FIFO.scala 45:24:@79892.4]
  wire  full; // @[FIFO.scala 46:23:@79893.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@81060.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@81061.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@79869.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@79879.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@79894.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@79867.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@79868.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@79890.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@79891.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@79892.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@79893.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@81060.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@81061.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@81067.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@81065.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@80099.4]
  assign enqCounter_clock = clock; // @[:@79870.4]
  assign enqCounter_reset = reset; // @[:@79871.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@79877.4]
  assign deqCounter_clock = clock; // @[:@79880.4]
  assign deqCounter_reset = reset; // @[:@79881.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@79887.4]
  assign FFRAM_clock = clock; // @[:@79895.4]
  assign FFRAM_reset = reset; // @[:@79896.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@80095.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@80096.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@80097.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@80098.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@80101.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@80100.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@80104.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@80103.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@80107.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@80106.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@80110.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@80109.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@80113.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@80112.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@80116.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@80115.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@80119.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@80118.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@80122.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@80121.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@80125.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@80124.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@80128.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@80127.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@80131.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@80130.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@80134.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@80133.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@80137.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@80136.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@80140.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@80139.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@80143.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@80142.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@80146.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@80145.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@80149.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@80148.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@80152.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@80151.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@80155.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@80154.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@80158.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@80157.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@80161.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@80160.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@80164.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@80163.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@80167.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@80166.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@80170.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@80169.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@80173.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@80172.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@80176.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@80175.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@80179.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@80178.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@80182.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@80181.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@80185.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@80184.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@80188.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@80187.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@80191.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@80190.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@80194.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@80193.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@80197.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@80196.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@80200.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@80199.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@80203.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@80202.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@80206.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@80205.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@80209.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@80208.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@80212.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@80211.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@80215.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@80214.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@80218.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@80217.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@80221.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@80220.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@80224.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@80223.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@80227.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@80226.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@80230.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@80229.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@80233.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@80232.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@80236.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@80235.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@80239.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@80238.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@80242.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@80241.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@80245.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@80244.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@80248.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@80247.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@80251.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@80250.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@80254.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@80253.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@80257.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@80256.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@80260.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@80259.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@80263.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@80262.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@80266.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@80265.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@80269.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@80268.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@80272.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@80271.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@80275.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@80274.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@80278.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@80277.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@80281.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@80280.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@80284.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@80283.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@80287.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@80286.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@80290.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@80289.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@81069.2]
  input         clock, // @[:@81070.4]
  input         reset, // @[:@81071.4]
  input         io_dram_cmd_ready, // @[:@81072.4]
  output        io_dram_cmd_valid, // @[:@81072.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@81072.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@81072.4]
  input         io_dram_wdata_ready, // @[:@81072.4]
  output        io_dram_wdata_valid, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@81072.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@81072.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@81072.4]
  output        io_dram_wresp_ready, // @[:@81072.4]
  input         io_dram_wresp_valid, // @[:@81072.4]
  output        io_store_cmd_ready, // @[:@81072.4]
  input         io_store_cmd_valid, // @[:@81072.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@81072.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@81072.4]
  output        io_store_data_ready, // @[:@81072.4]
  input         io_store_data_valid, // @[:@81072.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@81072.4]
  input         io_store_data_bits_wstrb, // @[:@81072.4]
  input         io_store_wresp_ready, // @[:@81072.4]
  output        io_store_wresp_valid, // @[:@81072.4]
  output        io_store_wresp_bits // @[:@81072.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@81197.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@81197.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@81197.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@81197.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@81197.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@81197.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@81197.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@81197.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@81197.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@81197.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@81603.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@81603.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@81603.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@81603.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@81603.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@81603.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@81603.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@81603.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@81603.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@81844.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@81844.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@81600.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@81197.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@81603.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@81844.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@81600.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@81597.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@81598.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@81601.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@81633.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@81634.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@81635.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@81636.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@81637.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@81638.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@81639.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@81640.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@81641.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@81642.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@81643.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@81644.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@81645.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@81646.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@81647.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@81648.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@81649.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@81779.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@81780.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@81781.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@81782.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@81783.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@81784.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@81785.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@81786.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@81787.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@81788.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@81789.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@81790.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@81791.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@81792.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@81793.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@81794.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@81795.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@81796.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@81797.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@81798.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@81799.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@81800.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@81801.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@81802.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@81803.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@81804.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@81805.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@81806.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@81807.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@81808.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@81809.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@81810.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@81811.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@81812.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@81813.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@81814.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@81815.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@81816.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@81817.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@81818.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@81819.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@81820.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@81821.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@81822.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@81823.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@81824.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@81825.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@81826.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@81827.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@81828.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@81829.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@81830.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@81831.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@81832.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@81833.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@81834.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@81835.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@81836.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@81837.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@81838.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@81839.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@81840.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@81841.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@81842.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@82111.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@81595.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@81632.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@82112.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@82113.4]
  assign cmd_clock = clock; // @[:@81198.4]
  assign cmd_reset = reset; // @[:@81199.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@81592.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@81594.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@81593.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@81596.4]
  assign wdata_clock = clock; // @[:@81604.4]
  assign wdata_reset = reset; // @[:@81605.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@81629.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@81630.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@81631.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@81843.4]
  assign wresp_clock = clock; // @[:@81845.4]
  assign wresp_reset = reset; // @[:@81846.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@82109.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@82110.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@82114.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@82180.2]
  output        io_in_ready, // @[:@82183.4]
  input         io_in_valid, // @[:@82183.4]
  input  [63:0] io_in_bits_0_addr, // @[:@82183.4]
  input  [31:0] io_in_bits_0_size, // @[:@82183.4]
  input         io_in_bits_0_isWr, // @[:@82183.4]
  input  [31:0] io_in_bits_0_tag, // @[:@82183.4]
  input         io_out_ready, // @[:@82183.4]
  output        io_out_valid, // @[:@82183.4]
  output [63:0] io_out_bits_addr, // @[:@82183.4]
  output [31:0] io_out_bits_size, // @[:@82183.4]
  output        io_out_bits_isWr, // @[:@82183.4]
  output [31:0] io_out_bits_tag // @[:@82183.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@82185.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@82185.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@82194.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@82193.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@82199.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@82198.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@82196.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@82195.4]
endmodule
module MuxPipe_1( // @[:@82201.2]
  output        io_in_ready, // @[:@82204.4]
  input         io_in_valid, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@82204.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@82204.4]
  input         io_in_bits_0_wstrb_0, // @[:@82204.4]
  input         io_in_bits_0_wstrb_1, // @[:@82204.4]
  input         io_in_bits_0_wstrb_2, // @[:@82204.4]
  input         io_in_bits_0_wstrb_3, // @[:@82204.4]
  input         io_in_bits_0_wstrb_4, // @[:@82204.4]
  input         io_in_bits_0_wstrb_5, // @[:@82204.4]
  input         io_in_bits_0_wstrb_6, // @[:@82204.4]
  input         io_in_bits_0_wstrb_7, // @[:@82204.4]
  input         io_in_bits_0_wstrb_8, // @[:@82204.4]
  input         io_in_bits_0_wstrb_9, // @[:@82204.4]
  input         io_in_bits_0_wstrb_10, // @[:@82204.4]
  input         io_in_bits_0_wstrb_11, // @[:@82204.4]
  input         io_in_bits_0_wstrb_12, // @[:@82204.4]
  input         io_in_bits_0_wstrb_13, // @[:@82204.4]
  input         io_in_bits_0_wstrb_14, // @[:@82204.4]
  input         io_in_bits_0_wstrb_15, // @[:@82204.4]
  input         io_in_bits_0_wstrb_16, // @[:@82204.4]
  input         io_in_bits_0_wstrb_17, // @[:@82204.4]
  input         io_in_bits_0_wstrb_18, // @[:@82204.4]
  input         io_in_bits_0_wstrb_19, // @[:@82204.4]
  input         io_in_bits_0_wstrb_20, // @[:@82204.4]
  input         io_in_bits_0_wstrb_21, // @[:@82204.4]
  input         io_in_bits_0_wstrb_22, // @[:@82204.4]
  input         io_in_bits_0_wstrb_23, // @[:@82204.4]
  input         io_in_bits_0_wstrb_24, // @[:@82204.4]
  input         io_in_bits_0_wstrb_25, // @[:@82204.4]
  input         io_in_bits_0_wstrb_26, // @[:@82204.4]
  input         io_in_bits_0_wstrb_27, // @[:@82204.4]
  input         io_in_bits_0_wstrb_28, // @[:@82204.4]
  input         io_in_bits_0_wstrb_29, // @[:@82204.4]
  input         io_in_bits_0_wstrb_30, // @[:@82204.4]
  input         io_in_bits_0_wstrb_31, // @[:@82204.4]
  input         io_in_bits_0_wstrb_32, // @[:@82204.4]
  input         io_in_bits_0_wstrb_33, // @[:@82204.4]
  input         io_in_bits_0_wstrb_34, // @[:@82204.4]
  input         io_in_bits_0_wstrb_35, // @[:@82204.4]
  input         io_in_bits_0_wstrb_36, // @[:@82204.4]
  input         io_in_bits_0_wstrb_37, // @[:@82204.4]
  input         io_in_bits_0_wstrb_38, // @[:@82204.4]
  input         io_in_bits_0_wstrb_39, // @[:@82204.4]
  input         io_in_bits_0_wstrb_40, // @[:@82204.4]
  input         io_in_bits_0_wstrb_41, // @[:@82204.4]
  input         io_in_bits_0_wstrb_42, // @[:@82204.4]
  input         io_in_bits_0_wstrb_43, // @[:@82204.4]
  input         io_in_bits_0_wstrb_44, // @[:@82204.4]
  input         io_in_bits_0_wstrb_45, // @[:@82204.4]
  input         io_in_bits_0_wstrb_46, // @[:@82204.4]
  input         io_in_bits_0_wstrb_47, // @[:@82204.4]
  input         io_in_bits_0_wstrb_48, // @[:@82204.4]
  input         io_in_bits_0_wstrb_49, // @[:@82204.4]
  input         io_in_bits_0_wstrb_50, // @[:@82204.4]
  input         io_in_bits_0_wstrb_51, // @[:@82204.4]
  input         io_in_bits_0_wstrb_52, // @[:@82204.4]
  input         io_in_bits_0_wstrb_53, // @[:@82204.4]
  input         io_in_bits_0_wstrb_54, // @[:@82204.4]
  input         io_in_bits_0_wstrb_55, // @[:@82204.4]
  input         io_in_bits_0_wstrb_56, // @[:@82204.4]
  input         io_in_bits_0_wstrb_57, // @[:@82204.4]
  input         io_in_bits_0_wstrb_58, // @[:@82204.4]
  input         io_in_bits_0_wstrb_59, // @[:@82204.4]
  input         io_in_bits_0_wstrb_60, // @[:@82204.4]
  input         io_in_bits_0_wstrb_61, // @[:@82204.4]
  input         io_in_bits_0_wstrb_62, // @[:@82204.4]
  input         io_in_bits_0_wstrb_63, // @[:@82204.4]
  input         io_out_ready, // @[:@82204.4]
  output        io_out_valid, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_0, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_1, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_2, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_3, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_4, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_5, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_6, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_7, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_8, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_9, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_10, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_11, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_12, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_13, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_14, // @[:@82204.4]
  output [31:0] io_out_bits_wdata_15, // @[:@82204.4]
  output        io_out_bits_wstrb_0, // @[:@82204.4]
  output        io_out_bits_wstrb_1, // @[:@82204.4]
  output        io_out_bits_wstrb_2, // @[:@82204.4]
  output        io_out_bits_wstrb_3, // @[:@82204.4]
  output        io_out_bits_wstrb_4, // @[:@82204.4]
  output        io_out_bits_wstrb_5, // @[:@82204.4]
  output        io_out_bits_wstrb_6, // @[:@82204.4]
  output        io_out_bits_wstrb_7, // @[:@82204.4]
  output        io_out_bits_wstrb_8, // @[:@82204.4]
  output        io_out_bits_wstrb_9, // @[:@82204.4]
  output        io_out_bits_wstrb_10, // @[:@82204.4]
  output        io_out_bits_wstrb_11, // @[:@82204.4]
  output        io_out_bits_wstrb_12, // @[:@82204.4]
  output        io_out_bits_wstrb_13, // @[:@82204.4]
  output        io_out_bits_wstrb_14, // @[:@82204.4]
  output        io_out_bits_wstrb_15, // @[:@82204.4]
  output        io_out_bits_wstrb_16, // @[:@82204.4]
  output        io_out_bits_wstrb_17, // @[:@82204.4]
  output        io_out_bits_wstrb_18, // @[:@82204.4]
  output        io_out_bits_wstrb_19, // @[:@82204.4]
  output        io_out_bits_wstrb_20, // @[:@82204.4]
  output        io_out_bits_wstrb_21, // @[:@82204.4]
  output        io_out_bits_wstrb_22, // @[:@82204.4]
  output        io_out_bits_wstrb_23, // @[:@82204.4]
  output        io_out_bits_wstrb_24, // @[:@82204.4]
  output        io_out_bits_wstrb_25, // @[:@82204.4]
  output        io_out_bits_wstrb_26, // @[:@82204.4]
  output        io_out_bits_wstrb_27, // @[:@82204.4]
  output        io_out_bits_wstrb_28, // @[:@82204.4]
  output        io_out_bits_wstrb_29, // @[:@82204.4]
  output        io_out_bits_wstrb_30, // @[:@82204.4]
  output        io_out_bits_wstrb_31, // @[:@82204.4]
  output        io_out_bits_wstrb_32, // @[:@82204.4]
  output        io_out_bits_wstrb_33, // @[:@82204.4]
  output        io_out_bits_wstrb_34, // @[:@82204.4]
  output        io_out_bits_wstrb_35, // @[:@82204.4]
  output        io_out_bits_wstrb_36, // @[:@82204.4]
  output        io_out_bits_wstrb_37, // @[:@82204.4]
  output        io_out_bits_wstrb_38, // @[:@82204.4]
  output        io_out_bits_wstrb_39, // @[:@82204.4]
  output        io_out_bits_wstrb_40, // @[:@82204.4]
  output        io_out_bits_wstrb_41, // @[:@82204.4]
  output        io_out_bits_wstrb_42, // @[:@82204.4]
  output        io_out_bits_wstrb_43, // @[:@82204.4]
  output        io_out_bits_wstrb_44, // @[:@82204.4]
  output        io_out_bits_wstrb_45, // @[:@82204.4]
  output        io_out_bits_wstrb_46, // @[:@82204.4]
  output        io_out_bits_wstrb_47, // @[:@82204.4]
  output        io_out_bits_wstrb_48, // @[:@82204.4]
  output        io_out_bits_wstrb_49, // @[:@82204.4]
  output        io_out_bits_wstrb_50, // @[:@82204.4]
  output        io_out_bits_wstrb_51, // @[:@82204.4]
  output        io_out_bits_wstrb_52, // @[:@82204.4]
  output        io_out_bits_wstrb_53, // @[:@82204.4]
  output        io_out_bits_wstrb_54, // @[:@82204.4]
  output        io_out_bits_wstrb_55, // @[:@82204.4]
  output        io_out_bits_wstrb_56, // @[:@82204.4]
  output        io_out_bits_wstrb_57, // @[:@82204.4]
  output        io_out_bits_wstrb_58, // @[:@82204.4]
  output        io_out_bits_wstrb_59, // @[:@82204.4]
  output        io_out_bits_wstrb_60, // @[:@82204.4]
  output        io_out_bits_wstrb_61, // @[:@82204.4]
  output        io_out_bits_wstrb_62, // @[:@82204.4]
  output        io_out_bits_wstrb_63 // @[:@82204.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@82206.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@82206.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@82291.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@82290.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@82357.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@82358.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@82359.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@82360.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@82361.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@82362.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@82363.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@82364.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@82365.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@82366.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@82367.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@82368.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@82369.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@82370.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@82371.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@82372.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@82293.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@82294.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@82295.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@82296.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@82297.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@82298.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@82299.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@82300.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@82301.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@82302.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@82303.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@82304.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@82305.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@82306.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@82307.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@82308.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@82309.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@82310.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@82311.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@82312.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@82313.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@82314.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@82315.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@82316.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@82317.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@82318.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@82319.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@82320.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@82321.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@82322.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@82323.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@82324.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@82325.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@82326.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@82327.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@82328.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@82329.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@82330.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@82331.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@82332.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@82333.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@82334.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@82335.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@82336.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@82337.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@82338.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@82339.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@82340.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@82341.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@82342.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@82343.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@82344.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@82345.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@82346.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@82347.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@82348.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@82349.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@82350.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@82351.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@82352.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@82353.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@82354.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@82355.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@82356.4]
endmodule
module ElementCounter( // @[:@82374.2]
  input         clock, // @[:@82375.4]
  input         reset, // @[:@82376.4]
  input         io_reset, // @[:@82377.4]
  input         io_enable, // @[:@82377.4]
  output [31:0] io_out // @[:@82377.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@82379.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@82380.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@82381.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@82386.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@82382.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@82380.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@82381.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@82386.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@82382.4]
  assign io_out = count; // @[Counter.scala 47:10:@82389.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@82391.2]
  input         clock, // @[:@82392.4]
  input         reset, // @[:@82393.4]
  output        io_app_0_cmd_ready, // @[:@82394.4]
  input         io_app_0_cmd_valid, // @[:@82394.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@82394.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@82394.4]
  input         io_app_0_cmd_bits_isWr, // @[:@82394.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@82394.4]
  output        io_app_0_wdata_ready, // @[:@82394.4]
  input         io_app_0_wdata_valid, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@82394.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@82394.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@82394.4]
  input         io_app_0_rresp_ready, // @[:@82394.4]
  input         io_app_0_wresp_ready, // @[:@82394.4]
  output        io_app_0_wresp_valid, // @[:@82394.4]
  input         io_dram_cmd_ready, // @[:@82394.4]
  output        io_dram_cmd_valid, // @[:@82394.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@82394.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@82394.4]
  output        io_dram_cmd_bits_isWr, // @[:@82394.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@82394.4]
  input         io_dram_wdata_ready, // @[:@82394.4]
  output        io_dram_wdata_valid, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@82394.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@82394.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@82394.4]
  output        io_dram_rresp_ready, // @[:@82394.4]
  output        io_dram_wresp_ready, // @[:@82394.4]
  input         io_dram_wresp_valid, // @[:@82394.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@82394.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@82623.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@82623.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@82623.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@82623.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@82623.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@82630.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@82630.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@82630.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@82630.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@82630.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@82640.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@82640.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@82640.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@82640.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@82640.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@82640.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@82640.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@82640.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@82640.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@82640.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@82640.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@82640.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@82663.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@82663.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@82666.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@82666.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@82666.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@82666.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@82666.4]
  wire  _T_346; // @[package.scala 96:25:@82635.4 package.scala 96:25:@82636.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@82637.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@82639.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@82655.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@82657.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@82660.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@82669.4]
  wire [31:0] _T_365; // @[:@82673.4 :@82674.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@82675.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@82681.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@82684.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@82685.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@82872.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@82879.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@82884.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@82888.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@82889.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@82913.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@82623.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@82630.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@82640.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@82663.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@82666.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@82635.4 package.scala 96:25:@82636.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@82637.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@82639.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@82655.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@82657.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@82660.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@82669.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@82673.4 :@82674.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@82675.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@82681.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@82684.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@82685.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@82872.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@82879.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@82884.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@82888.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@82889.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@82913.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@82886.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@82892.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@82915.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@82775.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@82774.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@82773.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@82771.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@82770.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@82858.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@82842.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@82843.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@82844.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@82845.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@82846.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@82847.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@82848.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@82849.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@82850.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@82851.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@82852.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@82853.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@82854.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@82855.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@82856.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@82857.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@82778.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@82779.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@82780.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@82781.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@82782.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@82783.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@82784.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@82785.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@82786.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@82787.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@82788.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@82789.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@82790.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@82791.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@82792.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@82793.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@82794.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@82795.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@82796.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@82797.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@82798.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@82799.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@82800.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@82801.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@82802.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@82803.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@82804.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@82805.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@82806.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@82807.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@82808.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@82809.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@82810.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@82811.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@82812.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@82813.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@82814.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@82815.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@82816.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@82817.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@82818.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@82819.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@82820.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@82821.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@82822.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@82823.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@82824.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@82825.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@82826.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@82827.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@82828.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@82829.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@82830.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@82831.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@82832.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@82833.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@82834.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@82835.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@82836.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@82837.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@82838.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@82839.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@82840.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@82841.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@82919.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@82922.4]
  assign RetimeWrapper_clock = clock; // @[:@82624.4]
  assign RetimeWrapper_reset = reset; // @[:@82625.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@82627.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@82626.4]
  assign RetimeWrapper_1_clock = clock; // @[:@82631.4]
  assign RetimeWrapper_1_reset = reset; // @[:@82632.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@82634.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@82633.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@82643.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@82649.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@82648.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@82646.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@82645.4 FringeBundles.scala 115:32:@82662.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@82776.4 StreamArbiter.scala 57:23:@82882.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@82687.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@82754.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@82755.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@82756.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@82757.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@82758.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@82759.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@82760.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@82761.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@82762.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@82763.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@82764.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@82765.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@82766.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@82767.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@82768.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@82769.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@82690.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@82691.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@82692.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@82693.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@82694.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@82695.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@82696.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@82697.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@82698.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@82699.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@82700.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@82701.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@82702.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@82703.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@82704.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@82705.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@82706.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@82707.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@82708.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@82709.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@82710.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@82711.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@82712.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@82713.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@82714.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@82715.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@82716.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@82717.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@82718.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@82719.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@82720.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@82721.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@82722.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@82723.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@82724.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@82725.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@82726.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@82727.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@82728.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@82729.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@82730.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@82731.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@82732.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@82733.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@82734.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@82735.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@82736.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@82737.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@82738.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@82739.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@82740.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@82741.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@82742.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@82743.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@82744.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@82745.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@82746.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@82747.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@82748.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@82749.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@82750.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@82751.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@82752.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@82753.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@82859.4 StreamArbiter.scala 58:25:@82883.4]
  assign elementCtr_clock = clock; // @[:@82667.4]
  assign elementCtr_reset = reset; // @[:@82668.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@82671.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@82670.4]
endmodule
module Counter_72( // @[:@82924.2]
  input         clock, // @[:@82925.4]
  input         reset, // @[:@82926.4]
  input         io_reset, // @[:@82927.4]
  input         io_enable, // @[:@82927.4]
  input  [31:0] io_stride, // @[:@82927.4]
  output [31:0] io_out, // @[:@82927.4]
  output [31:0] io_next // @[:@82927.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@82929.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@82930.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@82931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@82936.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@82932.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@82930.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@82931.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@82936.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@82932.4]
  assign io_out = count; // @[Counter.scala 25:10:@82939.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@82940.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@82942.2]
  input         clock, // @[:@82943.4]
  input         reset, // @[:@82944.4]
  output        io_in_cmd_ready, // @[:@82945.4]
  input         io_in_cmd_valid, // @[:@82945.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@82945.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@82945.4]
  input         io_in_cmd_bits_isWr, // @[:@82945.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@82945.4]
  output        io_in_wdata_ready, // @[:@82945.4]
  input         io_in_wdata_valid, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@82945.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@82945.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@82945.4]
  input         io_in_rresp_ready, // @[:@82945.4]
  input         io_in_wresp_ready, // @[:@82945.4]
  output        io_in_wresp_valid, // @[:@82945.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@82945.4]
  input         io_out_cmd_ready, // @[:@82945.4]
  output        io_out_cmd_valid, // @[:@82945.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@82945.4]
  output [31:0] io_out_cmd_bits_size, // @[:@82945.4]
  output        io_out_cmd_bits_isWr, // @[:@82945.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@82945.4]
  input         io_out_wdata_ready, // @[:@82945.4]
  output        io_out_wdata_valid, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@82945.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@82945.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@82945.4]
  output        io_out_rresp_ready, // @[:@82945.4]
  output        io_out_wresp_ready, // @[:@82945.4]
  input         io_out_wresp_valid, // @[:@82945.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@82945.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@83059.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@83059.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@83059.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@83059.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@83059.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@83059.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@83059.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@83062.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@83063.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@83064.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@83065.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@83068.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@83068.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@83069.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@83069.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@83070.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@83073.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@83080.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@83084.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@83087.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@83090.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@83101.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@83059.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@83062.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@83063.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@83064.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@83065.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@83068.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@83068.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@83069.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@83069.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@83070.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@83073.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@83080.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@83084.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@83087.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@83090.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@83101.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@83058.4 AXIProtocol.scala 38:19:@83092.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@83051.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@82948.4 AXIProtocol.scala 46:21:@83106.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@82947.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@83057.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@83056.4 AXIProtocol.scala 29:24:@83075.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@83055.4 AXIProtocol.scala 25:24:@83067.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@83053.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@83052.4 FringeBundles.scala 115:32:@83089.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@83050.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@83034.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@83035.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@83036.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@83037.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@83038.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@83039.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@83040.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@83041.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@83042.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@83043.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@83044.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@83045.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@83046.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@83047.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@83048.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@83049.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@82970.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@82971.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@82972.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@82973.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@82974.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@82975.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@82976.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@82977.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@82978.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@82979.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@82980.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@82981.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@82982.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@82983.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@82984.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@82985.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@82986.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@82987.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@82988.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@82989.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@82990.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@82991.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@82992.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@82993.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@82994.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@82995.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@82996.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@82997.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@82998.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@82999.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@83000.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@83001.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@83002.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@83003.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@83004.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@83005.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@83006.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@83007.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@83008.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@83009.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@83010.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@83011.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@83012.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@83013.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@83014.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@83015.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@83016.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@83017.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@83018.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@83019.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@83020.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@83021.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@83022.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@83023.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@83024.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@83025.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@83026.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@83027.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@83028.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@83029.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@83030.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@83031.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@83032.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@83033.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@82968.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@82949.4 AXIProtocol.scala 47:22:@83108.4]
  assign cmdSizeCounter_clock = clock; // @[:@83060.4]
  assign cmdSizeCounter_reset = reset; // @[:@83061.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@83093.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@83094.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@83095.4]
endmodule
module AXICmdIssue( // @[:@83128.2]
  input         clock, // @[:@83129.4]
  input         reset, // @[:@83130.4]
  output        io_in_cmd_ready, // @[:@83131.4]
  input         io_in_cmd_valid, // @[:@83131.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@83131.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@83131.4]
  input         io_in_cmd_bits_isWr, // @[:@83131.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@83131.4]
  output        io_in_wdata_ready, // @[:@83131.4]
  input         io_in_wdata_valid, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@83131.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@83131.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@83131.4]
  input         io_in_rresp_ready, // @[:@83131.4]
  input         io_in_wresp_ready, // @[:@83131.4]
  output        io_in_wresp_valid, // @[:@83131.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@83131.4]
  input         io_out_cmd_ready, // @[:@83131.4]
  output        io_out_cmd_valid, // @[:@83131.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@83131.4]
  output [31:0] io_out_cmd_bits_size, // @[:@83131.4]
  output        io_out_cmd_bits_isWr, // @[:@83131.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@83131.4]
  input         io_out_wdata_ready, // @[:@83131.4]
  output        io_out_wdata_valid, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@83131.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@83131.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@83131.4]
  output        io_out_wdata_bits_wlast, // @[:@83131.4]
  output        io_out_rresp_ready, // @[:@83131.4]
  output        io_out_wresp_ready, // @[:@83131.4]
  input         io_out_wresp_valid, // @[:@83131.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@83131.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@83245.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@83245.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@83245.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@83245.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@83245.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@83245.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@83245.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@83248.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@83249.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@83250.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@83251.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@83252.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@83258.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@83259.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@83254.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@83268.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@83269.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@83245.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@83249.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@83250.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@83251.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@83252.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@83258.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@83259.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@83254.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@83268.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@83269.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@83244.4 AXIProtocol.scala 81:19:@83266.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@83237.4 AXIProtocol.scala 82:21:@83267.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@83134.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@83133.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@83243.4 AXIProtocol.scala 84:20:@83271.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@83242.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@83241.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@83239.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@83238.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@83236.4 AXIProtocol.scala 86:22:@83273.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@83220.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@83221.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@83222.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@83223.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@83224.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@83225.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@83226.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@83227.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@83228.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@83229.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@83230.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@83231.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@83232.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@83233.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@83234.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@83235.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@83156.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@83157.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@83158.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@83159.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@83160.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@83161.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@83162.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@83163.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@83164.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@83165.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@83166.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@83167.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@83168.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@83169.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@83170.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@83171.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@83172.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@83173.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@83174.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@83175.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@83176.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@83177.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@83178.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@83179.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@83180.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@83181.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@83182.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@83183.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@83184.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@83185.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@83186.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@83187.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@83188.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@83189.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@83190.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@83191.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@83192.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@83193.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@83194.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@83195.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@83196.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@83197.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@83198.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@83199.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@83200.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@83201.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@83202.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@83203.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@83204.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@83205.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@83206.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@83207.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@83208.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@83209.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@83210.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@83211.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@83212.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@83213.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@83214.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@83215.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@83216.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@83217.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@83218.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@83219.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@83155.4 AXIProtocol.scala 87:27:@83274.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@83154.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@83135.4]
  assign wdataCounter_clock = clock; // @[:@83246.4]
  assign wdataCounter_reset = reset; // @[:@83247.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@83262.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@83263.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@83264.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@83276.2]
  input         clock, // @[:@83277.4]
  input         reset, // @[:@83278.4]
  input         io_enable, // @[:@83279.4]
  output        io_app_stores_0_cmd_ready, // @[:@83279.4]
  input         io_app_stores_0_cmd_valid, // @[:@83279.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@83279.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@83279.4]
  output        io_app_stores_0_data_ready, // @[:@83279.4]
  input         io_app_stores_0_data_valid, // @[:@83279.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@83279.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@83279.4]
  input         io_app_stores_0_wresp_ready, // @[:@83279.4]
  output        io_app_stores_0_wresp_valid, // @[:@83279.4]
  output        io_app_stores_0_wresp_bits, // @[:@83279.4]
  input         io_dram_cmd_ready, // @[:@83279.4]
  output        io_dram_cmd_valid, // @[:@83279.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@83279.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@83279.4]
  output        io_dram_cmd_bits_isWr, // @[:@83279.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@83279.4]
  input         io_dram_wdata_ready, // @[:@83279.4]
  output        io_dram_wdata_valid, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@83279.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@83279.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@83279.4]
  output        io_dram_wdata_bits_wlast, // @[:@83279.4]
  output        io_dram_rresp_ready, // @[:@83279.4]
  output        io_dram_wresp_ready, // @[:@83279.4]
  input         io_dram_wresp_valid, // @[:@83279.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@83279.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@84165.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@84179.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@84407.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@84522.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@84522.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@84165.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@84179.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@84407.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@84522.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@84178.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@84174.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@84169.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@84168.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@84747.4 DRAMArbiter.scala 100:23:@84750.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@84746.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@84745.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@84743.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@84742.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@84740.4 DRAMArbiter.scala 101:25:@84752.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@84724.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@84725.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@84726.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@84727.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@84728.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@84729.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@84730.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@84731.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@84732.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@84733.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@84734.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@84735.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@84736.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@84737.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@84738.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@84739.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@84660.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@84661.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@84662.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@84663.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@84664.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@84665.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@84666.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@84667.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@84668.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@84669.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@84670.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@84671.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@84672.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@84673.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@84674.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@84675.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@84676.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@84677.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@84678.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@84679.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@84680.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@84681.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@84682.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@84683.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@84684.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@84685.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@84686.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@84687.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@84688.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@84689.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@84690.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@84691.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@84692.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@84693.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@84694.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@84695.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@84696.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@84697.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@84698.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@84699.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@84700.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@84701.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@84702.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@84703.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@84704.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@84705.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@84706.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@84707.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@84708.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@84709.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@84710.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@84711.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@84712.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@84713.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@84714.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@84715.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@84716.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@84717.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@84718.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@84719.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@84720.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@84721.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@84722.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@84723.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@84659.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@84658.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@84639.4]
  assign StreamControllerStore_clock = clock; // @[:@84166.4]
  assign StreamControllerStore_reset = reset; // @[:@84167.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@84294.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@84287.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@84184.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@84177.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@84176.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@84175.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@84173.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@84172.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@84171.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@84170.4]
  assign StreamArbiter_clock = clock; // @[:@84180.4]
  assign StreamArbiter_reset = reset; // @[:@84181.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@84405.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@84404.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@84403.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@84401.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@84400.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@84398.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@84382.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@84383.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@84384.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@84385.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@84386.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@84387.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@84388.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@84389.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@84390.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@84391.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@84392.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@84393.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@84394.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@84395.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@84396.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@84397.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@84318.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@84319.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@84320.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@84321.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@84322.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@84323.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@84324.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@84325.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@84326.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@84327.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@84328.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@84329.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@84330.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@84331.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@84332.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@84333.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@84334.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@84335.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@84336.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@84337.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@84338.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@84339.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@84340.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@84341.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@84342.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@84343.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@84344.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@84345.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@84346.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@84347.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@84348.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@84349.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@84350.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@84351.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@84352.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@84353.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@84354.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@84355.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@84356.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@84357.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@84358.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@84359.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@84360.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@84361.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@84362.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@84363.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@84364.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@84365.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@84366.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@84367.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@84368.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@84369.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@84370.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@84371.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@84372.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@84373.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@84374.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@84375.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@84376.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@84377.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@84378.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@84379.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@84380.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@84381.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@84316.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@84297.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@84521.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@84514.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@84411.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@84410.4]
  assign AXICmdSplit_clock = clock; // @[:@84408.4]
  assign AXICmdSplit_reset = reset; // @[:@84409.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@84520.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@84519.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@84518.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@84516.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@84515.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@84513.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@84497.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@84498.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@84499.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@84500.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@84501.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@84502.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@84503.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@84504.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@84505.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@84506.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@84507.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@84508.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@84509.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@84510.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@84511.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@84512.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@84433.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@84434.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@84435.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@84436.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@84437.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@84438.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@84439.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@84440.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@84441.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@84442.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@84443.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@84444.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@84445.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@84446.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@84447.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@84448.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@84449.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@84450.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@84451.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@84452.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@84453.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@84454.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@84455.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@84456.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@84457.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@84458.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@84459.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@84460.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@84461.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@84462.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@84463.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@84464.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@84465.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@84466.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@84467.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@84468.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@84469.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@84470.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@84471.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@84472.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@84473.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@84474.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@84475.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@84476.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@84477.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@84478.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@84479.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@84480.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@84481.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@84482.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@84483.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@84484.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@84485.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@84486.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@84487.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@84488.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@84489.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@84490.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@84491.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@84492.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@84493.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@84494.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@84495.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@84496.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@84431.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@84412.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@84636.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@84629.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@84526.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@84525.4]
  assign AXICmdIssue_clock = clock; // @[:@84523.4]
  assign AXICmdIssue_reset = reset; // @[:@84524.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@84635.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@84634.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@84633.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@84631.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@84630.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@84628.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@84612.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@84613.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@84614.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@84615.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@84616.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@84617.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@84618.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@84619.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@84620.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@84621.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@84622.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@84623.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@84624.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@84625.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@84626.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@84627.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@84548.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@84549.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@84550.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@84551.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@84552.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@84553.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@84554.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@84555.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@84556.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@84557.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@84558.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@84559.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@84560.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@84561.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@84562.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@84563.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@84564.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@84565.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@84566.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@84567.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@84568.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@84569.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@84570.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@84571.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@84572.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@84573.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@84574.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@84575.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@84576.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@84577.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@84578.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@84579.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@84580.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@84581.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@84582.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@84583.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@84584.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@84585.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@84586.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@84587.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@84588.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@84589.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@84590.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@84591.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@84592.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@84593.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@84594.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@84595.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@84596.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@84597.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@84598.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@84599.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@84600.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@84601.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@84602.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@84603.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@84604.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@84605.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@84606.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@84607.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@84608.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@84609.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@84610.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@84611.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@84546.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@84527.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@84748.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@84741.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@84638.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@84637.4]
endmodule
module DRAMArbiter_1( // @[:@98977.2]
  input         clock, // @[:@98978.4]
  input         reset, // @[:@98979.4]
  input         io_enable, // @[:@98980.4]
  input         io_dram_cmd_ready, // @[:@98980.4]
  output        io_dram_cmd_valid, // @[:@98980.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@98980.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@98980.4]
  output        io_dram_cmd_bits_isWr, // @[:@98980.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@98980.4]
  input         io_dram_wdata_ready, // @[:@98980.4]
  output        io_dram_wdata_valid, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@98980.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@98980.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@98980.4]
  output        io_dram_wdata_bits_wlast, // @[:@98980.4]
  output        io_dram_rresp_ready, // @[:@98980.4]
  output        io_dram_wresp_ready, // @[:@98980.4]
  input         io_dram_wresp_valid, // @[:@98980.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@98980.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@99866.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@99880.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@100108.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@100223.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@100223.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@99866.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@99880.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@100108.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@100223.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@100448.4 DRAMArbiter.scala 100:23:@100451.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@100447.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@100446.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@100444.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@100443.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@100441.4 DRAMArbiter.scala 101:25:@100453.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@100425.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@100426.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@100427.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@100428.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@100429.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@100430.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@100431.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@100432.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@100433.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@100434.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@100435.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@100436.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@100437.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@100438.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@100439.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@100440.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@100361.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@100362.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@100363.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@100364.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@100365.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@100366.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@100367.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@100368.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@100369.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@100370.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@100371.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@100372.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@100373.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@100374.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@100375.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@100376.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@100377.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@100378.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@100379.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@100380.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@100381.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@100382.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@100383.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@100384.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@100385.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@100386.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@100387.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@100388.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@100389.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@100390.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@100391.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@100392.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@100393.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@100394.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@100395.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@100396.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@100397.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@100398.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@100399.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@100400.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@100401.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@100402.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@100403.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@100404.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@100405.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@100406.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@100407.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@100408.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@100409.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@100410.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@100411.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@100412.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@100413.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@100414.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@100415.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@100416.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@100417.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@100418.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@100419.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@100420.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@100421.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@100422.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@100423.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@100424.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@100360.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@100359.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@100340.4]
  assign StreamControllerStore_clock = clock; // @[:@99867.4]
  assign StreamControllerStore_reset = reset; // @[:@99868.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@99995.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@99988.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@99885.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@99878.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@99877.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@99876.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@99874.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@99873.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@99872.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@99871.4]
  assign StreamArbiter_clock = clock; // @[:@99881.4]
  assign StreamArbiter_reset = reset; // @[:@99882.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@100106.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@100105.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@100104.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@100102.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@100101.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@100099.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@100083.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@100084.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@100085.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@100086.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@100087.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@100088.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@100089.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@100090.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@100091.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@100092.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@100093.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@100094.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@100095.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@100096.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@100097.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@100098.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@100019.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@100020.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@100021.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@100022.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@100023.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@100024.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@100025.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@100026.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@100027.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@100028.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@100029.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@100030.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@100031.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@100032.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@100033.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@100034.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@100035.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@100036.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@100037.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@100038.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@100039.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@100040.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@100041.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@100042.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@100043.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@100044.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@100045.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@100046.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@100047.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@100048.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@100049.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@100050.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@100051.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@100052.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@100053.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@100054.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@100055.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@100056.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@100057.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@100058.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@100059.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@100060.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@100061.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@100062.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@100063.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@100064.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@100065.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@100066.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@100067.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@100068.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@100069.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@100070.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@100071.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@100072.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@100073.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@100074.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@100075.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@100076.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@100077.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@100078.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@100079.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@100080.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@100081.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@100082.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@100017.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@99998.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@100222.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@100215.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@100112.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@100111.4]
  assign AXICmdSplit_clock = clock; // @[:@100109.4]
  assign AXICmdSplit_reset = reset; // @[:@100110.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@100221.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@100220.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@100219.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@100217.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@100216.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@100214.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@100198.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@100199.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@100200.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@100201.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@100202.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@100203.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@100204.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@100205.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@100206.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@100207.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@100208.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@100209.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@100210.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@100211.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@100212.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@100213.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@100134.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@100135.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@100136.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@100137.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@100138.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@100139.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@100140.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@100141.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@100142.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@100143.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@100144.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@100145.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@100146.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@100147.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@100148.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@100149.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@100150.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@100151.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@100152.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@100153.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@100154.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@100155.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@100156.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@100157.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@100158.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@100159.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@100160.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@100161.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@100162.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@100163.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@100164.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@100165.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@100166.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@100167.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@100168.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@100169.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@100170.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@100171.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@100172.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@100173.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@100174.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@100175.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@100176.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@100177.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@100178.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@100179.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@100180.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@100181.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@100182.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@100183.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@100184.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@100185.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@100186.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@100187.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@100188.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@100189.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@100190.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@100191.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@100192.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@100193.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@100194.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@100195.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@100196.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@100197.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@100132.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@100113.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@100337.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@100330.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@100227.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@100226.4]
  assign AXICmdIssue_clock = clock; // @[:@100224.4]
  assign AXICmdIssue_reset = reset; // @[:@100225.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@100336.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@100335.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@100334.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@100332.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@100331.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@100329.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@100313.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@100314.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@100315.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@100316.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@100317.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@100318.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@100319.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@100320.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@100321.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@100322.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@100323.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@100324.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@100325.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@100326.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@100327.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@100328.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@100249.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@100250.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@100251.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@100252.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@100253.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@100254.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@100255.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@100256.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@100257.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@100258.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@100259.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@100260.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@100261.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@100262.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@100263.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@100264.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@100265.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@100266.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@100267.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@100268.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@100269.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@100270.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@100271.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@100272.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@100273.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@100274.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@100275.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@100276.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@100277.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@100278.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@100279.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@100280.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@100281.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@100282.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@100283.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@100284.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@100285.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@100286.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@100287.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@100288.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@100289.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@100290.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@100291.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@100292.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@100293.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@100294.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@100295.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@100296.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@100297.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@100298.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@100299.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@100300.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@100301.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@100302.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@100303.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@100304.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@100305.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@100306.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@100307.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@100308.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@100309.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@100310.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@100311.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@100312.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@100247.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@100228.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@100449.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@100442.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@100339.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@100338.4]
endmodule
module DRAMHeap( // @[:@131085.2]
  input         io_accel_0_req_valid, // @[:@131088.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@131088.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@131088.4]
  output        io_accel_0_resp_valid, // @[:@131088.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@131088.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@131088.4]
  output        io_host_0_req_valid, // @[:@131088.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@131088.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@131088.4]
  input         io_host_0_resp_valid, // @[:@131088.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@131088.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@131088.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@131095.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@131097.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@131096.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@131092.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@131091.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@131090.4]
endmodule
module RetimeWrapper_719( // @[:@131111.2]
  input         clock, // @[:@131112.4]
  input         reset, // @[:@131113.4]
  input         io_flow, // @[:@131114.4]
  input  [63:0] io_in, // @[:@131114.4]
  output [63:0] io_out // @[:@131114.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@131116.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@131116.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@131116.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@131116.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@131116.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@131116.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@131116.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@131129.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@131128.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@131127.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@131126.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@131125.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@131123.4]
endmodule
module FringeFF( // @[:@131131.2]
  input         clock, // @[:@131132.4]
  input         reset, // @[:@131133.4]
  input  [63:0] io_in, // @[:@131134.4]
  input         io_reset, // @[:@131134.4]
  output [63:0] io_out, // @[:@131134.4]
  input         io_enable // @[:@131134.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@131137.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@131137.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@131137.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@131137.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@131137.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@131142.4 package.scala 96:25:@131143.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@131148.6]
  RetimeWrapper_719 RetimeWrapper ( // @[package.scala 93:22:@131137.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@131142.4 package.scala 96:25:@131143.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@131148.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@131154.4]
  assign RetimeWrapper_clock = clock; // @[:@131138.4]
  assign RetimeWrapper_reset = reset; // @[:@131139.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@131141.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@131140.4]
endmodule
module MuxN( // @[:@159770.2]
  input  [63:0] io_ins_0, // @[:@159773.4]
  input  [63:0] io_ins_1, // @[:@159773.4]
  input  [63:0] io_ins_2, // @[:@159773.4]
  input  [63:0] io_ins_3, // @[:@159773.4]
  input  [63:0] io_ins_4, // @[:@159773.4]
  input  [63:0] io_ins_5, // @[:@159773.4]
  input  [63:0] io_ins_6, // @[:@159773.4]
  input  [63:0] io_ins_7, // @[:@159773.4]
  input  [63:0] io_ins_8, // @[:@159773.4]
  input  [63:0] io_ins_9, // @[:@159773.4]
  input  [63:0] io_ins_10, // @[:@159773.4]
  input  [63:0] io_ins_11, // @[:@159773.4]
  input  [63:0] io_ins_12, // @[:@159773.4]
  input  [63:0] io_ins_13, // @[:@159773.4]
  input  [63:0] io_ins_14, // @[:@159773.4]
  input  [63:0] io_ins_15, // @[:@159773.4]
  input  [63:0] io_ins_16, // @[:@159773.4]
  input  [63:0] io_ins_17, // @[:@159773.4]
  input  [63:0] io_ins_18, // @[:@159773.4]
  input  [63:0] io_ins_19, // @[:@159773.4]
  input  [63:0] io_ins_20, // @[:@159773.4]
  input  [63:0] io_ins_21, // @[:@159773.4]
  input  [63:0] io_ins_22, // @[:@159773.4]
  input  [63:0] io_ins_23, // @[:@159773.4]
  input  [63:0] io_ins_24, // @[:@159773.4]
  input  [63:0] io_ins_25, // @[:@159773.4]
  input  [63:0] io_ins_26, // @[:@159773.4]
  input  [63:0] io_ins_27, // @[:@159773.4]
  input  [63:0] io_ins_28, // @[:@159773.4]
  input  [63:0] io_ins_29, // @[:@159773.4]
  input  [63:0] io_ins_30, // @[:@159773.4]
  input  [63:0] io_ins_31, // @[:@159773.4]
  input  [63:0] io_ins_32, // @[:@159773.4]
  input  [63:0] io_ins_33, // @[:@159773.4]
  input  [63:0] io_ins_34, // @[:@159773.4]
  input  [63:0] io_ins_35, // @[:@159773.4]
  input  [63:0] io_ins_36, // @[:@159773.4]
  input  [63:0] io_ins_37, // @[:@159773.4]
  input  [63:0] io_ins_38, // @[:@159773.4]
  input  [63:0] io_ins_39, // @[:@159773.4]
  input  [63:0] io_ins_40, // @[:@159773.4]
  input  [63:0] io_ins_41, // @[:@159773.4]
  input  [63:0] io_ins_42, // @[:@159773.4]
  input  [63:0] io_ins_43, // @[:@159773.4]
  input  [63:0] io_ins_44, // @[:@159773.4]
  input  [63:0] io_ins_45, // @[:@159773.4]
  input  [63:0] io_ins_46, // @[:@159773.4]
  input  [63:0] io_ins_47, // @[:@159773.4]
  input  [63:0] io_ins_48, // @[:@159773.4]
  input  [63:0] io_ins_49, // @[:@159773.4]
  input  [63:0] io_ins_50, // @[:@159773.4]
  input  [63:0] io_ins_51, // @[:@159773.4]
  input  [63:0] io_ins_52, // @[:@159773.4]
  input  [63:0] io_ins_53, // @[:@159773.4]
  input  [63:0] io_ins_54, // @[:@159773.4]
  input  [63:0] io_ins_55, // @[:@159773.4]
  input  [63:0] io_ins_56, // @[:@159773.4]
  input  [63:0] io_ins_57, // @[:@159773.4]
  input  [63:0] io_ins_58, // @[:@159773.4]
  input  [63:0] io_ins_59, // @[:@159773.4]
  input  [63:0] io_ins_60, // @[:@159773.4]
  input  [63:0] io_ins_61, // @[:@159773.4]
  input  [63:0] io_ins_62, // @[:@159773.4]
  input  [63:0] io_ins_63, // @[:@159773.4]
  input  [63:0] io_ins_64, // @[:@159773.4]
  input  [63:0] io_ins_65, // @[:@159773.4]
  input  [63:0] io_ins_66, // @[:@159773.4]
  input  [63:0] io_ins_67, // @[:@159773.4]
  input  [63:0] io_ins_68, // @[:@159773.4]
  input  [63:0] io_ins_69, // @[:@159773.4]
  input  [63:0] io_ins_70, // @[:@159773.4]
  input  [63:0] io_ins_71, // @[:@159773.4]
  input  [63:0] io_ins_72, // @[:@159773.4]
  input  [63:0] io_ins_73, // @[:@159773.4]
  input  [63:0] io_ins_74, // @[:@159773.4]
  input  [63:0] io_ins_75, // @[:@159773.4]
  input  [63:0] io_ins_76, // @[:@159773.4]
  input  [63:0] io_ins_77, // @[:@159773.4]
  input  [63:0] io_ins_78, // @[:@159773.4]
  input  [63:0] io_ins_79, // @[:@159773.4]
  input  [63:0] io_ins_80, // @[:@159773.4]
  input  [63:0] io_ins_81, // @[:@159773.4]
  input  [63:0] io_ins_82, // @[:@159773.4]
  input  [63:0] io_ins_83, // @[:@159773.4]
  input  [63:0] io_ins_84, // @[:@159773.4]
  input  [63:0] io_ins_85, // @[:@159773.4]
  input  [63:0] io_ins_86, // @[:@159773.4]
  input  [63:0] io_ins_87, // @[:@159773.4]
  input  [63:0] io_ins_88, // @[:@159773.4]
  input  [63:0] io_ins_89, // @[:@159773.4]
  input  [63:0] io_ins_90, // @[:@159773.4]
  input  [63:0] io_ins_91, // @[:@159773.4]
  input  [63:0] io_ins_92, // @[:@159773.4]
  input  [63:0] io_ins_93, // @[:@159773.4]
  input  [63:0] io_ins_94, // @[:@159773.4]
  input  [63:0] io_ins_95, // @[:@159773.4]
  input  [63:0] io_ins_96, // @[:@159773.4]
  input  [63:0] io_ins_97, // @[:@159773.4]
  input  [63:0] io_ins_98, // @[:@159773.4]
  input  [63:0] io_ins_99, // @[:@159773.4]
  input  [63:0] io_ins_100, // @[:@159773.4]
  input  [63:0] io_ins_101, // @[:@159773.4]
  input  [63:0] io_ins_102, // @[:@159773.4]
  input  [63:0] io_ins_103, // @[:@159773.4]
  input  [63:0] io_ins_104, // @[:@159773.4]
  input  [63:0] io_ins_105, // @[:@159773.4]
  input  [63:0] io_ins_106, // @[:@159773.4]
  input  [63:0] io_ins_107, // @[:@159773.4]
  input  [63:0] io_ins_108, // @[:@159773.4]
  input  [63:0] io_ins_109, // @[:@159773.4]
  input  [63:0] io_ins_110, // @[:@159773.4]
  input  [63:0] io_ins_111, // @[:@159773.4]
  input  [63:0] io_ins_112, // @[:@159773.4]
  input  [63:0] io_ins_113, // @[:@159773.4]
  input  [63:0] io_ins_114, // @[:@159773.4]
  input  [63:0] io_ins_115, // @[:@159773.4]
  input  [63:0] io_ins_116, // @[:@159773.4]
  input  [63:0] io_ins_117, // @[:@159773.4]
  input  [63:0] io_ins_118, // @[:@159773.4]
  input  [63:0] io_ins_119, // @[:@159773.4]
  input  [63:0] io_ins_120, // @[:@159773.4]
  input  [63:0] io_ins_121, // @[:@159773.4]
  input  [63:0] io_ins_122, // @[:@159773.4]
  input  [63:0] io_ins_123, // @[:@159773.4]
  input  [63:0] io_ins_124, // @[:@159773.4]
  input  [63:0] io_ins_125, // @[:@159773.4]
  input  [63:0] io_ins_126, // @[:@159773.4]
  input  [63:0] io_ins_127, // @[:@159773.4]
  input  [63:0] io_ins_128, // @[:@159773.4]
  input  [63:0] io_ins_129, // @[:@159773.4]
  input  [63:0] io_ins_130, // @[:@159773.4]
  input  [63:0] io_ins_131, // @[:@159773.4]
  input  [63:0] io_ins_132, // @[:@159773.4]
  input  [63:0] io_ins_133, // @[:@159773.4]
  input  [63:0] io_ins_134, // @[:@159773.4]
  input  [63:0] io_ins_135, // @[:@159773.4]
  input  [63:0] io_ins_136, // @[:@159773.4]
  input  [63:0] io_ins_137, // @[:@159773.4]
  input  [63:0] io_ins_138, // @[:@159773.4]
  input  [63:0] io_ins_139, // @[:@159773.4]
  input  [63:0] io_ins_140, // @[:@159773.4]
  input  [63:0] io_ins_141, // @[:@159773.4]
  input  [63:0] io_ins_142, // @[:@159773.4]
  input  [63:0] io_ins_143, // @[:@159773.4]
  input  [63:0] io_ins_144, // @[:@159773.4]
  input  [63:0] io_ins_145, // @[:@159773.4]
  input  [63:0] io_ins_146, // @[:@159773.4]
  input  [63:0] io_ins_147, // @[:@159773.4]
  input  [63:0] io_ins_148, // @[:@159773.4]
  input  [63:0] io_ins_149, // @[:@159773.4]
  input  [63:0] io_ins_150, // @[:@159773.4]
  input  [63:0] io_ins_151, // @[:@159773.4]
  input  [63:0] io_ins_152, // @[:@159773.4]
  input  [63:0] io_ins_153, // @[:@159773.4]
  input  [63:0] io_ins_154, // @[:@159773.4]
  input  [63:0] io_ins_155, // @[:@159773.4]
  input  [63:0] io_ins_156, // @[:@159773.4]
  input  [63:0] io_ins_157, // @[:@159773.4]
  input  [63:0] io_ins_158, // @[:@159773.4]
  input  [63:0] io_ins_159, // @[:@159773.4]
  input  [63:0] io_ins_160, // @[:@159773.4]
  input  [63:0] io_ins_161, // @[:@159773.4]
  input  [63:0] io_ins_162, // @[:@159773.4]
  input  [63:0] io_ins_163, // @[:@159773.4]
  input  [63:0] io_ins_164, // @[:@159773.4]
  input  [63:0] io_ins_165, // @[:@159773.4]
  input  [63:0] io_ins_166, // @[:@159773.4]
  input  [63:0] io_ins_167, // @[:@159773.4]
  input  [63:0] io_ins_168, // @[:@159773.4]
  input  [63:0] io_ins_169, // @[:@159773.4]
  input  [63:0] io_ins_170, // @[:@159773.4]
  input  [63:0] io_ins_171, // @[:@159773.4]
  input  [63:0] io_ins_172, // @[:@159773.4]
  input  [63:0] io_ins_173, // @[:@159773.4]
  input  [63:0] io_ins_174, // @[:@159773.4]
  input  [63:0] io_ins_175, // @[:@159773.4]
  input  [63:0] io_ins_176, // @[:@159773.4]
  input  [63:0] io_ins_177, // @[:@159773.4]
  input  [63:0] io_ins_178, // @[:@159773.4]
  input  [63:0] io_ins_179, // @[:@159773.4]
  input  [63:0] io_ins_180, // @[:@159773.4]
  input  [63:0] io_ins_181, // @[:@159773.4]
  input  [63:0] io_ins_182, // @[:@159773.4]
  input  [63:0] io_ins_183, // @[:@159773.4]
  input  [63:0] io_ins_184, // @[:@159773.4]
  input  [63:0] io_ins_185, // @[:@159773.4]
  input  [63:0] io_ins_186, // @[:@159773.4]
  input  [63:0] io_ins_187, // @[:@159773.4]
  input  [63:0] io_ins_188, // @[:@159773.4]
  input  [63:0] io_ins_189, // @[:@159773.4]
  input  [63:0] io_ins_190, // @[:@159773.4]
  input  [63:0] io_ins_191, // @[:@159773.4]
  input  [63:0] io_ins_192, // @[:@159773.4]
  input  [63:0] io_ins_193, // @[:@159773.4]
  input  [63:0] io_ins_194, // @[:@159773.4]
  input  [63:0] io_ins_195, // @[:@159773.4]
  input  [63:0] io_ins_196, // @[:@159773.4]
  input  [63:0] io_ins_197, // @[:@159773.4]
  input  [63:0] io_ins_198, // @[:@159773.4]
  input  [63:0] io_ins_199, // @[:@159773.4]
  input  [63:0] io_ins_200, // @[:@159773.4]
  input  [63:0] io_ins_201, // @[:@159773.4]
  input  [63:0] io_ins_202, // @[:@159773.4]
  input  [63:0] io_ins_203, // @[:@159773.4]
  input  [63:0] io_ins_204, // @[:@159773.4]
  input  [63:0] io_ins_205, // @[:@159773.4]
  input  [63:0] io_ins_206, // @[:@159773.4]
  input  [63:0] io_ins_207, // @[:@159773.4]
  input  [63:0] io_ins_208, // @[:@159773.4]
  input  [63:0] io_ins_209, // @[:@159773.4]
  input  [63:0] io_ins_210, // @[:@159773.4]
  input  [63:0] io_ins_211, // @[:@159773.4]
  input  [63:0] io_ins_212, // @[:@159773.4]
  input  [63:0] io_ins_213, // @[:@159773.4]
  input  [63:0] io_ins_214, // @[:@159773.4]
  input  [63:0] io_ins_215, // @[:@159773.4]
  input  [63:0] io_ins_216, // @[:@159773.4]
  input  [63:0] io_ins_217, // @[:@159773.4]
  input  [63:0] io_ins_218, // @[:@159773.4]
  input  [63:0] io_ins_219, // @[:@159773.4]
  input  [63:0] io_ins_220, // @[:@159773.4]
  input  [63:0] io_ins_221, // @[:@159773.4]
  input  [63:0] io_ins_222, // @[:@159773.4]
  input  [63:0] io_ins_223, // @[:@159773.4]
  input  [63:0] io_ins_224, // @[:@159773.4]
  input  [63:0] io_ins_225, // @[:@159773.4]
  input  [63:0] io_ins_226, // @[:@159773.4]
  input  [63:0] io_ins_227, // @[:@159773.4]
  input  [63:0] io_ins_228, // @[:@159773.4]
  input  [63:0] io_ins_229, // @[:@159773.4]
  input  [63:0] io_ins_230, // @[:@159773.4]
  input  [63:0] io_ins_231, // @[:@159773.4]
  input  [63:0] io_ins_232, // @[:@159773.4]
  input  [63:0] io_ins_233, // @[:@159773.4]
  input  [63:0] io_ins_234, // @[:@159773.4]
  input  [63:0] io_ins_235, // @[:@159773.4]
  input  [63:0] io_ins_236, // @[:@159773.4]
  input  [63:0] io_ins_237, // @[:@159773.4]
  input  [63:0] io_ins_238, // @[:@159773.4]
  input  [63:0] io_ins_239, // @[:@159773.4]
  input  [63:0] io_ins_240, // @[:@159773.4]
  input  [63:0] io_ins_241, // @[:@159773.4]
  input  [63:0] io_ins_242, // @[:@159773.4]
  input  [63:0] io_ins_243, // @[:@159773.4]
  input  [63:0] io_ins_244, // @[:@159773.4]
  input  [63:0] io_ins_245, // @[:@159773.4]
  input  [63:0] io_ins_246, // @[:@159773.4]
  input  [63:0] io_ins_247, // @[:@159773.4]
  input  [63:0] io_ins_248, // @[:@159773.4]
  input  [63:0] io_ins_249, // @[:@159773.4]
  input  [63:0] io_ins_250, // @[:@159773.4]
  input  [63:0] io_ins_251, // @[:@159773.4]
  input  [63:0] io_ins_252, // @[:@159773.4]
  input  [63:0] io_ins_253, // @[:@159773.4]
  input  [63:0] io_ins_254, // @[:@159773.4]
  input  [63:0] io_ins_255, // @[:@159773.4]
  input  [63:0] io_ins_256, // @[:@159773.4]
  input  [63:0] io_ins_257, // @[:@159773.4]
  input  [63:0] io_ins_258, // @[:@159773.4]
  input  [63:0] io_ins_259, // @[:@159773.4]
  input  [63:0] io_ins_260, // @[:@159773.4]
  input  [63:0] io_ins_261, // @[:@159773.4]
  input  [63:0] io_ins_262, // @[:@159773.4]
  input  [63:0] io_ins_263, // @[:@159773.4]
  input  [63:0] io_ins_264, // @[:@159773.4]
  input  [63:0] io_ins_265, // @[:@159773.4]
  input  [63:0] io_ins_266, // @[:@159773.4]
  input  [63:0] io_ins_267, // @[:@159773.4]
  input  [63:0] io_ins_268, // @[:@159773.4]
  input  [63:0] io_ins_269, // @[:@159773.4]
  input  [63:0] io_ins_270, // @[:@159773.4]
  input  [63:0] io_ins_271, // @[:@159773.4]
  input  [63:0] io_ins_272, // @[:@159773.4]
  input  [63:0] io_ins_273, // @[:@159773.4]
  input  [63:0] io_ins_274, // @[:@159773.4]
  input  [63:0] io_ins_275, // @[:@159773.4]
  input  [63:0] io_ins_276, // @[:@159773.4]
  input  [63:0] io_ins_277, // @[:@159773.4]
  input  [63:0] io_ins_278, // @[:@159773.4]
  input  [63:0] io_ins_279, // @[:@159773.4]
  input  [63:0] io_ins_280, // @[:@159773.4]
  input  [63:0] io_ins_281, // @[:@159773.4]
  input  [63:0] io_ins_282, // @[:@159773.4]
  input  [63:0] io_ins_283, // @[:@159773.4]
  input  [63:0] io_ins_284, // @[:@159773.4]
  input  [63:0] io_ins_285, // @[:@159773.4]
  input  [63:0] io_ins_286, // @[:@159773.4]
  input  [63:0] io_ins_287, // @[:@159773.4]
  input  [63:0] io_ins_288, // @[:@159773.4]
  input  [63:0] io_ins_289, // @[:@159773.4]
  input  [63:0] io_ins_290, // @[:@159773.4]
  input  [63:0] io_ins_291, // @[:@159773.4]
  input  [63:0] io_ins_292, // @[:@159773.4]
  input  [63:0] io_ins_293, // @[:@159773.4]
  input  [63:0] io_ins_294, // @[:@159773.4]
  input  [63:0] io_ins_295, // @[:@159773.4]
  input  [63:0] io_ins_296, // @[:@159773.4]
  input  [63:0] io_ins_297, // @[:@159773.4]
  input  [63:0] io_ins_298, // @[:@159773.4]
  input  [63:0] io_ins_299, // @[:@159773.4]
  input  [63:0] io_ins_300, // @[:@159773.4]
  input  [63:0] io_ins_301, // @[:@159773.4]
  input  [63:0] io_ins_302, // @[:@159773.4]
  input  [63:0] io_ins_303, // @[:@159773.4]
  input  [63:0] io_ins_304, // @[:@159773.4]
  input  [63:0] io_ins_305, // @[:@159773.4]
  input  [63:0] io_ins_306, // @[:@159773.4]
  input  [63:0] io_ins_307, // @[:@159773.4]
  input  [63:0] io_ins_308, // @[:@159773.4]
  input  [63:0] io_ins_309, // @[:@159773.4]
  input  [63:0] io_ins_310, // @[:@159773.4]
  input  [63:0] io_ins_311, // @[:@159773.4]
  input  [63:0] io_ins_312, // @[:@159773.4]
  input  [63:0] io_ins_313, // @[:@159773.4]
  input  [63:0] io_ins_314, // @[:@159773.4]
  input  [63:0] io_ins_315, // @[:@159773.4]
  input  [63:0] io_ins_316, // @[:@159773.4]
  input  [63:0] io_ins_317, // @[:@159773.4]
  input  [63:0] io_ins_318, // @[:@159773.4]
  input  [63:0] io_ins_319, // @[:@159773.4]
  input  [63:0] io_ins_320, // @[:@159773.4]
  input  [63:0] io_ins_321, // @[:@159773.4]
  input  [63:0] io_ins_322, // @[:@159773.4]
  input  [63:0] io_ins_323, // @[:@159773.4]
  input  [63:0] io_ins_324, // @[:@159773.4]
  input  [63:0] io_ins_325, // @[:@159773.4]
  input  [63:0] io_ins_326, // @[:@159773.4]
  input  [63:0] io_ins_327, // @[:@159773.4]
  input  [63:0] io_ins_328, // @[:@159773.4]
  input  [63:0] io_ins_329, // @[:@159773.4]
  input  [63:0] io_ins_330, // @[:@159773.4]
  input  [63:0] io_ins_331, // @[:@159773.4]
  input  [63:0] io_ins_332, // @[:@159773.4]
  input  [63:0] io_ins_333, // @[:@159773.4]
  input  [63:0] io_ins_334, // @[:@159773.4]
  input  [63:0] io_ins_335, // @[:@159773.4]
  input  [63:0] io_ins_336, // @[:@159773.4]
  input  [63:0] io_ins_337, // @[:@159773.4]
  input  [63:0] io_ins_338, // @[:@159773.4]
  input  [63:0] io_ins_339, // @[:@159773.4]
  input  [63:0] io_ins_340, // @[:@159773.4]
  input  [63:0] io_ins_341, // @[:@159773.4]
  input  [63:0] io_ins_342, // @[:@159773.4]
  input  [63:0] io_ins_343, // @[:@159773.4]
  input  [63:0] io_ins_344, // @[:@159773.4]
  input  [63:0] io_ins_345, // @[:@159773.4]
  input  [63:0] io_ins_346, // @[:@159773.4]
  input  [63:0] io_ins_347, // @[:@159773.4]
  input  [63:0] io_ins_348, // @[:@159773.4]
  input  [63:0] io_ins_349, // @[:@159773.4]
  input  [63:0] io_ins_350, // @[:@159773.4]
  input  [63:0] io_ins_351, // @[:@159773.4]
  input  [63:0] io_ins_352, // @[:@159773.4]
  input  [63:0] io_ins_353, // @[:@159773.4]
  input  [63:0] io_ins_354, // @[:@159773.4]
  input  [63:0] io_ins_355, // @[:@159773.4]
  input  [63:0] io_ins_356, // @[:@159773.4]
  input  [63:0] io_ins_357, // @[:@159773.4]
  input  [63:0] io_ins_358, // @[:@159773.4]
  input  [63:0] io_ins_359, // @[:@159773.4]
  input  [63:0] io_ins_360, // @[:@159773.4]
  input  [63:0] io_ins_361, // @[:@159773.4]
  input  [63:0] io_ins_362, // @[:@159773.4]
  input  [63:0] io_ins_363, // @[:@159773.4]
  input  [63:0] io_ins_364, // @[:@159773.4]
  input  [63:0] io_ins_365, // @[:@159773.4]
  input  [63:0] io_ins_366, // @[:@159773.4]
  input  [63:0] io_ins_367, // @[:@159773.4]
  input  [63:0] io_ins_368, // @[:@159773.4]
  input  [63:0] io_ins_369, // @[:@159773.4]
  input  [63:0] io_ins_370, // @[:@159773.4]
  input  [63:0] io_ins_371, // @[:@159773.4]
  input  [63:0] io_ins_372, // @[:@159773.4]
  input  [63:0] io_ins_373, // @[:@159773.4]
  input  [63:0] io_ins_374, // @[:@159773.4]
  input  [63:0] io_ins_375, // @[:@159773.4]
  input  [63:0] io_ins_376, // @[:@159773.4]
  input  [63:0] io_ins_377, // @[:@159773.4]
  input  [63:0] io_ins_378, // @[:@159773.4]
  input  [63:0] io_ins_379, // @[:@159773.4]
  input  [63:0] io_ins_380, // @[:@159773.4]
  input  [63:0] io_ins_381, // @[:@159773.4]
  input  [63:0] io_ins_382, // @[:@159773.4]
  input  [63:0] io_ins_383, // @[:@159773.4]
  input  [63:0] io_ins_384, // @[:@159773.4]
  input  [63:0] io_ins_385, // @[:@159773.4]
  input  [63:0] io_ins_386, // @[:@159773.4]
  input  [63:0] io_ins_387, // @[:@159773.4]
  input  [63:0] io_ins_388, // @[:@159773.4]
  input  [63:0] io_ins_389, // @[:@159773.4]
  input  [63:0] io_ins_390, // @[:@159773.4]
  input  [63:0] io_ins_391, // @[:@159773.4]
  input  [63:0] io_ins_392, // @[:@159773.4]
  input  [63:0] io_ins_393, // @[:@159773.4]
  input  [63:0] io_ins_394, // @[:@159773.4]
  input  [63:0] io_ins_395, // @[:@159773.4]
  input  [63:0] io_ins_396, // @[:@159773.4]
  input  [63:0] io_ins_397, // @[:@159773.4]
  input  [63:0] io_ins_398, // @[:@159773.4]
  input  [63:0] io_ins_399, // @[:@159773.4]
  input  [63:0] io_ins_400, // @[:@159773.4]
  input  [63:0] io_ins_401, // @[:@159773.4]
  input  [63:0] io_ins_402, // @[:@159773.4]
  input  [63:0] io_ins_403, // @[:@159773.4]
  input  [63:0] io_ins_404, // @[:@159773.4]
  input  [63:0] io_ins_405, // @[:@159773.4]
  input  [63:0] io_ins_406, // @[:@159773.4]
  input  [63:0] io_ins_407, // @[:@159773.4]
  input  [63:0] io_ins_408, // @[:@159773.4]
  input  [63:0] io_ins_409, // @[:@159773.4]
  input  [63:0] io_ins_410, // @[:@159773.4]
  input  [63:0] io_ins_411, // @[:@159773.4]
  input  [63:0] io_ins_412, // @[:@159773.4]
  input  [63:0] io_ins_413, // @[:@159773.4]
  input  [63:0] io_ins_414, // @[:@159773.4]
  input  [63:0] io_ins_415, // @[:@159773.4]
  input  [63:0] io_ins_416, // @[:@159773.4]
  input  [63:0] io_ins_417, // @[:@159773.4]
  input  [63:0] io_ins_418, // @[:@159773.4]
  input  [63:0] io_ins_419, // @[:@159773.4]
  input  [63:0] io_ins_420, // @[:@159773.4]
  input  [63:0] io_ins_421, // @[:@159773.4]
  input  [63:0] io_ins_422, // @[:@159773.4]
  input  [63:0] io_ins_423, // @[:@159773.4]
  input  [63:0] io_ins_424, // @[:@159773.4]
  input  [63:0] io_ins_425, // @[:@159773.4]
  input  [63:0] io_ins_426, // @[:@159773.4]
  input  [63:0] io_ins_427, // @[:@159773.4]
  input  [63:0] io_ins_428, // @[:@159773.4]
  input  [63:0] io_ins_429, // @[:@159773.4]
  input  [63:0] io_ins_430, // @[:@159773.4]
  input  [63:0] io_ins_431, // @[:@159773.4]
  input  [63:0] io_ins_432, // @[:@159773.4]
  input  [63:0] io_ins_433, // @[:@159773.4]
  input  [63:0] io_ins_434, // @[:@159773.4]
  input  [63:0] io_ins_435, // @[:@159773.4]
  input  [63:0] io_ins_436, // @[:@159773.4]
  input  [63:0] io_ins_437, // @[:@159773.4]
  input  [63:0] io_ins_438, // @[:@159773.4]
  input  [63:0] io_ins_439, // @[:@159773.4]
  input  [63:0] io_ins_440, // @[:@159773.4]
  input  [63:0] io_ins_441, // @[:@159773.4]
  input  [63:0] io_ins_442, // @[:@159773.4]
  input  [63:0] io_ins_443, // @[:@159773.4]
  input  [63:0] io_ins_444, // @[:@159773.4]
  input  [63:0] io_ins_445, // @[:@159773.4]
  input  [63:0] io_ins_446, // @[:@159773.4]
  input  [63:0] io_ins_447, // @[:@159773.4]
  input  [63:0] io_ins_448, // @[:@159773.4]
  input  [63:0] io_ins_449, // @[:@159773.4]
  input  [63:0] io_ins_450, // @[:@159773.4]
  input  [63:0] io_ins_451, // @[:@159773.4]
  input  [63:0] io_ins_452, // @[:@159773.4]
  input  [63:0] io_ins_453, // @[:@159773.4]
  input  [63:0] io_ins_454, // @[:@159773.4]
  input  [63:0] io_ins_455, // @[:@159773.4]
  input  [63:0] io_ins_456, // @[:@159773.4]
  input  [63:0] io_ins_457, // @[:@159773.4]
  input  [63:0] io_ins_458, // @[:@159773.4]
  input  [63:0] io_ins_459, // @[:@159773.4]
  input  [63:0] io_ins_460, // @[:@159773.4]
  input  [63:0] io_ins_461, // @[:@159773.4]
  input  [63:0] io_ins_462, // @[:@159773.4]
  input  [63:0] io_ins_463, // @[:@159773.4]
  input  [63:0] io_ins_464, // @[:@159773.4]
  input  [63:0] io_ins_465, // @[:@159773.4]
  input  [63:0] io_ins_466, // @[:@159773.4]
  input  [63:0] io_ins_467, // @[:@159773.4]
  input  [63:0] io_ins_468, // @[:@159773.4]
  input  [63:0] io_ins_469, // @[:@159773.4]
  input  [63:0] io_ins_470, // @[:@159773.4]
  input  [63:0] io_ins_471, // @[:@159773.4]
  input  [63:0] io_ins_472, // @[:@159773.4]
  input  [63:0] io_ins_473, // @[:@159773.4]
  input  [63:0] io_ins_474, // @[:@159773.4]
  input  [63:0] io_ins_475, // @[:@159773.4]
  input  [63:0] io_ins_476, // @[:@159773.4]
  input  [63:0] io_ins_477, // @[:@159773.4]
  input  [63:0] io_ins_478, // @[:@159773.4]
  input  [63:0] io_ins_479, // @[:@159773.4]
  input  [63:0] io_ins_480, // @[:@159773.4]
  input  [63:0] io_ins_481, // @[:@159773.4]
  input  [63:0] io_ins_482, // @[:@159773.4]
  input  [63:0] io_ins_483, // @[:@159773.4]
  input  [63:0] io_ins_484, // @[:@159773.4]
  input  [63:0] io_ins_485, // @[:@159773.4]
  input  [63:0] io_ins_486, // @[:@159773.4]
  input  [63:0] io_ins_487, // @[:@159773.4]
  input  [63:0] io_ins_488, // @[:@159773.4]
  input  [63:0] io_ins_489, // @[:@159773.4]
  input  [63:0] io_ins_490, // @[:@159773.4]
  input  [63:0] io_ins_491, // @[:@159773.4]
  input  [63:0] io_ins_492, // @[:@159773.4]
  input  [63:0] io_ins_493, // @[:@159773.4]
  input  [63:0] io_ins_494, // @[:@159773.4]
  input  [63:0] io_ins_495, // @[:@159773.4]
  input  [63:0] io_ins_496, // @[:@159773.4]
  input  [63:0] io_ins_497, // @[:@159773.4]
  input  [63:0] io_ins_498, // @[:@159773.4]
  input  [63:0] io_ins_499, // @[:@159773.4]
  input  [63:0] io_ins_500, // @[:@159773.4]
  input  [63:0] io_ins_501, // @[:@159773.4]
  input  [63:0] io_ins_502, // @[:@159773.4]
  input  [8:0]  io_sel, // @[:@159773.4]
  output [63:0] io_out // @[:@159773.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@159775.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@159775.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@159775.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@159775.4]
endmodule
module RegFile( // @[:@159777.2]
  input         clock, // @[:@159778.4]
  input         reset, // @[:@159779.4]
  input  [31:0] io_raddr, // @[:@159780.4]
  input         io_wen, // @[:@159780.4]
  input  [31:0] io_waddr, // @[:@159780.4]
  input  [63:0] io_wdata, // @[:@159780.4]
  output [63:0] io_rdata, // @[:@159780.4]
  input         io_reset, // @[:@159780.4]
  output [63:0] io_argIns_0, // @[:@159780.4]
  output [63:0] io_argIns_1, // @[:@159780.4]
  output [63:0] io_argIns_2, // @[:@159780.4]
  output [63:0] io_argIns_3, // @[:@159780.4]
  input         io_argOuts_0_valid, // @[:@159780.4]
  input  [63:0] io_argOuts_0_bits, // @[:@159780.4]
  input         io_argOuts_1_valid, // @[:@159780.4]
  input  [63:0] io_argOuts_1_bits // @[:@159780.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@161790.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@161790.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@161790.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@161790.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@161790.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@161790.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@161802.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@161802.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@161802.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@161802.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@161802.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@161802.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@161821.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@161821.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@161821.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@161821.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@161821.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@161821.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@161833.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@161833.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@161833.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@161833.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@161833.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@161833.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@161845.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@161845.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@161845.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@161845.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@161845.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@161845.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@161859.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@161859.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@161859.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@161859.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@161859.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@161859.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@161873.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@161873.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@161873.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@161873.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@161873.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@161873.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@161887.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@161887.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@161887.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@161887.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@161887.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@161887.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@161901.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@161901.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@161901.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@161901.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@161901.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@161901.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@161915.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@161915.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@161915.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@161915.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@161915.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@161915.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@161929.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@161929.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@161929.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@161929.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@161929.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@161929.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@161943.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@161943.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@161943.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@161943.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@161943.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@161943.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@161957.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@161957.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@161957.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@161957.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@161957.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@161957.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@161971.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@161971.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@161971.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@161971.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@161971.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@161971.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@161985.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@161985.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@161985.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@161985.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@161985.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@161985.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@161999.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@161999.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@161999.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@161999.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@161999.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@161999.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@162013.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@162013.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@162013.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@162013.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@162013.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@162013.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@162027.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@162027.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@162027.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@162027.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@162027.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@162027.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@162041.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@162041.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@162041.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@162041.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@162041.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@162041.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@162055.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@162055.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@162055.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@162055.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@162055.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@162055.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@162069.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@162069.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@162069.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@162069.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@162069.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@162069.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@162083.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@162083.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@162083.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@162083.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@162083.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@162083.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@162097.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@162097.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@162097.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@162097.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@162097.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@162097.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@162111.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@162111.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@162111.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@162111.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@162111.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@162111.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@162125.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@162125.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@162125.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@162125.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@162125.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@162125.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@162139.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@162139.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@162139.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@162139.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@162139.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@162139.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@162153.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@162153.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@162153.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@162153.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@162153.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@162153.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@162167.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@162167.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@162167.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@162167.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@162167.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@162167.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@162181.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@162181.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@162181.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@162181.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@162181.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@162181.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@162195.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@162195.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@162195.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@162195.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@162195.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@162195.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@162209.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@162209.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@162209.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@162209.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@162209.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@162209.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@162223.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@162223.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@162223.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@162223.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@162223.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@162223.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@162237.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@162237.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@162237.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@162237.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@162237.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@162237.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@162251.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@162251.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@162251.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@162251.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@162251.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@162251.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@162265.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@162265.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@162265.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@162265.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@162265.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@162265.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@162279.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@162279.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@162279.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@162279.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@162279.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@162279.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@162293.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@162293.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@162293.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@162293.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@162293.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@162293.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@162307.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@162307.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@162307.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@162307.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@162307.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@162307.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@162321.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@162321.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@162321.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@162321.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@162321.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@162321.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@162335.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@162335.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@162335.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@162335.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@162335.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@162335.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@162349.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@162349.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@162349.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@162349.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@162349.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@162349.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@162363.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@162363.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@162363.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@162363.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@162363.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@162363.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@162377.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@162377.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@162377.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@162377.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@162377.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@162377.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@162391.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@162391.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@162391.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@162391.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@162391.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@162391.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@162405.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@162405.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@162405.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@162405.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@162405.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@162405.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@162419.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@162419.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@162419.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@162419.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@162419.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@162419.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@162433.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@162433.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@162433.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@162433.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@162433.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@162433.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@162447.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@162447.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@162447.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@162447.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@162447.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@162447.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@162461.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@162461.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@162461.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@162461.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@162461.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@162461.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@162475.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@162475.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@162475.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@162475.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@162475.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@162475.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@162489.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@162489.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@162489.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@162489.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@162489.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@162489.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@162503.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@162503.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@162503.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@162503.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@162503.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@162503.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@162517.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@162517.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@162517.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@162517.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@162517.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@162517.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@162531.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@162531.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@162531.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@162531.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@162531.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@162531.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@162545.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@162545.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@162545.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@162545.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@162545.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@162545.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@162559.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@162559.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@162559.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@162559.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@162559.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@162559.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@162573.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@162573.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@162573.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@162573.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@162573.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@162573.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@162587.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@162587.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@162587.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@162587.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@162587.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@162587.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@162601.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@162601.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@162601.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@162601.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@162601.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@162601.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@162615.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@162615.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@162615.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@162615.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@162615.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@162615.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@162629.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@162629.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@162629.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@162629.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@162629.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@162629.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@162643.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@162643.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@162643.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@162643.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@162643.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@162643.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@162657.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@162657.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@162657.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@162657.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@162657.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@162657.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@162671.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@162671.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@162671.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@162671.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@162671.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@162671.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@162685.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@162685.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@162685.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@162685.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@162685.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@162685.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@162699.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@162699.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@162699.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@162699.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@162699.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@162699.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@162713.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@162713.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@162713.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@162713.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@162713.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@162713.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@162727.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@162727.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@162727.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@162727.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@162727.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@162727.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@162741.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@162741.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@162741.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@162741.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@162741.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@162741.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@162755.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@162755.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@162755.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@162755.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@162755.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@162755.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@162769.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@162769.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@162769.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@162769.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@162769.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@162769.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@162783.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@162783.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@162783.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@162783.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@162783.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@162783.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@162797.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@162797.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@162797.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@162797.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@162797.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@162797.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@162811.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@162811.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@162811.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@162811.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@162811.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@162811.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@162825.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@162825.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@162825.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@162825.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@162825.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@162825.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@162839.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@162839.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@162839.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@162839.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@162839.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@162839.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@162853.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@162853.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@162853.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@162853.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@162853.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@162853.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@162867.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@162867.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@162867.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@162867.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@162867.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@162867.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@162881.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@162881.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@162881.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@162881.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@162881.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@162881.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@162895.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@162895.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@162895.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@162895.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@162895.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@162895.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@162909.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@162909.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@162909.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@162909.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@162909.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@162909.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@162923.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@162923.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@162923.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@162923.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@162923.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@162923.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@162937.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@162937.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@162937.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@162937.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@162937.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@162937.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@162951.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@162951.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@162951.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@162951.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@162951.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@162951.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@162965.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@162965.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@162965.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@162965.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@162965.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@162965.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@162979.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@162979.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@162979.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@162979.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@162979.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@162979.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@162993.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@162993.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@162993.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@162993.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@162993.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@162993.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@163007.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@163007.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@163007.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@163007.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@163007.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@163007.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@163021.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@163021.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@163021.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@163021.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@163021.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@163021.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@163035.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@163035.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@163035.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@163035.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@163035.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@163035.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@163049.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@163049.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@163049.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@163049.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@163049.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@163049.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@163063.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@163063.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@163063.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@163063.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@163063.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@163063.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@163077.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@163077.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@163077.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@163077.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@163077.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@163077.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@163091.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@163091.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@163091.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@163091.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@163091.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@163091.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@163105.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@163105.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@163105.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@163105.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@163105.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@163105.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@163119.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@163119.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@163119.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@163119.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@163119.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@163119.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@163133.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@163133.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@163133.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@163133.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@163133.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@163133.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@163147.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@163147.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@163147.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@163147.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@163147.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@163147.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@163161.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@163161.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@163161.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@163161.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@163161.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@163161.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@163175.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@163175.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@163175.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@163175.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@163175.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@163175.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@163189.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@163189.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@163189.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@163189.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@163189.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@163189.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@163203.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@163203.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@163203.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@163203.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@163203.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@163203.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@163217.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@163217.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@163217.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@163217.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@163217.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@163217.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@163231.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@163231.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@163231.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@163231.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@163231.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@163231.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@163245.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@163245.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@163245.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@163245.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@163245.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@163245.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@163259.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@163259.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@163259.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@163259.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@163259.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@163259.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@163273.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@163273.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@163273.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@163273.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@163273.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@163273.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@163287.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@163287.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@163287.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@163287.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@163287.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@163287.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@163301.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@163301.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@163301.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@163301.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@163301.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@163301.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@163315.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@163315.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@163315.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@163315.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@163315.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@163315.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@163329.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@163329.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@163329.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@163329.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@163329.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@163329.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@163343.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@163343.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@163343.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@163343.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@163343.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@163343.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@163357.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@163357.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@163357.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@163357.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@163357.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@163357.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@163371.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@163371.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@163371.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@163371.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@163371.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@163371.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@163385.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@163385.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@163385.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@163385.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@163385.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@163385.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@163399.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@163399.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@163399.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@163399.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@163399.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@163399.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@163413.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@163413.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@163413.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@163413.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@163413.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@163413.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@163427.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@163427.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@163427.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@163427.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@163427.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@163427.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@163441.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@163441.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@163441.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@163441.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@163441.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@163441.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@163455.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@163455.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@163455.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@163455.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@163455.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@163455.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@163469.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@163469.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@163469.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@163469.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@163469.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@163469.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@163483.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@163483.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@163483.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@163483.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@163483.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@163483.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@163497.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@163497.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@163497.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@163497.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@163497.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@163497.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@163511.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@163511.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@163511.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@163511.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@163511.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@163511.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@163525.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@163525.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@163525.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@163525.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@163525.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@163525.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@163539.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@163539.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@163539.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@163539.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@163539.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@163539.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@163553.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@163553.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@163553.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@163553.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@163553.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@163553.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@163567.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@163567.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@163567.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@163567.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@163567.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@163567.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@163581.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@163581.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@163581.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@163581.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@163581.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@163581.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@163595.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@163595.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@163595.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@163595.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@163595.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@163595.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@163609.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@163609.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@163609.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@163609.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@163609.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@163609.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@163623.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@163623.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@163623.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@163623.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@163623.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@163623.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@163637.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@163637.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@163637.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@163637.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@163637.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@163637.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@163651.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@163651.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@163651.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@163651.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@163651.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@163651.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@163665.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@163665.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@163665.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@163665.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@163665.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@163665.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@163679.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@163679.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@163679.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@163679.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@163679.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@163679.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@163693.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@163693.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@163693.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@163693.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@163693.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@163693.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@163707.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@163707.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@163707.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@163707.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@163707.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@163707.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@163721.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@163721.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@163721.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@163721.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@163721.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@163721.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@163735.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@163735.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@163735.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@163735.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@163735.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@163735.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@163749.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@163749.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@163749.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@163749.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@163749.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@163749.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@163763.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@163763.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@163763.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@163763.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@163763.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@163763.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@163777.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@163777.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@163777.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@163777.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@163777.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@163777.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@163791.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@163791.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@163791.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@163791.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@163791.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@163791.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@163805.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@163805.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@163805.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@163805.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@163805.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@163805.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@163819.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@163819.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@163819.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@163819.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@163819.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@163819.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@163833.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@163833.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@163833.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@163833.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@163833.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@163833.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@163847.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@163847.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@163847.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@163847.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@163847.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@163847.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@163861.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@163861.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@163861.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@163861.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@163861.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@163861.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@163875.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@163875.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@163875.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@163875.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@163875.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@163875.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@163889.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@163889.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@163889.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@163889.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@163889.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@163889.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@163903.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@163903.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@163903.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@163903.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@163903.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@163903.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@163917.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@163917.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@163917.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@163917.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@163917.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@163917.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@163931.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@163931.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@163931.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@163931.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@163931.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@163931.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@163945.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@163945.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@163945.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@163945.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@163945.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@163945.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@163959.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@163959.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@163959.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@163959.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@163959.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@163959.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@163973.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@163973.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@163973.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@163973.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@163973.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@163973.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@163987.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@163987.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@163987.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@163987.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@163987.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@163987.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@164001.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@164001.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@164001.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@164001.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@164001.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@164001.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@164015.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@164015.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@164015.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@164015.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@164015.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@164015.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@164029.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@164029.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@164029.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@164029.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@164029.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@164029.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@164043.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@164043.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@164043.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@164043.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@164043.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@164043.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@164057.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@164057.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@164057.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@164057.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@164057.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@164057.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@164071.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@164071.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@164071.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@164071.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@164071.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@164071.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@164085.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@164085.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@164085.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@164085.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@164085.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@164085.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@164099.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@164099.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@164099.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@164099.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@164099.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@164099.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@164113.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@164113.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@164113.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@164113.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@164113.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@164113.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@164127.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@164127.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@164127.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@164127.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@164127.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@164127.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@164141.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@164141.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@164141.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@164141.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@164141.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@164141.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@164155.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@164155.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@164155.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@164155.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@164155.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@164155.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@164169.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@164169.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@164169.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@164169.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@164169.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@164169.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@164183.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@164183.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@164183.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@164183.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@164183.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@164183.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@164197.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@164197.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@164197.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@164197.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@164197.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@164197.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@164211.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@164211.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@164211.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@164211.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@164211.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@164211.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@164225.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@164225.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@164225.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@164225.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@164225.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@164225.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@164239.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@164239.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@164239.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@164239.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@164239.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@164239.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@164253.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@164253.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@164253.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@164253.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@164253.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@164253.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@164267.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@164267.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@164267.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@164267.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@164267.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@164267.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@164281.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@164281.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@164281.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@164281.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@164281.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@164281.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@164295.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@164295.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@164295.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@164295.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@164295.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@164295.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@164309.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@164309.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@164309.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@164309.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@164309.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@164309.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@164323.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@164323.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@164323.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@164323.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@164323.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@164323.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@164337.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@164337.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@164337.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@164337.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@164337.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@164337.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@164351.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@164351.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@164351.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@164351.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@164351.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@164351.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@164365.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@164365.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@164365.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@164365.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@164365.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@164365.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@164379.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@164379.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@164379.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@164379.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@164379.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@164379.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@164393.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@164393.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@164393.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@164393.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@164393.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@164393.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@164407.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@164407.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@164407.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@164407.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@164407.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@164407.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@164421.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@164421.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@164421.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@164421.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@164421.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@164421.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@164435.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@164435.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@164435.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@164435.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@164435.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@164435.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@164449.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@164449.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@164449.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@164449.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@164449.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@164449.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@164463.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@164463.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@164463.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@164463.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@164463.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@164463.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@164477.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@164477.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@164477.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@164477.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@164477.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@164477.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@164491.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@164491.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@164491.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@164491.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@164491.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@164491.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@164505.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@164505.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@164505.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@164505.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@164505.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@164505.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@164519.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@164519.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@164519.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@164519.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@164519.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@164519.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@164533.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@164533.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@164533.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@164533.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@164533.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@164533.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@164547.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@164547.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@164547.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@164547.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@164547.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@164547.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@164561.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@164561.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@164561.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@164561.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@164561.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@164561.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@164575.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@164575.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@164575.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@164575.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@164575.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@164575.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@164589.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@164589.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@164589.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@164589.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@164589.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@164589.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@164603.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@164603.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@164603.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@164603.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@164603.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@164603.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@164617.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@164617.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@164617.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@164617.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@164617.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@164617.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@164631.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@164631.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@164631.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@164631.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@164631.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@164631.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@164645.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@164645.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@164645.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@164645.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@164645.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@164645.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@164659.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@164659.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@164659.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@164659.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@164659.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@164659.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@164673.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@164673.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@164673.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@164673.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@164673.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@164673.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@164687.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@164687.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@164687.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@164687.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@164687.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@164687.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@164701.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@164701.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@164701.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@164701.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@164701.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@164701.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@164715.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@164715.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@164715.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@164715.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@164715.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@164715.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@164729.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@164729.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@164729.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@164729.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@164729.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@164729.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@164743.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@164743.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@164743.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@164743.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@164743.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@164743.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@164757.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@164757.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@164757.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@164757.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@164757.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@164757.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@164771.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@164771.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@164771.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@164771.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@164771.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@164771.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@164785.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@164785.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@164785.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@164785.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@164785.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@164785.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@164799.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@164799.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@164799.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@164799.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@164799.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@164799.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@164813.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@164813.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@164813.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@164813.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@164813.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@164813.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@164827.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@164827.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@164827.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@164827.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@164827.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@164827.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@164841.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@164841.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@164841.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@164841.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@164841.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@164841.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@164855.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@164855.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@164855.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@164855.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@164855.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@164855.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@164869.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@164869.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@164869.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@164869.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@164869.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@164869.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@164883.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@164883.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@164883.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@164883.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@164883.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@164883.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@164897.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@164897.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@164897.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@164897.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@164897.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@164897.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@164911.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@164911.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@164911.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@164911.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@164911.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@164911.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@164925.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@164925.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@164925.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@164925.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@164925.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@164925.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@164939.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@164939.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@164939.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@164939.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@164939.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@164939.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@164953.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@164953.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@164953.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@164953.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@164953.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@164953.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@164967.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@164967.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@164967.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@164967.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@164967.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@164967.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@164981.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@164981.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@164981.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@164981.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@164981.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@164981.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@164995.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@164995.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@164995.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@164995.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@164995.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@164995.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@165009.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@165009.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@165009.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@165009.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@165009.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@165009.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@165023.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@165023.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@165023.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@165023.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@165023.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@165023.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@165037.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@165037.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@165037.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@165037.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@165037.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@165037.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@165051.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@165051.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@165051.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@165051.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@165051.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@165051.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@165065.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@165065.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@165065.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@165065.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@165065.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@165065.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@165079.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@165079.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@165079.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@165079.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@165079.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@165079.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@165093.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@165093.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@165093.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@165093.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@165093.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@165093.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@165107.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@165107.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@165107.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@165107.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@165107.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@165107.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@165121.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@165121.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@165121.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@165121.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@165121.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@165121.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@165135.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@165135.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@165135.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@165135.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@165135.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@165135.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@165149.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@165149.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@165149.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@165149.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@165149.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@165149.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@165163.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@165163.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@165163.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@165163.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@165163.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@165163.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@165177.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@165177.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@165177.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@165177.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@165177.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@165177.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@165191.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@165191.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@165191.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@165191.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@165191.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@165191.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@165205.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@165205.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@165205.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@165205.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@165205.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@165205.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@165219.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@165219.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@165219.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@165219.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@165219.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@165219.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@165233.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@165233.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@165233.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@165233.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@165233.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@165233.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@165247.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@165247.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@165247.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@165247.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@165247.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@165247.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@165261.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@165261.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@165261.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@165261.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@165261.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@165261.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@165275.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@165275.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@165275.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@165275.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@165275.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@165275.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@165289.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@165289.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@165289.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@165289.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@165289.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@165289.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@165303.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@165303.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@165303.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@165303.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@165303.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@165303.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@165317.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@165317.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@165317.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@165317.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@165317.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@165317.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@165331.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@165331.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@165331.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@165331.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@165331.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@165331.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@165345.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@165345.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@165345.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@165345.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@165345.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@165345.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@165359.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@165359.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@165359.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@165359.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@165359.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@165359.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@165373.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@165373.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@165373.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@165373.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@165373.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@165373.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@165387.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@165387.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@165387.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@165387.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@165387.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@165387.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@165401.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@165401.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@165401.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@165401.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@165401.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@165401.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@165415.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@165415.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@165415.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@165415.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@165415.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@165415.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@165429.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@165429.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@165429.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@165429.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@165429.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@165429.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@165443.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@165443.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@165443.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@165443.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@165443.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@165443.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@165457.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@165457.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@165457.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@165457.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@165457.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@165457.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@165471.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@165471.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@165471.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@165471.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@165471.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@165471.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@165485.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@165485.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@165485.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@165485.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@165485.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@165485.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@165499.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@165499.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@165499.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@165499.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@165499.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@165499.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@165513.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@165513.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@165513.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@165513.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@165513.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@165513.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@165527.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@165527.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@165527.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@165527.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@165527.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@165527.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@165541.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@165541.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@165541.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@165541.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@165541.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@165541.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@165555.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@165555.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@165555.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@165555.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@165555.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@165555.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@165569.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@165569.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@165569.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@165569.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@165569.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@165569.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@165583.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@165583.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@165583.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@165583.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@165583.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@165583.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@165597.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@165597.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@165597.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@165597.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@165597.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@165597.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@165611.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@165611.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@165611.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@165611.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@165611.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@165611.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@165625.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@165625.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@165625.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@165625.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@165625.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@165625.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@165639.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@165639.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@165639.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@165639.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@165639.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@165639.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@165653.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@165653.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@165653.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@165653.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@165653.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@165653.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@165667.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@165667.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@165667.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@165667.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@165667.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@165667.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@165681.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@165681.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@165681.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@165681.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@165681.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@165681.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@165695.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@165695.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@165695.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@165695.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@165695.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@165695.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@165709.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@165709.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@165709.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@165709.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@165709.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@165709.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@165723.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@165723.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@165723.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@165723.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@165723.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@165723.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@165737.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@165737.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@165737.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@165737.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@165737.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@165737.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@165751.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@165751.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@165751.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@165751.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@165751.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@165751.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@165765.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@165765.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@165765.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@165765.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@165765.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@165765.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@165779.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@165779.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@165779.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@165779.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@165779.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@165779.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@165793.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@165793.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@165793.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@165793.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@165793.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@165793.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@165807.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@165807.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@165807.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@165807.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@165807.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@165807.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@165821.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@165821.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@165821.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@165821.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@165821.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@165821.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@165835.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@165835.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@165835.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@165835.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@165835.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@165835.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@165849.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@165849.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@165849.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@165849.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@165849.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@165849.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@165863.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@165863.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@165863.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@165863.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@165863.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@165863.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@165877.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@165877.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@165877.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@165877.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@165877.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@165877.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@165891.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@165891.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@165891.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@165891.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@165891.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@165891.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@165905.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@165905.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@165905.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@165905.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@165905.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@165905.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@165919.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@165919.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@165919.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@165919.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@165919.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@165919.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@165933.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@165933.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@165933.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@165933.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@165933.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@165933.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@165947.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@165947.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@165947.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@165947.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@165947.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@165947.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@165961.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@165961.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@165961.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@165961.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@165961.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@165961.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@165975.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@165975.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@165975.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@165975.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@165975.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@165975.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@165989.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@165989.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@165989.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@165989.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@165989.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@165989.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@166003.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@166003.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@166003.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@166003.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@166003.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@166003.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@166017.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@166017.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@166017.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@166017.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@166017.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@166017.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@166031.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@166031.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@166031.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@166031.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@166031.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@166031.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@166045.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@166045.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@166045.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@166045.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@166045.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@166045.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@166059.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@166059.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@166059.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@166059.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@166059.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@166059.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@166073.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@166073.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@166073.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@166073.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@166073.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@166073.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@166087.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@166087.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@166087.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@166087.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@166087.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@166087.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@166101.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@166101.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@166101.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@166101.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@166101.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@166101.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@166115.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@166115.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@166115.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@166115.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@166115.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@166115.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@166129.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@166129.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@166129.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@166129.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@166129.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@166129.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@166143.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@166143.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@166143.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@166143.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@166143.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@166143.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@166157.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@166157.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@166157.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@166157.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@166157.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@166157.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@166171.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@166171.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@166171.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@166171.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@166171.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@166171.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@166185.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@166185.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@166185.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@166185.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@166185.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@166185.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@166199.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@166199.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@166199.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@166199.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@166199.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@166199.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@166213.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@166213.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@166213.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@166213.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@166213.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@166213.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@166227.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@166227.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@166227.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@166227.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@166227.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@166227.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@166241.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@166241.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@166241.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@166241.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@166241.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@166241.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@166255.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@166255.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@166255.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@166255.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@166255.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@166255.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@166269.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@166269.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@166269.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@166269.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@166269.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@166269.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@166283.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@166283.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@166283.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@166283.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@166283.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@166283.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@166297.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@166297.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@166297.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@166297.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@166297.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@166297.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@166311.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@166311.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@166311.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@166311.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@166311.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@166311.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@166325.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@166325.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@166325.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@166325.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@166325.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@166325.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@166339.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@166339.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@166339.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@166339.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@166339.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@166339.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@166353.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@166353.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@166353.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@166353.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@166353.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@166353.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@166367.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@166367.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@166367.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@166367.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@166367.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@166367.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@166381.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@166381.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@166381.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@166381.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@166381.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@166381.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@166395.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@166395.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@166395.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@166395.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@166395.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@166395.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@166409.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@166409.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@166409.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@166409.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@166409.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@166409.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@166423.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@166423.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@166423.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@166423.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@166423.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@166423.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@166437.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@166437.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@166437.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@166437.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@166437.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@166437.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@166451.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@166451.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@166451.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@166451.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@166451.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@166451.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@166465.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@166465.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@166465.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@166465.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@166465.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@166465.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@166479.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@166479.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@166479.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@166479.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@166479.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@166479.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@166493.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@166493.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@166493.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@166493.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@166493.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@166493.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@166507.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@166507.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@166507.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@166507.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@166507.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@166507.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@166521.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@166521.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@166521.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@166521.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@166521.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@166521.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@166535.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@166535.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@166535.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@166535.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@166535.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@166535.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@166549.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@166549.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@166549.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@166549.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@166549.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@166549.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@166563.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@166563.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@166563.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@166563.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@166563.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@166563.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@166577.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@166577.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@166577.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@166577.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@166577.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@166577.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@166591.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@166591.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@166591.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@166591.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@166591.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@166591.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@166605.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@166605.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@166605.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@166605.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@166605.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@166605.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@166619.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@166619.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@166619.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@166619.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@166619.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@166619.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@166633.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@166633.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@166633.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@166633.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@166633.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@166633.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@166647.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@166647.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@166647.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@166647.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@166647.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@166647.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@166661.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@166661.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@166661.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@166661.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@166661.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@166661.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@166675.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@166675.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@166675.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@166675.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@166675.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@166675.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@166689.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@166689.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@166689.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@166689.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@166689.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@166689.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@166703.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@166703.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@166703.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@166703.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@166703.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@166703.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@166717.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@166717.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@166717.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@166717.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@166717.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@166717.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@166731.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@166731.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@166731.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@166731.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@166731.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@166731.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@166745.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@166745.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@166745.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@166745.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@166745.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@166745.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@166759.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@166759.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@166759.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@166759.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@166759.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@166759.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@166773.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@166773.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@166773.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@166773.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@166773.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@166773.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@166787.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@166787.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@166787.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@166787.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@166787.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@166787.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@166801.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@166801.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@166801.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@166801.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@166801.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@166801.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@166815.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@166815.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@166815.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@166815.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@166815.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@166815.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@166829.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@166829.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@166829.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@166829.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@166829.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@166829.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@166843.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@166843.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@166843.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@166843.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@166843.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@166843.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@166857.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@166857.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@166857.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@166857.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@166857.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@166857.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@166871.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@166871.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@166871.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@166871.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@166871.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@166871.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@166885.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@166885.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@166885.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@166885.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@166885.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@166885.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@166899.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@166899.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@166899.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@166899.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@166899.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@166899.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@166913.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@166913.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@166913.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@166913.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@166913.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@166913.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@166927.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@166927.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@166927.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@166927.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@166927.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@166927.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@166941.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@166941.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@166941.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@166941.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@166941.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@166941.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@166955.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@166955.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@166955.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@166955.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@166955.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@166955.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@166969.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@166969.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@166969.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@166969.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@166969.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@166969.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@166983.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@166983.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@166983.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@166983.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@166983.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@166983.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@166997.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@166997.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@166997.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@166997.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@166997.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@166997.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@167011.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@167011.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@167011.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@167011.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@167011.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@167011.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@167025.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@167025.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@167025.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@167025.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@167025.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@167025.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@167039.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@167039.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@167039.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@167039.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@167039.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@167039.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@167053.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@167053.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@167053.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@167053.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@167053.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@167053.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@167067.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@167067.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@167067.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@167067.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@167067.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@167067.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@167081.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@167081.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@167081.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@167081.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@167081.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@167081.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@167095.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@167095.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@167095.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@167095.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@167095.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@167095.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@167109.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@167109.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@167109.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@167109.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@167109.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@167109.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@167123.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@167123.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@167123.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@167123.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@167123.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@167123.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@167137.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@167137.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@167137.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@167137.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@167137.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@167137.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@167151.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@167151.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@167151.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@167151.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@167151.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@167151.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@167165.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@167165.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@167165.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@167165.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@167165.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@167165.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@167179.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@167179.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@167179.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@167179.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@167179.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@167179.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@167193.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@167193.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@167193.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@167193.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@167193.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@167193.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@167207.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@167207.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@167207.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@167207.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@167207.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@167207.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@167221.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@167221.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@167221.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@167221.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@167221.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@167221.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@167235.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@167235.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@167235.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@167235.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@167235.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@167235.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@167249.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@167249.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@167249.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@167249.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@167249.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@167249.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@167263.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@167263.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@167263.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@167263.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@167263.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@167263.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@167277.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@167277.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@167277.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@167277.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@167277.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@167277.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@167291.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@167291.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@167291.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@167291.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@167291.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@167291.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@167305.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@167305.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@167305.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@167305.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@167305.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@167305.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@167319.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@167319.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@167319.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@167319.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@167319.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@167319.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@167333.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@167333.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@167333.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@167333.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@167333.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@167333.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@167347.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@167347.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@167347.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@167347.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@167347.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@167347.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@167361.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@167361.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@167361.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@167361.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@167361.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@167361.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@167375.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@167375.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@167375.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@167375.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@167375.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@167375.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@167389.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@167389.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@167389.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@167389.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@167389.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@167389.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@167403.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@167403.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@167403.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@167403.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@167403.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@167403.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@167417.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@167417.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@167417.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@167417.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@167417.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@167417.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@167431.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@167431.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@167431.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@167431.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@167431.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@167431.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@167445.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@167445.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@167445.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@167445.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@167445.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@167445.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@167459.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@167459.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@167459.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@167459.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@167459.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@167459.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@167473.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@167473.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@167473.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@167473.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@167473.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@167473.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@167487.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@167487.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@167487.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@167487.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@167487.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@167487.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@167501.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@167501.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@167501.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@167501.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@167501.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@167501.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@167515.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@167515.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@167515.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@167515.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@167515.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@167515.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@167529.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@167529.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@167529.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@167529.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@167529.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@167529.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@167543.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@167543.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@167543.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@167543.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@167543.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@167543.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@167557.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@167557.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@167557.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@167557.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@167557.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@167557.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@167571.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@167571.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@167571.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@167571.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@167571.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@167571.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@167585.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@167585.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@167585.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@167585.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@167585.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@167585.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@167599.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@167599.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@167599.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@167599.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@167599.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@167599.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@167613.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@167613.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@167613.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@167613.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@167613.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@167613.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@167627.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@167627.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@167627.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@167627.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@167627.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@167627.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@167641.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@167641.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@167641.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@167641.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@167641.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@167641.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@167655.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@167655.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@167655.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@167655.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@167655.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@167655.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@167669.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@167669.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@167669.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@167669.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@167669.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@167669.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@167683.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@167683.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@167683.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@167683.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@167683.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@167683.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@167697.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@167697.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@167697.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@167697.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@167697.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@167697.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@167711.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@167711.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@167711.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@167711.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@167711.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@167711.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@167725.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@167725.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@167725.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@167725.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@167725.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@167725.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@167739.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@167739.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@167739.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@167739.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@167739.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@167739.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@167753.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@167753.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@167753.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@167753.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@167753.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@167753.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@167767.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@167767.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@167767.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@167767.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@167767.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@167767.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@167781.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@167781.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@167781.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@167781.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@167781.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@167781.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@167795.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@167795.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@167795.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@167795.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@167795.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@167795.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@167809.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@167809.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@167809.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@167809.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@167809.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@167809.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@167823.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@167823.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@167823.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@167823.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@167823.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@167823.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@167837.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@167837.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@167837.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@167837.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@167837.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@167837.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@167851.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@167851.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@167851.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@167851.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@167851.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@167851.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@167865.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@167865.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@167865.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@167865.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@167865.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@167865.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@167879.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@167879.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@167879.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@167879.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@167879.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@167879.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@167893.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@167893.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@167893.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@167893.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@167893.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@167893.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@167907.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@167907.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@167907.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@167907.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@167907.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@167907.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@167921.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@167921.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@167921.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@167921.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@167921.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@167921.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@167935.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@167935.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@167935.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@167935.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@167935.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@167935.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@167949.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@167949.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@167949.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@167949.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@167949.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@167949.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@167963.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@167963.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@167963.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@167963.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@167963.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@167963.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@167977.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@167977.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@167977.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@167977.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@167977.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@167977.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@167991.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@167991.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@167991.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@167991.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@167991.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@167991.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@168005.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@168005.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@168005.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@168005.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@168005.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@168005.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@168019.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@168019.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@168019.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@168019.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@168019.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@168019.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@168033.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@168033.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@168033.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@168033.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@168033.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@168033.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@168047.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@168047.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@168047.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@168047.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@168047.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@168047.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@168061.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@168061.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@168061.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@168061.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@168061.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@168061.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@168075.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@168075.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@168075.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@168075.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@168075.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@168075.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@168089.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@168089.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@168089.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@168089.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@168089.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@168089.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@168103.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@168103.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@168103.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@168103.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@168103.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@168103.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@168117.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@168117.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@168117.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@168117.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@168117.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@168117.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@168131.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@168131.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@168131.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@168131.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@168131.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@168131.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@168145.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@168145.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@168145.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@168145.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@168145.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@168145.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@168159.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@168159.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@168159.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@168159.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@168159.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@168159.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@168173.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@168173.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@168173.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@168173.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@168173.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@168173.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@168187.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@168187.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@168187.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@168187.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@168187.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@168187.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@168201.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@168201.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@168201.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@168201.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@168201.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@168201.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@168215.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@168215.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@168215.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@168215.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@168215.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@168215.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@168229.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@168229.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@168229.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@168229.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@168229.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@168229.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@168243.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@168243.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@168243.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@168243.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@168243.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@168243.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@168257.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@168257.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@168257.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@168257.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@168257.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@168257.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@168271.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@168271.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@168271.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@168271.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@168271.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@168271.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@168285.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@168285.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@168285.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@168285.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@168285.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@168285.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@168299.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@168299.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@168299.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@168299.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@168299.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@168299.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@168313.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@168313.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@168313.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@168313.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@168313.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@168313.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@168327.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@168327.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@168327.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@168327.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@168327.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@168327.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@168341.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@168341.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@168341.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@168341.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@168341.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@168341.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@168355.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@168355.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@168355.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@168355.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@168355.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@168355.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@168369.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@168369.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@168369.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@168369.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@168369.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@168369.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@168383.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@168383.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@168383.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@168383.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@168383.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@168383.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@168397.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@168397.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@168397.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@168397.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@168397.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@168397.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@168411.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@168411.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@168411.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@168411.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@168411.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@168411.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@168425.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@168425.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@168425.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@168425.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@168425.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@168425.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@168439.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@168439.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@168439.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@168439.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@168439.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@168439.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@168453.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@168453.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@168453.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@168453.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@168453.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@168453.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@168467.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@168467.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@168467.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@168467.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@168467.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@168467.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@168481.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@168481.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@168481.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@168481.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@168481.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@168481.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@168495.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@168495.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@168495.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@168495.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@168495.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@168495.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@168509.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@168509.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@168509.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@168509.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@168509.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@168509.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@168523.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@168523.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@168523.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@168523.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@168523.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@168523.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@168537.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@168537.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@168537.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@168537.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@168537.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@168537.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@168551.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@168551.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@168551.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@168551.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@168551.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@168551.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@168565.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@168565.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@168565.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@168565.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@168565.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@168565.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@168579.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@168579.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@168579.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@168579.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@168579.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@168579.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@168593.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@168593.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@168593.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@168593.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@168593.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@168593.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@168607.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@168607.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@168607.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@168607.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@168607.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@168607.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@168621.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@168621.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@168621.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@168621.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@168621.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@168621.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@168635.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@168635.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@168635.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@168635.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@168635.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@168635.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@168649.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@168649.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@168649.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@168649.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@168649.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@168649.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@168663.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@168663.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@168663.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@168663.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@168663.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@168663.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@168677.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@168677.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@168677.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@168677.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@168677.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@168677.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@168691.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@168691.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@168691.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@168691.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@168691.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@168691.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@168705.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@168705.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@168705.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@168705.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@168705.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@168705.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@168719.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@168719.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@168719.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@168719.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@168719.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@168719.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@168733.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@168733.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@168733.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@168733.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@168733.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@168733.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@168747.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@168747.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@168747.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@168747.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@168747.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@168747.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@168761.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@168761.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@168761.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@168761.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@168761.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@168761.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@168775.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@168775.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@168775.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@168775.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@168775.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@168775.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@168789.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@168789.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@168789.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@168789.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@168789.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@168789.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@168803.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@168803.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@168803.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@168803.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@168803.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@168803.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@168817.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@168817.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@168817.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@168817.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@168817.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@168817.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@168831.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@168831.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@168831.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@161793.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@161805.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@161806.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@161824.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@161836.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@161848.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@161849.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@161790.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@161802.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@161821.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@161833.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@161845.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@161859.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@161873.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@161887.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@161901.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@161915.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@161929.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@161943.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@161957.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@161971.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@161985.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@161999.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@162013.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@162027.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@162041.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@162055.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@162069.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@162083.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@162097.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@162111.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@162125.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@162139.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@162153.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@162167.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@162181.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@162195.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@162209.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@162223.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@162237.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@162251.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@162265.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@162279.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@162293.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@162307.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@162321.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@162335.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@162349.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@162363.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@162377.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@162391.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@162405.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@162419.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@162433.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@162447.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@162461.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@162475.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@162489.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@162503.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@162517.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@162531.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@162545.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@162559.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@162573.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@162587.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@162601.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@162615.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@162629.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@162643.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@162657.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@162671.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@162685.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@162699.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@162713.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@162727.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@162741.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@162755.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@162769.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@162783.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@162797.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@162811.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@162825.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@162839.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@162853.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@162867.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@162881.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@162895.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@162909.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@162923.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@162937.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@162951.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@162965.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@162979.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@162993.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@163007.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@163021.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@163035.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@163049.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@163063.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@163077.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@163091.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@163105.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@163119.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@163133.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@163147.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@163161.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@163175.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@163189.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@163203.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@163217.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@163231.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@163245.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@163259.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@163273.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@163287.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@163301.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@163315.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@163329.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@163343.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@163357.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@163371.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@163385.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@163399.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@163413.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@163427.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@163441.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@163455.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@163469.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@163483.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@163497.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@163511.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@163525.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@163539.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@163553.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@163567.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@163581.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@163595.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@163609.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@163623.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@163637.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@163651.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@163665.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@163679.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@163693.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@163707.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@163721.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@163735.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@163749.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@163763.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@163777.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@163791.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@163805.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@163819.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@163833.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@163847.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@163861.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@163875.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@163889.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@163903.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@163917.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@163931.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@163945.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@163959.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@163973.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@163987.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@164001.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@164015.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@164029.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@164043.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@164057.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@164071.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@164085.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@164099.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@164113.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@164127.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@164141.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@164155.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@164169.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@164183.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@164197.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@164211.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@164225.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@164239.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@164253.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@164267.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@164281.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@164295.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@164309.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@164323.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@164337.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@164351.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@164365.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@164379.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@164393.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@164407.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@164421.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@164435.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@164449.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@164463.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@164477.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@164491.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@164505.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@164519.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@164533.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@164547.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@164561.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@164575.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@164589.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@164603.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@164617.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@164631.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@164645.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@164659.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@164673.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@164687.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@164701.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@164715.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@164729.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@164743.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@164757.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@164771.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@164785.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@164799.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@164813.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@164827.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@164841.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@164855.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@164869.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@164883.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@164897.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@164911.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@164925.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@164939.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@164953.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@164967.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@164981.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@164995.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@165009.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@165023.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@165037.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@165051.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@165065.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@165079.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@165093.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@165107.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@165121.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@165135.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@165149.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@165163.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@165177.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@165191.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@165205.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@165219.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@165233.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@165247.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@165261.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@165275.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@165289.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@165303.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@165317.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@165331.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@165345.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@165359.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@165373.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@165387.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@165401.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@165415.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@165429.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@165443.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@165457.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@165471.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@165485.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@165499.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@165513.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@165527.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@165541.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@165555.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@165569.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@165583.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@165597.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@165611.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@165625.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@165639.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@165653.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@165667.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@165681.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@165695.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@165709.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@165723.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@165737.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@165751.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@165765.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@165779.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@165793.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@165807.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@165821.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@165835.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@165849.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@165863.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@165877.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@165891.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@165905.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@165919.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@165933.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@165947.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@165961.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@165975.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@165989.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@166003.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@166017.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@166031.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@166045.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@166059.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@166073.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@166087.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@166101.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@166115.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@166129.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@166143.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@166157.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@166171.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@166185.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@166199.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@166213.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@166227.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@166241.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@166255.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@166269.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@166283.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@166297.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@166311.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@166325.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@166339.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@166353.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@166367.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@166381.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@166395.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@166409.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@166423.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@166437.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@166451.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@166465.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@166479.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@166493.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@166507.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@166521.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@166535.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@166549.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@166563.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@166577.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@166591.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@166605.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@166619.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@166633.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@166647.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@166661.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@166675.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@166689.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@166703.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@166717.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@166731.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@166745.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@166759.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@166773.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@166787.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@166801.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@166815.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@166829.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@166843.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@166857.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@166871.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@166885.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@166899.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@166913.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@166927.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@166941.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@166955.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@166969.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@166983.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@166997.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@167011.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@167025.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@167039.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@167053.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@167067.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@167081.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@167095.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@167109.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@167123.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@167137.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@167151.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@167165.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@167179.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@167193.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@167207.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@167221.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@167235.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@167249.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@167263.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@167277.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@167291.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@167305.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@167319.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@167333.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@167347.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@167361.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@167375.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@167389.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@167403.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@167417.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@167431.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@167445.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@167459.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@167473.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@167487.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@167501.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@167515.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@167529.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@167543.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@167557.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@167571.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@167585.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@167599.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@167613.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@167627.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@167641.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@167655.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@167669.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@167683.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@167697.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@167711.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@167725.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@167739.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@167753.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@167767.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@167781.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@167795.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@167809.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@167823.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@167837.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@167851.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@167865.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@167879.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@167893.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@167907.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@167921.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@167935.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@167949.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@167963.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@167977.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@167991.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@168005.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@168019.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@168033.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@168047.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@168061.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@168075.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@168089.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@168103.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@168117.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@168131.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@168145.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@168159.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@168173.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@168187.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@168201.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@168215.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@168229.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@168243.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@168257.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@168271.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@168285.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@168299.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@168313.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@168327.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@168341.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@168355.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@168369.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@168383.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@168397.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@168411.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@168425.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@168439.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@168453.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@168467.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@168481.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@168495.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@168509.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@168523.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@168537.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@168551.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@168565.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@168579.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@168593.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@168607.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@168621.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@168635.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@168649.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@168663.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@168677.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@168691.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@168705.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@168719.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@168733.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@168747.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@168761.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@168775.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@168789.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@168803.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@168817.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@168831.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@161793.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@161805.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@161806.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@161824.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@161836.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@161848.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@161849.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@169842.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@169848.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@169849.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@169850.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@169851.4]
  assign regs_0_clock = clock; // @[:@161791.4]
  assign regs_0_reset = reset; // @[:@161792.4 RegFile.scala 82:16:@161798.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@161796.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@161800.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@161795.4]
  assign regs_1_clock = clock; // @[:@161803.4]
  assign regs_1_reset = reset; // @[:@161804.4 RegFile.scala 70:16:@161816.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@161814.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@161819.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@161810.4]
  assign regs_2_clock = clock; // @[:@161822.4]
  assign regs_2_reset = reset; // @[:@161823.4 RegFile.scala 82:16:@161829.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@161827.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@161831.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@161826.4]
  assign regs_3_clock = clock; // @[:@161834.4]
  assign regs_3_reset = reset; // @[:@161835.4 RegFile.scala 82:16:@161841.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@161839.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@161843.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@161838.4]
  assign regs_4_clock = clock; // @[:@161846.4]
  assign regs_4_reset = io_reset; // @[:@161847.4 RegFile.scala 76:16:@161854.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@161853.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@161857.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@161851.4]
  assign regs_5_clock = clock; // @[:@161860.4]
  assign regs_5_reset = io_reset; // @[:@161861.4 RegFile.scala 76:16:@161868.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@161867.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@161871.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@161865.4]
  assign regs_6_clock = clock; // @[:@161874.4]
  assign regs_6_reset = io_reset; // @[:@161875.4 RegFile.scala 76:16:@161882.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@161881.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@161885.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@161879.4]
  assign regs_7_clock = clock; // @[:@161888.4]
  assign regs_7_reset = io_reset; // @[:@161889.4 RegFile.scala 76:16:@161896.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@161895.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@161899.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@161893.4]
  assign regs_8_clock = clock; // @[:@161902.4]
  assign regs_8_reset = io_reset; // @[:@161903.4 RegFile.scala 76:16:@161910.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@161909.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@161913.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@161907.4]
  assign regs_9_clock = clock; // @[:@161916.4]
  assign regs_9_reset = io_reset; // @[:@161917.4 RegFile.scala 76:16:@161924.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@161923.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@161927.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@161921.4]
  assign regs_10_clock = clock; // @[:@161930.4]
  assign regs_10_reset = io_reset; // @[:@161931.4 RegFile.scala 76:16:@161938.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@161937.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@161941.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@161935.4]
  assign regs_11_clock = clock; // @[:@161944.4]
  assign regs_11_reset = io_reset; // @[:@161945.4 RegFile.scala 76:16:@161952.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@161951.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@161955.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@161949.4]
  assign regs_12_clock = clock; // @[:@161958.4]
  assign regs_12_reset = io_reset; // @[:@161959.4 RegFile.scala 76:16:@161966.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@161965.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@161969.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@161963.4]
  assign regs_13_clock = clock; // @[:@161972.4]
  assign regs_13_reset = io_reset; // @[:@161973.4 RegFile.scala 76:16:@161980.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@161979.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@161983.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@161977.4]
  assign regs_14_clock = clock; // @[:@161986.4]
  assign regs_14_reset = io_reset; // @[:@161987.4 RegFile.scala 76:16:@161994.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@161993.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@161997.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@161991.4]
  assign regs_15_clock = clock; // @[:@162000.4]
  assign regs_15_reset = io_reset; // @[:@162001.4 RegFile.scala 76:16:@162008.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@162007.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@162011.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@162005.4]
  assign regs_16_clock = clock; // @[:@162014.4]
  assign regs_16_reset = io_reset; // @[:@162015.4 RegFile.scala 76:16:@162022.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@162021.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@162025.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@162019.4]
  assign regs_17_clock = clock; // @[:@162028.4]
  assign regs_17_reset = io_reset; // @[:@162029.4 RegFile.scala 76:16:@162036.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@162035.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@162039.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@162033.4]
  assign regs_18_clock = clock; // @[:@162042.4]
  assign regs_18_reset = io_reset; // @[:@162043.4 RegFile.scala 76:16:@162050.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@162049.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@162053.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@162047.4]
  assign regs_19_clock = clock; // @[:@162056.4]
  assign regs_19_reset = io_reset; // @[:@162057.4 RegFile.scala 76:16:@162064.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@162063.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@162067.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@162061.4]
  assign regs_20_clock = clock; // @[:@162070.4]
  assign regs_20_reset = io_reset; // @[:@162071.4 RegFile.scala 76:16:@162078.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@162077.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@162081.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@162075.4]
  assign regs_21_clock = clock; // @[:@162084.4]
  assign regs_21_reset = io_reset; // @[:@162085.4 RegFile.scala 76:16:@162092.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@162091.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@162095.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@162089.4]
  assign regs_22_clock = clock; // @[:@162098.4]
  assign regs_22_reset = io_reset; // @[:@162099.4 RegFile.scala 76:16:@162106.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@162105.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@162109.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@162103.4]
  assign regs_23_clock = clock; // @[:@162112.4]
  assign regs_23_reset = io_reset; // @[:@162113.4 RegFile.scala 76:16:@162120.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@162119.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@162123.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@162117.4]
  assign regs_24_clock = clock; // @[:@162126.4]
  assign regs_24_reset = io_reset; // @[:@162127.4 RegFile.scala 76:16:@162134.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@162133.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@162137.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@162131.4]
  assign regs_25_clock = clock; // @[:@162140.4]
  assign regs_25_reset = io_reset; // @[:@162141.4 RegFile.scala 76:16:@162148.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@162147.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@162151.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@162145.4]
  assign regs_26_clock = clock; // @[:@162154.4]
  assign regs_26_reset = io_reset; // @[:@162155.4 RegFile.scala 76:16:@162162.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@162161.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@162165.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@162159.4]
  assign regs_27_clock = clock; // @[:@162168.4]
  assign regs_27_reset = io_reset; // @[:@162169.4 RegFile.scala 76:16:@162176.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@162175.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@162179.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@162173.4]
  assign regs_28_clock = clock; // @[:@162182.4]
  assign regs_28_reset = io_reset; // @[:@162183.4 RegFile.scala 76:16:@162190.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@162189.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@162193.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@162187.4]
  assign regs_29_clock = clock; // @[:@162196.4]
  assign regs_29_reset = io_reset; // @[:@162197.4 RegFile.scala 76:16:@162204.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@162203.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@162207.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@162201.4]
  assign regs_30_clock = clock; // @[:@162210.4]
  assign regs_30_reset = io_reset; // @[:@162211.4 RegFile.scala 76:16:@162218.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@162217.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@162221.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@162215.4]
  assign regs_31_clock = clock; // @[:@162224.4]
  assign regs_31_reset = io_reset; // @[:@162225.4 RegFile.scala 76:16:@162232.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@162231.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@162235.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@162229.4]
  assign regs_32_clock = clock; // @[:@162238.4]
  assign regs_32_reset = io_reset; // @[:@162239.4 RegFile.scala 76:16:@162246.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@162245.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@162249.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@162243.4]
  assign regs_33_clock = clock; // @[:@162252.4]
  assign regs_33_reset = io_reset; // @[:@162253.4 RegFile.scala 76:16:@162260.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@162259.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@162263.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@162257.4]
  assign regs_34_clock = clock; // @[:@162266.4]
  assign regs_34_reset = io_reset; // @[:@162267.4 RegFile.scala 76:16:@162274.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@162273.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@162277.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@162271.4]
  assign regs_35_clock = clock; // @[:@162280.4]
  assign regs_35_reset = io_reset; // @[:@162281.4 RegFile.scala 76:16:@162288.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@162287.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@162291.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@162285.4]
  assign regs_36_clock = clock; // @[:@162294.4]
  assign regs_36_reset = io_reset; // @[:@162295.4 RegFile.scala 76:16:@162302.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@162301.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@162305.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@162299.4]
  assign regs_37_clock = clock; // @[:@162308.4]
  assign regs_37_reset = io_reset; // @[:@162309.4 RegFile.scala 76:16:@162316.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@162315.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@162319.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@162313.4]
  assign regs_38_clock = clock; // @[:@162322.4]
  assign regs_38_reset = io_reset; // @[:@162323.4 RegFile.scala 76:16:@162330.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@162329.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@162333.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@162327.4]
  assign regs_39_clock = clock; // @[:@162336.4]
  assign regs_39_reset = io_reset; // @[:@162337.4 RegFile.scala 76:16:@162344.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@162343.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@162347.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@162341.4]
  assign regs_40_clock = clock; // @[:@162350.4]
  assign regs_40_reset = io_reset; // @[:@162351.4 RegFile.scala 76:16:@162358.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@162357.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@162361.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@162355.4]
  assign regs_41_clock = clock; // @[:@162364.4]
  assign regs_41_reset = io_reset; // @[:@162365.4 RegFile.scala 76:16:@162372.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@162371.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@162375.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@162369.4]
  assign regs_42_clock = clock; // @[:@162378.4]
  assign regs_42_reset = io_reset; // @[:@162379.4 RegFile.scala 76:16:@162386.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@162385.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@162389.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@162383.4]
  assign regs_43_clock = clock; // @[:@162392.4]
  assign regs_43_reset = io_reset; // @[:@162393.4 RegFile.scala 76:16:@162400.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@162399.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@162403.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@162397.4]
  assign regs_44_clock = clock; // @[:@162406.4]
  assign regs_44_reset = io_reset; // @[:@162407.4 RegFile.scala 76:16:@162414.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@162413.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@162417.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@162411.4]
  assign regs_45_clock = clock; // @[:@162420.4]
  assign regs_45_reset = io_reset; // @[:@162421.4 RegFile.scala 76:16:@162428.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@162427.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@162431.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@162425.4]
  assign regs_46_clock = clock; // @[:@162434.4]
  assign regs_46_reset = io_reset; // @[:@162435.4 RegFile.scala 76:16:@162442.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@162441.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@162445.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@162439.4]
  assign regs_47_clock = clock; // @[:@162448.4]
  assign regs_47_reset = io_reset; // @[:@162449.4 RegFile.scala 76:16:@162456.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@162455.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@162459.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@162453.4]
  assign regs_48_clock = clock; // @[:@162462.4]
  assign regs_48_reset = io_reset; // @[:@162463.4 RegFile.scala 76:16:@162470.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@162469.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@162473.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@162467.4]
  assign regs_49_clock = clock; // @[:@162476.4]
  assign regs_49_reset = io_reset; // @[:@162477.4 RegFile.scala 76:16:@162484.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@162483.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@162487.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@162481.4]
  assign regs_50_clock = clock; // @[:@162490.4]
  assign regs_50_reset = io_reset; // @[:@162491.4 RegFile.scala 76:16:@162498.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@162497.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@162501.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@162495.4]
  assign regs_51_clock = clock; // @[:@162504.4]
  assign regs_51_reset = io_reset; // @[:@162505.4 RegFile.scala 76:16:@162512.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@162511.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@162515.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@162509.4]
  assign regs_52_clock = clock; // @[:@162518.4]
  assign regs_52_reset = io_reset; // @[:@162519.4 RegFile.scala 76:16:@162526.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@162525.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@162529.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@162523.4]
  assign regs_53_clock = clock; // @[:@162532.4]
  assign regs_53_reset = io_reset; // @[:@162533.4 RegFile.scala 76:16:@162540.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@162539.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@162543.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@162537.4]
  assign regs_54_clock = clock; // @[:@162546.4]
  assign regs_54_reset = io_reset; // @[:@162547.4 RegFile.scala 76:16:@162554.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@162553.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@162557.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@162551.4]
  assign regs_55_clock = clock; // @[:@162560.4]
  assign regs_55_reset = io_reset; // @[:@162561.4 RegFile.scala 76:16:@162568.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@162567.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@162571.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@162565.4]
  assign regs_56_clock = clock; // @[:@162574.4]
  assign regs_56_reset = io_reset; // @[:@162575.4 RegFile.scala 76:16:@162582.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@162581.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@162585.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@162579.4]
  assign regs_57_clock = clock; // @[:@162588.4]
  assign regs_57_reset = io_reset; // @[:@162589.4 RegFile.scala 76:16:@162596.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@162595.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@162599.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@162593.4]
  assign regs_58_clock = clock; // @[:@162602.4]
  assign regs_58_reset = io_reset; // @[:@162603.4 RegFile.scala 76:16:@162610.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@162609.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@162613.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@162607.4]
  assign regs_59_clock = clock; // @[:@162616.4]
  assign regs_59_reset = io_reset; // @[:@162617.4 RegFile.scala 76:16:@162624.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@162623.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@162627.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@162621.4]
  assign regs_60_clock = clock; // @[:@162630.4]
  assign regs_60_reset = io_reset; // @[:@162631.4 RegFile.scala 76:16:@162638.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@162637.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@162641.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@162635.4]
  assign regs_61_clock = clock; // @[:@162644.4]
  assign regs_61_reset = io_reset; // @[:@162645.4 RegFile.scala 76:16:@162652.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@162651.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@162655.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@162649.4]
  assign regs_62_clock = clock; // @[:@162658.4]
  assign regs_62_reset = io_reset; // @[:@162659.4 RegFile.scala 76:16:@162666.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@162665.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@162669.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@162663.4]
  assign regs_63_clock = clock; // @[:@162672.4]
  assign regs_63_reset = io_reset; // @[:@162673.4 RegFile.scala 76:16:@162680.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@162679.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@162683.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@162677.4]
  assign regs_64_clock = clock; // @[:@162686.4]
  assign regs_64_reset = io_reset; // @[:@162687.4 RegFile.scala 76:16:@162694.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@162693.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@162697.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@162691.4]
  assign regs_65_clock = clock; // @[:@162700.4]
  assign regs_65_reset = io_reset; // @[:@162701.4 RegFile.scala 76:16:@162708.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@162707.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@162711.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@162705.4]
  assign regs_66_clock = clock; // @[:@162714.4]
  assign regs_66_reset = io_reset; // @[:@162715.4 RegFile.scala 76:16:@162722.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@162721.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@162725.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@162719.4]
  assign regs_67_clock = clock; // @[:@162728.4]
  assign regs_67_reset = io_reset; // @[:@162729.4 RegFile.scala 76:16:@162736.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@162735.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@162739.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@162733.4]
  assign regs_68_clock = clock; // @[:@162742.4]
  assign regs_68_reset = io_reset; // @[:@162743.4 RegFile.scala 76:16:@162750.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@162749.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@162753.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@162747.4]
  assign regs_69_clock = clock; // @[:@162756.4]
  assign regs_69_reset = io_reset; // @[:@162757.4 RegFile.scala 76:16:@162764.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@162763.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@162767.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@162761.4]
  assign regs_70_clock = clock; // @[:@162770.4]
  assign regs_70_reset = io_reset; // @[:@162771.4 RegFile.scala 76:16:@162778.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@162777.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@162781.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@162775.4]
  assign regs_71_clock = clock; // @[:@162784.4]
  assign regs_71_reset = io_reset; // @[:@162785.4 RegFile.scala 76:16:@162792.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@162791.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@162795.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@162789.4]
  assign regs_72_clock = clock; // @[:@162798.4]
  assign regs_72_reset = io_reset; // @[:@162799.4 RegFile.scala 76:16:@162806.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@162805.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@162809.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@162803.4]
  assign regs_73_clock = clock; // @[:@162812.4]
  assign regs_73_reset = io_reset; // @[:@162813.4 RegFile.scala 76:16:@162820.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@162819.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@162823.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@162817.4]
  assign regs_74_clock = clock; // @[:@162826.4]
  assign regs_74_reset = io_reset; // @[:@162827.4 RegFile.scala 76:16:@162834.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@162833.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@162837.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@162831.4]
  assign regs_75_clock = clock; // @[:@162840.4]
  assign regs_75_reset = io_reset; // @[:@162841.4 RegFile.scala 76:16:@162848.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@162847.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@162851.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@162845.4]
  assign regs_76_clock = clock; // @[:@162854.4]
  assign regs_76_reset = io_reset; // @[:@162855.4 RegFile.scala 76:16:@162862.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@162861.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@162865.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@162859.4]
  assign regs_77_clock = clock; // @[:@162868.4]
  assign regs_77_reset = io_reset; // @[:@162869.4 RegFile.scala 76:16:@162876.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@162875.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@162879.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@162873.4]
  assign regs_78_clock = clock; // @[:@162882.4]
  assign regs_78_reset = io_reset; // @[:@162883.4 RegFile.scala 76:16:@162890.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@162889.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@162893.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@162887.4]
  assign regs_79_clock = clock; // @[:@162896.4]
  assign regs_79_reset = io_reset; // @[:@162897.4 RegFile.scala 76:16:@162904.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@162903.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@162907.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@162901.4]
  assign regs_80_clock = clock; // @[:@162910.4]
  assign regs_80_reset = io_reset; // @[:@162911.4 RegFile.scala 76:16:@162918.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@162917.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@162921.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@162915.4]
  assign regs_81_clock = clock; // @[:@162924.4]
  assign regs_81_reset = io_reset; // @[:@162925.4 RegFile.scala 76:16:@162932.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@162931.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@162935.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@162929.4]
  assign regs_82_clock = clock; // @[:@162938.4]
  assign regs_82_reset = io_reset; // @[:@162939.4 RegFile.scala 76:16:@162946.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@162945.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@162949.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@162943.4]
  assign regs_83_clock = clock; // @[:@162952.4]
  assign regs_83_reset = io_reset; // @[:@162953.4 RegFile.scala 76:16:@162960.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@162959.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@162963.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@162957.4]
  assign regs_84_clock = clock; // @[:@162966.4]
  assign regs_84_reset = io_reset; // @[:@162967.4 RegFile.scala 76:16:@162974.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@162973.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@162977.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@162971.4]
  assign regs_85_clock = clock; // @[:@162980.4]
  assign regs_85_reset = io_reset; // @[:@162981.4 RegFile.scala 76:16:@162988.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@162987.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@162991.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@162985.4]
  assign regs_86_clock = clock; // @[:@162994.4]
  assign regs_86_reset = io_reset; // @[:@162995.4 RegFile.scala 76:16:@163002.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@163001.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@163005.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@162999.4]
  assign regs_87_clock = clock; // @[:@163008.4]
  assign regs_87_reset = io_reset; // @[:@163009.4 RegFile.scala 76:16:@163016.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@163015.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@163019.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@163013.4]
  assign regs_88_clock = clock; // @[:@163022.4]
  assign regs_88_reset = io_reset; // @[:@163023.4 RegFile.scala 76:16:@163030.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@163029.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@163033.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@163027.4]
  assign regs_89_clock = clock; // @[:@163036.4]
  assign regs_89_reset = io_reset; // @[:@163037.4 RegFile.scala 76:16:@163044.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@163043.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@163047.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@163041.4]
  assign regs_90_clock = clock; // @[:@163050.4]
  assign regs_90_reset = io_reset; // @[:@163051.4 RegFile.scala 76:16:@163058.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@163057.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@163061.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@163055.4]
  assign regs_91_clock = clock; // @[:@163064.4]
  assign regs_91_reset = io_reset; // @[:@163065.4 RegFile.scala 76:16:@163072.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@163071.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@163075.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@163069.4]
  assign regs_92_clock = clock; // @[:@163078.4]
  assign regs_92_reset = io_reset; // @[:@163079.4 RegFile.scala 76:16:@163086.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@163085.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@163089.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@163083.4]
  assign regs_93_clock = clock; // @[:@163092.4]
  assign regs_93_reset = io_reset; // @[:@163093.4 RegFile.scala 76:16:@163100.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@163099.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@163103.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@163097.4]
  assign regs_94_clock = clock; // @[:@163106.4]
  assign regs_94_reset = io_reset; // @[:@163107.4 RegFile.scala 76:16:@163114.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@163113.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@163117.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@163111.4]
  assign regs_95_clock = clock; // @[:@163120.4]
  assign regs_95_reset = io_reset; // @[:@163121.4 RegFile.scala 76:16:@163128.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@163127.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@163131.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@163125.4]
  assign regs_96_clock = clock; // @[:@163134.4]
  assign regs_96_reset = io_reset; // @[:@163135.4 RegFile.scala 76:16:@163142.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@163141.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@163145.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@163139.4]
  assign regs_97_clock = clock; // @[:@163148.4]
  assign regs_97_reset = io_reset; // @[:@163149.4 RegFile.scala 76:16:@163156.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@163155.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@163159.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@163153.4]
  assign regs_98_clock = clock; // @[:@163162.4]
  assign regs_98_reset = io_reset; // @[:@163163.4 RegFile.scala 76:16:@163170.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@163169.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@163173.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@163167.4]
  assign regs_99_clock = clock; // @[:@163176.4]
  assign regs_99_reset = io_reset; // @[:@163177.4 RegFile.scala 76:16:@163184.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@163183.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@163187.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@163181.4]
  assign regs_100_clock = clock; // @[:@163190.4]
  assign regs_100_reset = io_reset; // @[:@163191.4 RegFile.scala 76:16:@163198.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@163197.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@163201.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@163195.4]
  assign regs_101_clock = clock; // @[:@163204.4]
  assign regs_101_reset = io_reset; // @[:@163205.4 RegFile.scala 76:16:@163212.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@163211.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@163215.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@163209.4]
  assign regs_102_clock = clock; // @[:@163218.4]
  assign regs_102_reset = io_reset; // @[:@163219.4 RegFile.scala 76:16:@163226.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@163225.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@163229.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@163223.4]
  assign regs_103_clock = clock; // @[:@163232.4]
  assign regs_103_reset = io_reset; // @[:@163233.4 RegFile.scala 76:16:@163240.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@163239.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@163243.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@163237.4]
  assign regs_104_clock = clock; // @[:@163246.4]
  assign regs_104_reset = io_reset; // @[:@163247.4 RegFile.scala 76:16:@163254.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@163253.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@163257.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@163251.4]
  assign regs_105_clock = clock; // @[:@163260.4]
  assign regs_105_reset = io_reset; // @[:@163261.4 RegFile.scala 76:16:@163268.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@163267.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@163271.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@163265.4]
  assign regs_106_clock = clock; // @[:@163274.4]
  assign regs_106_reset = io_reset; // @[:@163275.4 RegFile.scala 76:16:@163282.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@163281.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@163285.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@163279.4]
  assign regs_107_clock = clock; // @[:@163288.4]
  assign regs_107_reset = io_reset; // @[:@163289.4 RegFile.scala 76:16:@163296.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@163295.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@163299.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@163293.4]
  assign regs_108_clock = clock; // @[:@163302.4]
  assign regs_108_reset = io_reset; // @[:@163303.4 RegFile.scala 76:16:@163310.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@163309.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@163313.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@163307.4]
  assign regs_109_clock = clock; // @[:@163316.4]
  assign regs_109_reset = io_reset; // @[:@163317.4 RegFile.scala 76:16:@163324.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@163323.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@163327.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@163321.4]
  assign regs_110_clock = clock; // @[:@163330.4]
  assign regs_110_reset = io_reset; // @[:@163331.4 RegFile.scala 76:16:@163338.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@163337.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@163341.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@163335.4]
  assign regs_111_clock = clock; // @[:@163344.4]
  assign regs_111_reset = io_reset; // @[:@163345.4 RegFile.scala 76:16:@163352.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@163351.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@163355.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@163349.4]
  assign regs_112_clock = clock; // @[:@163358.4]
  assign regs_112_reset = io_reset; // @[:@163359.4 RegFile.scala 76:16:@163366.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@163365.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@163369.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@163363.4]
  assign regs_113_clock = clock; // @[:@163372.4]
  assign regs_113_reset = io_reset; // @[:@163373.4 RegFile.scala 76:16:@163380.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@163379.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@163383.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@163377.4]
  assign regs_114_clock = clock; // @[:@163386.4]
  assign regs_114_reset = io_reset; // @[:@163387.4 RegFile.scala 76:16:@163394.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@163393.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@163397.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@163391.4]
  assign regs_115_clock = clock; // @[:@163400.4]
  assign regs_115_reset = io_reset; // @[:@163401.4 RegFile.scala 76:16:@163408.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@163407.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@163411.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@163405.4]
  assign regs_116_clock = clock; // @[:@163414.4]
  assign regs_116_reset = io_reset; // @[:@163415.4 RegFile.scala 76:16:@163422.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@163421.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@163425.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@163419.4]
  assign regs_117_clock = clock; // @[:@163428.4]
  assign regs_117_reset = io_reset; // @[:@163429.4 RegFile.scala 76:16:@163436.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@163435.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@163439.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@163433.4]
  assign regs_118_clock = clock; // @[:@163442.4]
  assign regs_118_reset = io_reset; // @[:@163443.4 RegFile.scala 76:16:@163450.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@163449.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@163453.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@163447.4]
  assign regs_119_clock = clock; // @[:@163456.4]
  assign regs_119_reset = io_reset; // @[:@163457.4 RegFile.scala 76:16:@163464.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@163463.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@163467.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@163461.4]
  assign regs_120_clock = clock; // @[:@163470.4]
  assign regs_120_reset = io_reset; // @[:@163471.4 RegFile.scala 76:16:@163478.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@163477.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@163481.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@163475.4]
  assign regs_121_clock = clock; // @[:@163484.4]
  assign regs_121_reset = io_reset; // @[:@163485.4 RegFile.scala 76:16:@163492.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@163491.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@163495.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@163489.4]
  assign regs_122_clock = clock; // @[:@163498.4]
  assign regs_122_reset = io_reset; // @[:@163499.4 RegFile.scala 76:16:@163506.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@163505.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@163509.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@163503.4]
  assign regs_123_clock = clock; // @[:@163512.4]
  assign regs_123_reset = io_reset; // @[:@163513.4 RegFile.scala 76:16:@163520.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@163519.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@163523.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@163517.4]
  assign regs_124_clock = clock; // @[:@163526.4]
  assign regs_124_reset = io_reset; // @[:@163527.4 RegFile.scala 76:16:@163534.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@163533.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@163537.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@163531.4]
  assign regs_125_clock = clock; // @[:@163540.4]
  assign regs_125_reset = io_reset; // @[:@163541.4 RegFile.scala 76:16:@163548.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@163547.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@163551.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@163545.4]
  assign regs_126_clock = clock; // @[:@163554.4]
  assign regs_126_reset = io_reset; // @[:@163555.4 RegFile.scala 76:16:@163562.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@163561.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@163565.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@163559.4]
  assign regs_127_clock = clock; // @[:@163568.4]
  assign regs_127_reset = io_reset; // @[:@163569.4 RegFile.scala 76:16:@163576.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@163575.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@163579.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@163573.4]
  assign regs_128_clock = clock; // @[:@163582.4]
  assign regs_128_reset = io_reset; // @[:@163583.4 RegFile.scala 76:16:@163590.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@163589.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@163593.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@163587.4]
  assign regs_129_clock = clock; // @[:@163596.4]
  assign regs_129_reset = io_reset; // @[:@163597.4 RegFile.scala 76:16:@163604.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@163603.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@163607.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@163601.4]
  assign regs_130_clock = clock; // @[:@163610.4]
  assign regs_130_reset = io_reset; // @[:@163611.4 RegFile.scala 76:16:@163618.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@163617.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@163621.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@163615.4]
  assign regs_131_clock = clock; // @[:@163624.4]
  assign regs_131_reset = io_reset; // @[:@163625.4 RegFile.scala 76:16:@163632.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@163631.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@163635.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@163629.4]
  assign regs_132_clock = clock; // @[:@163638.4]
  assign regs_132_reset = io_reset; // @[:@163639.4 RegFile.scala 76:16:@163646.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@163645.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@163649.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@163643.4]
  assign regs_133_clock = clock; // @[:@163652.4]
  assign regs_133_reset = io_reset; // @[:@163653.4 RegFile.scala 76:16:@163660.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@163659.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@163663.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@163657.4]
  assign regs_134_clock = clock; // @[:@163666.4]
  assign regs_134_reset = io_reset; // @[:@163667.4 RegFile.scala 76:16:@163674.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@163673.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@163677.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@163671.4]
  assign regs_135_clock = clock; // @[:@163680.4]
  assign regs_135_reset = io_reset; // @[:@163681.4 RegFile.scala 76:16:@163688.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@163687.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@163691.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@163685.4]
  assign regs_136_clock = clock; // @[:@163694.4]
  assign regs_136_reset = io_reset; // @[:@163695.4 RegFile.scala 76:16:@163702.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@163701.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@163705.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@163699.4]
  assign regs_137_clock = clock; // @[:@163708.4]
  assign regs_137_reset = io_reset; // @[:@163709.4 RegFile.scala 76:16:@163716.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@163715.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@163719.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@163713.4]
  assign regs_138_clock = clock; // @[:@163722.4]
  assign regs_138_reset = io_reset; // @[:@163723.4 RegFile.scala 76:16:@163730.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@163729.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@163733.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@163727.4]
  assign regs_139_clock = clock; // @[:@163736.4]
  assign regs_139_reset = io_reset; // @[:@163737.4 RegFile.scala 76:16:@163744.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@163743.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@163747.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@163741.4]
  assign regs_140_clock = clock; // @[:@163750.4]
  assign regs_140_reset = io_reset; // @[:@163751.4 RegFile.scala 76:16:@163758.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@163757.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@163761.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@163755.4]
  assign regs_141_clock = clock; // @[:@163764.4]
  assign regs_141_reset = io_reset; // @[:@163765.4 RegFile.scala 76:16:@163772.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@163771.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@163775.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@163769.4]
  assign regs_142_clock = clock; // @[:@163778.4]
  assign regs_142_reset = io_reset; // @[:@163779.4 RegFile.scala 76:16:@163786.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@163785.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@163789.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@163783.4]
  assign regs_143_clock = clock; // @[:@163792.4]
  assign regs_143_reset = io_reset; // @[:@163793.4 RegFile.scala 76:16:@163800.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@163799.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@163803.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@163797.4]
  assign regs_144_clock = clock; // @[:@163806.4]
  assign regs_144_reset = io_reset; // @[:@163807.4 RegFile.scala 76:16:@163814.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@163813.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@163817.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@163811.4]
  assign regs_145_clock = clock; // @[:@163820.4]
  assign regs_145_reset = io_reset; // @[:@163821.4 RegFile.scala 76:16:@163828.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@163827.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@163831.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@163825.4]
  assign regs_146_clock = clock; // @[:@163834.4]
  assign regs_146_reset = io_reset; // @[:@163835.4 RegFile.scala 76:16:@163842.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@163841.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@163845.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@163839.4]
  assign regs_147_clock = clock; // @[:@163848.4]
  assign regs_147_reset = io_reset; // @[:@163849.4 RegFile.scala 76:16:@163856.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@163855.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@163859.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@163853.4]
  assign regs_148_clock = clock; // @[:@163862.4]
  assign regs_148_reset = io_reset; // @[:@163863.4 RegFile.scala 76:16:@163870.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@163869.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@163873.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@163867.4]
  assign regs_149_clock = clock; // @[:@163876.4]
  assign regs_149_reset = io_reset; // @[:@163877.4 RegFile.scala 76:16:@163884.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@163883.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@163887.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@163881.4]
  assign regs_150_clock = clock; // @[:@163890.4]
  assign regs_150_reset = io_reset; // @[:@163891.4 RegFile.scala 76:16:@163898.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@163897.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@163901.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@163895.4]
  assign regs_151_clock = clock; // @[:@163904.4]
  assign regs_151_reset = io_reset; // @[:@163905.4 RegFile.scala 76:16:@163912.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@163911.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@163915.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@163909.4]
  assign regs_152_clock = clock; // @[:@163918.4]
  assign regs_152_reset = io_reset; // @[:@163919.4 RegFile.scala 76:16:@163926.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@163925.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@163929.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@163923.4]
  assign regs_153_clock = clock; // @[:@163932.4]
  assign regs_153_reset = io_reset; // @[:@163933.4 RegFile.scala 76:16:@163940.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@163939.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@163943.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@163937.4]
  assign regs_154_clock = clock; // @[:@163946.4]
  assign regs_154_reset = io_reset; // @[:@163947.4 RegFile.scala 76:16:@163954.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@163953.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@163957.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@163951.4]
  assign regs_155_clock = clock; // @[:@163960.4]
  assign regs_155_reset = io_reset; // @[:@163961.4 RegFile.scala 76:16:@163968.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@163967.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@163971.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@163965.4]
  assign regs_156_clock = clock; // @[:@163974.4]
  assign regs_156_reset = io_reset; // @[:@163975.4 RegFile.scala 76:16:@163982.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@163981.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@163985.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@163979.4]
  assign regs_157_clock = clock; // @[:@163988.4]
  assign regs_157_reset = io_reset; // @[:@163989.4 RegFile.scala 76:16:@163996.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@163995.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@163999.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@163993.4]
  assign regs_158_clock = clock; // @[:@164002.4]
  assign regs_158_reset = io_reset; // @[:@164003.4 RegFile.scala 76:16:@164010.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@164009.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@164013.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@164007.4]
  assign regs_159_clock = clock; // @[:@164016.4]
  assign regs_159_reset = io_reset; // @[:@164017.4 RegFile.scala 76:16:@164024.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@164023.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@164027.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@164021.4]
  assign regs_160_clock = clock; // @[:@164030.4]
  assign regs_160_reset = io_reset; // @[:@164031.4 RegFile.scala 76:16:@164038.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@164037.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@164041.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@164035.4]
  assign regs_161_clock = clock; // @[:@164044.4]
  assign regs_161_reset = io_reset; // @[:@164045.4 RegFile.scala 76:16:@164052.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@164051.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@164055.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@164049.4]
  assign regs_162_clock = clock; // @[:@164058.4]
  assign regs_162_reset = io_reset; // @[:@164059.4 RegFile.scala 76:16:@164066.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@164065.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@164069.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@164063.4]
  assign regs_163_clock = clock; // @[:@164072.4]
  assign regs_163_reset = io_reset; // @[:@164073.4 RegFile.scala 76:16:@164080.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@164079.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@164083.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@164077.4]
  assign regs_164_clock = clock; // @[:@164086.4]
  assign regs_164_reset = io_reset; // @[:@164087.4 RegFile.scala 76:16:@164094.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@164093.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@164097.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@164091.4]
  assign regs_165_clock = clock; // @[:@164100.4]
  assign regs_165_reset = io_reset; // @[:@164101.4 RegFile.scala 76:16:@164108.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@164107.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@164111.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@164105.4]
  assign regs_166_clock = clock; // @[:@164114.4]
  assign regs_166_reset = io_reset; // @[:@164115.4 RegFile.scala 76:16:@164122.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@164121.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@164125.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@164119.4]
  assign regs_167_clock = clock; // @[:@164128.4]
  assign regs_167_reset = io_reset; // @[:@164129.4 RegFile.scala 76:16:@164136.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@164135.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@164139.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@164133.4]
  assign regs_168_clock = clock; // @[:@164142.4]
  assign regs_168_reset = io_reset; // @[:@164143.4 RegFile.scala 76:16:@164150.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@164149.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@164153.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@164147.4]
  assign regs_169_clock = clock; // @[:@164156.4]
  assign regs_169_reset = io_reset; // @[:@164157.4 RegFile.scala 76:16:@164164.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@164163.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@164167.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@164161.4]
  assign regs_170_clock = clock; // @[:@164170.4]
  assign regs_170_reset = io_reset; // @[:@164171.4 RegFile.scala 76:16:@164178.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@164177.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@164181.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@164175.4]
  assign regs_171_clock = clock; // @[:@164184.4]
  assign regs_171_reset = io_reset; // @[:@164185.4 RegFile.scala 76:16:@164192.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@164191.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@164195.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@164189.4]
  assign regs_172_clock = clock; // @[:@164198.4]
  assign regs_172_reset = io_reset; // @[:@164199.4 RegFile.scala 76:16:@164206.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@164205.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@164209.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@164203.4]
  assign regs_173_clock = clock; // @[:@164212.4]
  assign regs_173_reset = io_reset; // @[:@164213.4 RegFile.scala 76:16:@164220.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@164219.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@164223.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@164217.4]
  assign regs_174_clock = clock; // @[:@164226.4]
  assign regs_174_reset = io_reset; // @[:@164227.4 RegFile.scala 76:16:@164234.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@164233.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@164237.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@164231.4]
  assign regs_175_clock = clock; // @[:@164240.4]
  assign regs_175_reset = io_reset; // @[:@164241.4 RegFile.scala 76:16:@164248.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@164247.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@164251.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@164245.4]
  assign regs_176_clock = clock; // @[:@164254.4]
  assign regs_176_reset = io_reset; // @[:@164255.4 RegFile.scala 76:16:@164262.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@164261.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@164265.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@164259.4]
  assign regs_177_clock = clock; // @[:@164268.4]
  assign regs_177_reset = io_reset; // @[:@164269.4 RegFile.scala 76:16:@164276.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@164275.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@164279.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@164273.4]
  assign regs_178_clock = clock; // @[:@164282.4]
  assign regs_178_reset = io_reset; // @[:@164283.4 RegFile.scala 76:16:@164290.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@164289.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@164293.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@164287.4]
  assign regs_179_clock = clock; // @[:@164296.4]
  assign regs_179_reset = io_reset; // @[:@164297.4 RegFile.scala 76:16:@164304.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@164303.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@164307.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@164301.4]
  assign regs_180_clock = clock; // @[:@164310.4]
  assign regs_180_reset = io_reset; // @[:@164311.4 RegFile.scala 76:16:@164318.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@164317.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@164321.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@164315.4]
  assign regs_181_clock = clock; // @[:@164324.4]
  assign regs_181_reset = io_reset; // @[:@164325.4 RegFile.scala 76:16:@164332.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@164331.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@164335.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@164329.4]
  assign regs_182_clock = clock; // @[:@164338.4]
  assign regs_182_reset = io_reset; // @[:@164339.4 RegFile.scala 76:16:@164346.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@164345.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@164349.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@164343.4]
  assign regs_183_clock = clock; // @[:@164352.4]
  assign regs_183_reset = io_reset; // @[:@164353.4 RegFile.scala 76:16:@164360.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@164359.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@164363.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@164357.4]
  assign regs_184_clock = clock; // @[:@164366.4]
  assign regs_184_reset = io_reset; // @[:@164367.4 RegFile.scala 76:16:@164374.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@164373.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@164377.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@164371.4]
  assign regs_185_clock = clock; // @[:@164380.4]
  assign regs_185_reset = io_reset; // @[:@164381.4 RegFile.scala 76:16:@164388.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@164387.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@164391.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@164385.4]
  assign regs_186_clock = clock; // @[:@164394.4]
  assign regs_186_reset = io_reset; // @[:@164395.4 RegFile.scala 76:16:@164402.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@164401.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@164405.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@164399.4]
  assign regs_187_clock = clock; // @[:@164408.4]
  assign regs_187_reset = io_reset; // @[:@164409.4 RegFile.scala 76:16:@164416.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@164415.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@164419.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@164413.4]
  assign regs_188_clock = clock; // @[:@164422.4]
  assign regs_188_reset = io_reset; // @[:@164423.4 RegFile.scala 76:16:@164430.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@164429.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@164433.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@164427.4]
  assign regs_189_clock = clock; // @[:@164436.4]
  assign regs_189_reset = io_reset; // @[:@164437.4 RegFile.scala 76:16:@164444.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@164443.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@164447.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@164441.4]
  assign regs_190_clock = clock; // @[:@164450.4]
  assign regs_190_reset = io_reset; // @[:@164451.4 RegFile.scala 76:16:@164458.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@164457.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@164461.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@164455.4]
  assign regs_191_clock = clock; // @[:@164464.4]
  assign regs_191_reset = io_reset; // @[:@164465.4 RegFile.scala 76:16:@164472.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@164471.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@164475.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@164469.4]
  assign regs_192_clock = clock; // @[:@164478.4]
  assign regs_192_reset = io_reset; // @[:@164479.4 RegFile.scala 76:16:@164486.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@164485.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@164489.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@164483.4]
  assign regs_193_clock = clock; // @[:@164492.4]
  assign regs_193_reset = io_reset; // @[:@164493.4 RegFile.scala 76:16:@164500.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@164499.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@164503.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@164497.4]
  assign regs_194_clock = clock; // @[:@164506.4]
  assign regs_194_reset = io_reset; // @[:@164507.4 RegFile.scala 76:16:@164514.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@164513.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@164517.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@164511.4]
  assign regs_195_clock = clock; // @[:@164520.4]
  assign regs_195_reset = io_reset; // @[:@164521.4 RegFile.scala 76:16:@164528.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@164527.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@164531.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@164525.4]
  assign regs_196_clock = clock; // @[:@164534.4]
  assign regs_196_reset = io_reset; // @[:@164535.4 RegFile.scala 76:16:@164542.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@164541.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@164545.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@164539.4]
  assign regs_197_clock = clock; // @[:@164548.4]
  assign regs_197_reset = io_reset; // @[:@164549.4 RegFile.scala 76:16:@164556.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@164555.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@164559.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@164553.4]
  assign regs_198_clock = clock; // @[:@164562.4]
  assign regs_198_reset = io_reset; // @[:@164563.4 RegFile.scala 76:16:@164570.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@164569.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@164573.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@164567.4]
  assign regs_199_clock = clock; // @[:@164576.4]
  assign regs_199_reset = io_reset; // @[:@164577.4 RegFile.scala 76:16:@164584.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@164583.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@164587.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@164581.4]
  assign regs_200_clock = clock; // @[:@164590.4]
  assign regs_200_reset = io_reset; // @[:@164591.4 RegFile.scala 76:16:@164598.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@164597.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@164601.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@164595.4]
  assign regs_201_clock = clock; // @[:@164604.4]
  assign regs_201_reset = io_reset; // @[:@164605.4 RegFile.scala 76:16:@164612.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@164611.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@164615.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@164609.4]
  assign regs_202_clock = clock; // @[:@164618.4]
  assign regs_202_reset = io_reset; // @[:@164619.4 RegFile.scala 76:16:@164626.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@164625.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@164629.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@164623.4]
  assign regs_203_clock = clock; // @[:@164632.4]
  assign regs_203_reset = io_reset; // @[:@164633.4 RegFile.scala 76:16:@164640.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@164639.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@164643.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@164637.4]
  assign regs_204_clock = clock; // @[:@164646.4]
  assign regs_204_reset = io_reset; // @[:@164647.4 RegFile.scala 76:16:@164654.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@164653.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@164657.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@164651.4]
  assign regs_205_clock = clock; // @[:@164660.4]
  assign regs_205_reset = io_reset; // @[:@164661.4 RegFile.scala 76:16:@164668.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@164667.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@164671.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@164665.4]
  assign regs_206_clock = clock; // @[:@164674.4]
  assign regs_206_reset = io_reset; // @[:@164675.4 RegFile.scala 76:16:@164682.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@164681.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@164685.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@164679.4]
  assign regs_207_clock = clock; // @[:@164688.4]
  assign regs_207_reset = io_reset; // @[:@164689.4 RegFile.scala 76:16:@164696.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@164695.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@164699.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@164693.4]
  assign regs_208_clock = clock; // @[:@164702.4]
  assign regs_208_reset = io_reset; // @[:@164703.4 RegFile.scala 76:16:@164710.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@164709.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@164713.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@164707.4]
  assign regs_209_clock = clock; // @[:@164716.4]
  assign regs_209_reset = io_reset; // @[:@164717.4 RegFile.scala 76:16:@164724.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@164723.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@164727.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@164721.4]
  assign regs_210_clock = clock; // @[:@164730.4]
  assign regs_210_reset = io_reset; // @[:@164731.4 RegFile.scala 76:16:@164738.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@164737.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@164741.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@164735.4]
  assign regs_211_clock = clock; // @[:@164744.4]
  assign regs_211_reset = io_reset; // @[:@164745.4 RegFile.scala 76:16:@164752.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@164751.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@164755.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@164749.4]
  assign regs_212_clock = clock; // @[:@164758.4]
  assign regs_212_reset = io_reset; // @[:@164759.4 RegFile.scala 76:16:@164766.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@164765.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@164769.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@164763.4]
  assign regs_213_clock = clock; // @[:@164772.4]
  assign regs_213_reset = io_reset; // @[:@164773.4 RegFile.scala 76:16:@164780.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@164779.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@164783.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@164777.4]
  assign regs_214_clock = clock; // @[:@164786.4]
  assign regs_214_reset = io_reset; // @[:@164787.4 RegFile.scala 76:16:@164794.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@164793.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@164797.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@164791.4]
  assign regs_215_clock = clock; // @[:@164800.4]
  assign regs_215_reset = io_reset; // @[:@164801.4 RegFile.scala 76:16:@164808.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@164807.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@164811.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@164805.4]
  assign regs_216_clock = clock; // @[:@164814.4]
  assign regs_216_reset = io_reset; // @[:@164815.4 RegFile.scala 76:16:@164822.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@164821.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@164825.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@164819.4]
  assign regs_217_clock = clock; // @[:@164828.4]
  assign regs_217_reset = io_reset; // @[:@164829.4 RegFile.scala 76:16:@164836.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@164835.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@164839.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@164833.4]
  assign regs_218_clock = clock; // @[:@164842.4]
  assign regs_218_reset = io_reset; // @[:@164843.4 RegFile.scala 76:16:@164850.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@164849.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@164853.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@164847.4]
  assign regs_219_clock = clock; // @[:@164856.4]
  assign regs_219_reset = io_reset; // @[:@164857.4 RegFile.scala 76:16:@164864.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@164863.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@164867.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@164861.4]
  assign regs_220_clock = clock; // @[:@164870.4]
  assign regs_220_reset = io_reset; // @[:@164871.4 RegFile.scala 76:16:@164878.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@164877.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@164881.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@164875.4]
  assign regs_221_clock = clock; // @[:@164884.4]
  assign regs_221_reset = io_reset; // @[:@164885.4 RegFile.scala 76:16:@164892.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@164891.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@164895.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@164889.4]
  assign regs_222_clock = clock; // @[:@164898.4]
  assign regs_222_reset = io_reset; // @[:@164899.4 RegFile.scala 76:16:@164906.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@164905.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@164909.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@164903.4]
  assign regs_223_clock = clock; // @[:@164912.4]
  assign regs_223_reset = io_reset; // @[:@164913.4 RegFile.scala 76:16:@164920.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@164919.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@164923.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@164917.4]
  assign regs_224_clock = clock; // @[:@164926.4]
  assign regs_224_reset = io_reset; // @[:@164927.4 RegFile.scala 76:16:@164934.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@164933.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@164937.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@164931.4]
  assign regs_225_clock = clock; // @[:@164940.4]
  assign regs_225_reset = io_reset; // @[:@164941.4 RegFile.scala 76:16:@164948.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@164947.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@164951.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@164945.4]
  assign regs_226_clock = clock; // @[:@164954.4]
  assign regs_226_reset = io_reset; // @[:@164955.4 RegFile.scala 76:16:@164962.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@164961.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@164965.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@164959.4]
  assign regs_227_clock = clock; // @[:@164968.4]
  assign regs_227_reset = io_reset; // @[:@164969.4 RegFile.scala 76:16:@164976.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@164975.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@164979.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@164973.4]
  assign regs_228_clock = clock; // @[:@164982.4]
  assign regs_228_reset = io_reset; // @[:@164983.4 RegFile.scala 76:16:@164990.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@164989.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@164993.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@164987.4]
  assign regs_229_clock = clock; // @[:@164996.4]
  assign regs_229_reset = io_reset; // @[:@164997.4 RegFile.scala 76:16:@165004.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@165003.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@165007.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@165001.4]
  assign regs_230_clock = clock; // @[:@165010.4]
  assign regs_230_reset = io_reset; // @[:@165011.4 RegFile.scala 76:16:@165018.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@165017.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@165021.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@165015.4]
  assign regs_231_clock = clock; // @[:@165024.4]
  assign regs_231_reset = io_reset; // @[:@165025.4 RegFile.scala 76:16:@165032.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@165031.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@165035.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@165029.4]
  assign regs_232_clock = clock; // @[:@165038.4]
  assign regs_232_reset = io_reset; // @[:@165039.4 RegFile.scala 76:16:@165046.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@165045.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@165049.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@165043.4]
  assign regs_233_clock = clock; // @[:@165052.4]
  assign regs_233_reset = io_reset; // @[:@165053.4 RegFile.scala 76:16:@165060.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@165059.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@165063.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@165057.4]
  assign regs_234_clock = clock; // @[:@165066.4]
  assign regs_234_reset = io_reset; // @[:@165067.4 RegFile.scala 76:16:@165074.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@165073.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@165077.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@165071.4]
  assign regs_235_clock = clock; // @[:@165080.4]
  assign regs_235_reset = io_reset; // @[:@165081.4 RegFile.scala 76:16:@165088.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@165087.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@165091.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@165085.4]
  assign regs_236_clock = clock; // @[:@165094.4]
  assign regs_236_reset = io_reset; // @[:@165095.4 RegFile.scala 76:16:@165102.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@165101.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@165105.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@165099.4]
  assign regs_237_clock = clock; // @[:@165108.4]
  assign regs_237_reset = io_reset; // @[:@165109.4 RegFile.scala 76:16:@165116.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@165115.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@165119.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@165113.4]
  assign regs_238_clock = clock; // @[:@165122.4]
  assign regs_238_reset = io_reset; // @[:@165123.4 RegFile.scala 76:16:@165130.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@165129.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@165133.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@165127.4]
  assign regs_239_clock = clock; // @[:@165136.4]
  assign regs_239_reset = io_reset; // @[:@165137.4 RegFile.scala 76:16:@165144.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@165143.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@165147.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@165141.4]
  assign regs_240_clock = clock; // @[:@165150.4]
  assign regs_240_reset = io_reset; // @[:@165151.4 RegFile.scala 76:16:@165158.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@165157.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@165161.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@165155.4]
  assign regs_241_clock = clock; // @[:@165164.4]
  assign regs_241_reset = io_reset; // @[:@165165.4 RegFile.scala 76:16:@165172.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@165171.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@165175.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@165169.4]
  assign regs_242_clock = clock; // @[:@165178.4]
  assign regs_242_reset = io_reset; // @[:@165179.4 RegFile.scala 76:16:@165186.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@165185.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@165189.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@165183.4]
  assign regs_243_clock = clock; // @[:@165192.4]
  assign regs_243_reset = io_reset; // @[:@165193.4 RegFile.scala 76:16:@165200.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@165199.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@165203.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@165197.4]
  assign regs_244_clock = clock; // @[:@165206.4]
  assign regs_244_reset = io_reset; // @[:@165207.4 RegFile.scala 76:16:@165214.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@165213.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@165217.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@165211.4]
  assign regs_245_clock = clock; // @[:@165220.4]
  assign regs_245_reset = io_reset; // @[:@165221.4 RegFile.scala 76:16:@165228.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@165227.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@165231.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@165225.4]
  assign regs_246_clock = clock; // @[:@165234.4]
  assign regs_246_reset = io_reset; // @[:@165235.4 RegFile.scala 76:16:@165242.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@165241.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@165245.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@165239.4]
  assign regs_247_clock = clock; // @[:@165248.4]
  assign regs_247_reset = io_reset; // @[:@165249.4 RegFile.scala 76:16:@165256.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@165255.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@165259.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@165253.4]
  assign regs_248_clock = clock; // @[:@165262.4]
  assign regs_248_reset = io_reset; // @[:@165263.4 RegFile.scala 76:16:@165270.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@165269.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@165273.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@165267.4]
  assign regs_249_clock = clock; // @[:@165276.4]
  assign regs_249_reset = io_reset; // @[:@165277.4 RegFile.scala 76:16:@165284.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@165283.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@165287.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@165281.4]
  assign regs_250_clock = clock; // @[:@165290.4]
  assign regs_250_reset = io_reset; // @[:@165291.4 RegFile.scala 76:16:@165298.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@165297.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@165301.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@165295.4]
  assign regs_251_clock = clock; // @[:@165304.4]
  assign regs_251_reset = io_reset; // @[:@165305.4 RegFile.scala 76:16:@165312.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@165311.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@165315.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@165309.4]
  assign regs_252_clock = clock; // @[:@165318.4]
  assign regs_252_reset = io_reset; // @[:@165319.4 RegFile.scala 76:16:@165326.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@165325.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@165329.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@165323.4]
  assign regs_253_clock = clock; // @[:@165332.4]
  assign regs_253_reset = io_reset; // @[:@165333.4 RegFile.scala 76:16:@165340.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@165339.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@165343.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@165337.4]
  assign regs_254_clock = clock; // @[:@165346.4]
  assign regs_254_reset = io_reset; // @[:@165347.4 RegFile.scala 76:16:@165354.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@165353.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@165357.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@165351.4]
  assign regs_255_clock = clock; // @[:@165360.4]
  assign regs_255_reset = io_reset; // @[:@165361.4 RegFile.scala 76:16:@165368.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@165367.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@165371.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@165365.4]
  assign regs_256_clock = clock; // @[:@165374.4]
  assign regs_256_reset = io_reset; // @[:@165375.4 RegFile.scala 76:16:@165382.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@165381.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@165385.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@165379.4]
  assign regs_257_clock = clock; // @[:@165388.4]
  assign regs_257_reset = io_reset; // @[:@165389.4 RegFile.scala 76:16:@165396.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@165395.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@165399.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@165393.4]
  assign regs_258_clock = clock; // @[:@165402.4]
  assign regs_258_reset = io_reset; // @[:@165403.4 RegFile.scala 76:16:@165410.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@165409.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@165413.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@165407.4]
  assign regs_259_clock = clock; // @[:@165416.4]
  assign regs_259_reset = io_reset; // @[:@165417.4 RegFile.scala 76:16:@165424.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@165423.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@165427.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@165421.4]
  assign regs_260_clock = clock; // @[:@165430.4]
  assign regs_260_reset = io_reset; // @[:@165431.4 RegFile.scala 76:16:@165438.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@165437.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@165441.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@165435.4]
  assign regs_261_clock = clock; // @[:@165444.4]
  assign regs_261_reset = io_reset; // @[:@165445.4 RegFile.scala 76:16:@165452.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@165451.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@165455.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@165449.4]
  assign regs_262_clock = clock; // @[:@165458.4]
  assign regs_262_reset = io_reset; // @[:@165459.4 RegFile.scala 76:16:@165466.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@165465.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@165469.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@165463.4]
  assign regs_263_clock = clock; // @[:@165472.4]
  assign regs_263_reset = io_reset; // @[:@165473.4 RegFile.scala 76:16:@165480.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@165479.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@165483.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@165477.4]
  assign regs_264_clock = clock; // @[:@165486.4]
  assign regs_264_reset = io_reset; // @[:@165487.4 RegFile.scala 76:16:@165494.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@165493.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@165497.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@165491.4]
  assign regs_265_clock = clock; // @[:@165500.4]
  assign regs_265_reset = io_reset; // @[:@165501.4 RegFile.scala 76:16:@165508.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@165507.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@165511.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@165505.4]
  assign regs_266_clock = clock; // @[:@165514.4]
  assign regs_266_reset = io_reset; // @[:@165515.4 RegFile.scala 76:16:@165522.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@165521.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@165525.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@165519.4]
  assign regs_267_clock = clock; // @[:@165528.4]
  assign regs_267_reset = io_reset; // @[:@165529.4 RegFile.scala 76:16:@165536.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@165535.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@165539.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@165533.4]
  assign regs_268_clock = clock; // @[:@165542.4]
  assign regs_268_reset = io_reset; // @[:@165543.4 RegFile.scala 76:16:@165550.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@165549.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@165553.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@165547.4]
  assign regs_269_clock = clock; // @[:@165556.4]
  assign regs_269_reset = io_reset; // @[:@165557.4 RegFile.scala 76:16:@165564.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@165563.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@165567.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@165561.4]
  assign regs_270_clock = clock; // @[:@165570.4]
  assign regs_270_reset = io_reset; // @[:@165571.4 RegFile.scala 76:16:@165578.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@165577.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@165581.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@165575.4]
  assign regs_271_clock = clock; // @[:@165584.4]
  assign regs_271_reset = io_reset; // @[:@165585.4 RegFile.scala 76:16:@165592.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@165591.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@165595.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@165589.4]
  assign regs_272_clock = clock; // @[:@165598.4]
  assign regs_272_reset = io_reset; // @[:@165599.4 RegFile.scala 76:16:@165606.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@165605.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@165609.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@165603.4]
  assign regs_273_clock = clock; // @[:@165612.4]
  assign regs_273_reset = io_reset; // @[:@165613.4 RegFile.scala 76:16:@165620.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@165619.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@165623.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@165617.4]
  assign regs_274_clock = clock; // @[:@165626.4]
  assign regs_274_reset = io_reset; // @[:@165627.4 RegFile.scala 76:16:@165634.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@165633.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@165637.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@165631.4]
  assign regs_275_clock = clock; // @[:@165640.4]
  assign regs_275_reset = io_reset; // @[:@165641.4 RegFile.scala 76:16:@165648.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@165647.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@165651.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@165645.4]
  assign regs_276_clock = clock; // @[:@165654.4]
  assign regs_276_reset = io_reset; // @[:@165655.4 RegFile.scala 76:16:@165662.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@165661.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@165665.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@165659.4]
  assign regs_277_clock = clock; // @[:@165668.4]
  assign regs_277_reset = io_reset; // @[:@165669.4 RegFile.scala 76:16:@165676.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@165675.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@165679.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@165673.4]
  assign regs_278_clock = clock; // @[:@165682.4]
  assign regs_278_reset = io_reset; // @[:@165683.4 RegFile.scala 76:16:@165690.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@165689.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@165693.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@165687.4]
  assign regs_279_clock = clock; // @[:@165696.4]
  assign regs_279_reset = io_reset; // @[:@165697.4 RegFile.scala 76:16:@165704.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@165703.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@165707.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@165701.4]
  assign regs_280_clock = clock; // @[:@165710.4]
  assign regs_280_reset = io_reset; // @[:@165711.4 RegFile.scala 76:16:@165718.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@165717.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@165721.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@165715.4]
  assign regs_281_clock = clock; // @[:@165724.4]
  assign regs_281_reset = io_reset; // @[:@165725.4 RegFile.scala 76:16:@165732.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@165731.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@165735.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@165729.4]
  assign regs_282_clock = clock; // @[:@165738.4]
  assign regs_282_reset = io_reset; // @[:@165739.4 RegFile.scala 76:16:@165746.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@165745.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@165749.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@165743.4]
  assign regs_283_clock = clock; // @[:@165752.4]
  assign regs_283_reset = io_reset; // @[:@165753.4 RegFile.scala 76:16:@165760.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@165759.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@165763.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@165757.4]
  assign regs_284_clock = clock; // @[:@165766.4]
  assign regs_284_reset = io_reset; // @[:@165767.4 RegFile.scala 76:16:@165774.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@165773.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@165777.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@165771.4]
  assign regs_285_clock = clock; // @[:@165780.4]
  assign regs_285_reset = io_reset; // @[:@165781.4 RegFile.scala 76:16:@165788.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@165787.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@165791.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@165785.4]
  assign regs_286_clock = clock; // @[:@165794.4]
  assign regs_286_reset = io_reset; // @[:@165795.4 RegFile.scala 76:16:@165802.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@165801.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@165805.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@165799.4]
  assign regs_287_clock = clock; // @[:@165808.4]
  assign regs_287_reset = io_reset; // @[:@165809.4 RegFile.scala 76:16:@165816.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@165815.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@165819.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@165813.4]
  assign regs_288_clock = clock; // @[:@165822.4]
  assign regs_288_reset = io_reset; // @[:@165823.4 RegFile.scala 76:16:@165830.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@165829.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@165833.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@165827.4]
  assign regs_289_clock = clock; // @[:@165836.4]
  assign regs_289_reset = io_reset; // @[:@165837.4 RegFile.scala 76:16:@165844.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@165843.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@165847.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@165841.4]
  assign regs_290_clock = clock; // @[:@165850.4]
  assign regs_290_reset = io_reset; // @[:@165851.4 RegFile.scala 76:16:@165858.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@165857.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@165861.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@165855.4]
  assign regs_291_clock = clock; // @[:@165864.4]
  assign regs_291_reset = io_reset; // @[:@165865.4 RegFile.scala 76:16:@165872.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@165871.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@165875.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@165869.4]
  assign regs_292_clock = clock; // @[:@165878.4]
  assign regs_292_reset = io_reset; // @[:@165879.4 RegFile.scala 76:16:@165886.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@165885.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@165889.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@165883.4]
  assign regs_293_clock = clock; // @[:@165892.4]
  assign regs_293_reset = io_reset; // @[:@165893.4 RegFile.scala 76:16:@165900.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@165899.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@165903.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@165897.4]
  assign regs_294_clock = clock; // @[:@165906.4]
  assign regs_294_reset = io_reset; // @[:@165907.4 RegFile.scala 76:16:@165914.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@165913.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@165917.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@165911.4]
  assign regs_295_clock = clock; // @[:@165920.4]
  assign regs_295_reset = io_reset; // @[:@165921.4 RegFile.scala 76:16:@165928.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@165927.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@165931.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@165925.4]
  assign regs_296_clock = clock; // @[:@165934.4]
  assign regs_296_reset = io_reset; // @[:@165935.4 RegFile.scala 76:16:@165942.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@165941.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@165945.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@165939.4]
  assign regs_297_clock = clock; // @[:@165948.4]
  assign regs_297_reset = io_reset; // @[:@165949.4 RegFile.scala 76:16:@165956.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@165955.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@165959.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@165953.4]
  assign regs_298_clock = clock; // @[:@165962.4]
  assign regs_298_reset = io_reset; // @[:@165963.4 RegFile.scala 76:16:@165970.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@165969.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@165973.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@165967.4]
  assign regs_299_clock = clock; // @[:@165976.4]
  assign regs_299_reset = io_reset; // @[:@165977.4 RegFile.scala 76:16:@165984.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@165983.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@165987.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@165981.4]
  assign regs_300_clock = clock; // @[:@165990.4]
  assign regs_300_reset = io_reset; // @[:@165991.4 RegFile.scala 76:16:@165998.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@165997.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@166001.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@165995.4]
  assign regs_301_clock = clock; // @[:@166004.4]
  assign regs_301_reset = io_reset; // @[:@166005.4 RegFile.scala 76:16:@166012.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@166011.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@166015.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@166009.4]
  assign regs_302_clock = clock; // @[:@166018.4]
  assign regs_302_reset = io_reset; // @[:@166019.4 RegFile.scala 76:16:@166026.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@166025.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@166029.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@166023.4]
  assign regs_303_clock = clock; // @[:@166032.4]
  assign regs_303_reset = io_reset; // @[:@166033.4 RegFile.scala 76:16:@166040.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@166039.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@166043.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@166037.4]
  assign regs_304_clock = clock; // @[:@166046.4]
  assign regs_304_reset = io_reset; // @[:@166047.4 RegFile.scala 76:16:@166054.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@166053.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@166057.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@166051.4]
  assign regs_305_clock = clock; // @[:@166060.4]
  assign regs_305_reset = io_reset; // @[:@166061.4 RegFile.scala 76:16:@166068.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@166067.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@166071.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@166065.4]
  assign regs_306_clock = clock; // @[:@166074.4]
  assign regs_306_reset = io_reset; // @[:@166075.4 RegFile.scala 76:16:@166082.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@166081.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@166085.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@166079.4]
  assign regs_307_clock = clock; // @[:@166088.4]
  assign regs_307_reset = io_reset; // @[:@166089.4 RegFile.scala 76:16:@166096.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@166095.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@166099.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@166093.4]
  assign regs_308_clock = clock; // @[:@166102.4]
  assign regs_308_reset = io_reset; // @[:@166103.4 RegFile.scala 76:16:@166110.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@166109.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@166113.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@166107.4]
  assign regs_309_clock = clock; // @[:@166116.4]
  assign regs_309_reset = io_reset; // @[:@166117.4 RegFile.scala 76:16:@166124.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@166123.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@166127.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@166121.4]
  assign regs_310_clock = clock; // @[:@166130.4]
  assign regs_310_reset = io_reset; // @[:@166131.4 RegFile.scala 76:16:@166138.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@166137.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@166141.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@166135.4]
  assign regs_311_clock = clock; // @[:@166144.4]
  assign regs_311_reset = io_reset; // @[:@166145.4 RegFile.scala 76:16:@166152.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@166151.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@166155.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@166149.4]
  assign regs_312_clock = clock; // @[:@166158.4]
  assign regs_312_reset = io_reset; // @[:@166159.4 RegFile.scala 76:16:@166166.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@166165.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@166169.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@166163.4]
  assign regs_313_clock = clock; // @[:@166172.4]
  assign regs_313_reset = io_reset; // @[:@166173.4 RegFile.scala 76:16:@166180.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@166179.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@166183.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@166177.4]
  assign regs_314_clock = clock; // @[:@166186.4]
  assign regs_314_reset = io_reset; // @[:@166187.4 RegFile.scala 76:16:@166194.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@166193.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@166197.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@166191.4]
  assign regs_315_clock = clock; // @[:@166200.4]
  assign regs_315_reset = io_reset; // @[:@166201.4 RegFile.scala 76:16:@166208.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@166207.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@166211.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@166205.4]
  assign regs_316_clock = clock; // @[:@166214.4]
  assign regs_316_reset = io_reset; // @[:@166215.4 RegFile.scala 76:16:@166222.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@166221.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@166225.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@166219.4]
  assign regs_317_clock = clock; // @[:@166228.4]
  assign regs_317_reset = io_reset; // @[:@166229.4 RegFile.scala 76:16:@166236.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@166235.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@166239.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@166233.4]
  assign regs_318_clock = clock; // @[:@166242.4]
  assign regs_318_reset = io_reset; // @[:@166243.4 RegFile.scala 76:16:@166250.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@166249.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@166253.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@166247.4]
  assign regs_319_clock = clock; // @[:@166256.4]
  assign regs_319_reset = io_reset; // @[:@166257.4 RegFile.scala 76:16:@166264.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@166263.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@166267.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@166261.4]
  assign regs_320_clock = clock; // @[:@166270.4]
  assign regs_320_reset = io_reset; // @[:@166271.4 RegFile.scala 76:16:@166278.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@166277.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@166281.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@166275.4]
  assign regs_321_clock = clock; // @[:@166284.4]
  assign regs_321_reset = io_reset; // @[:@166285.4 RegFile.scala 76:16:@166292.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@166291.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@166295.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@166289.4]
  assign regs_322_clock = clock; // @[:@166298.4]
  assign regs_322_reset = io_reset; // @[:@166299.4 RegFile.scala 76:16:@166306.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@166305.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@166309.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@166303.4]
  assign regs_323_clock = clock; // @[:@166312.4]
  assign regs_323_reset = io_reset; // @[:@166313.4 RegFile.scala 76:16:@166320.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@166319.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@166323.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@166317.4]
  assign regs_324_clock = clock; // @[:@166326.4]
  assign regs_324_reset = io_reset; // @[:@166327.4 RegFile.scala 76:16:@166334.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@166333.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@166337.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@166331.4]
  assign regs_325_clock = clock; // @[:@166340.4]
  assign regs_325_reset = io_reset; // @[:@166341.4 RegFile.scala 76:16:@166348.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@166347.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@166351.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@166345.4]
  assign regs_326_clock = clock; // @[:@166354.4]
  assign regs_326_reset = io_reset; // @[:@166355.4 RegFile.scala 76:16:@166362.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@166361.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@166365.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@166359.4]
  assign regs_327_clock = clock; // @[:@166368.4]
  assign regs_327_reset = io_reset; // @[:@166369.4 RegFile.scala 76:16:@166376.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@166375.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@166379.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@166373.4]
  assign regs_328_clock = clock; // @[:@166382.4]
  assign regs_328_reset = io_reset; // @[:@166383.4 RegFile.scala 76:16:@166390.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@166389.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@166393.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@166387.4]
  assign regs_329_clock = clock; // @[:@166396.4]
  assign regs_329_reset = io_reset; // @[:@166397.4 RegFile.scala 76:16:@166404.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@166403.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@166407.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@166401.4]
  assign regs_330_clock = clock; // @[:@166410.4]
  assign regs_330_reset = io_reset; // @[:@166411.4 RegFile.scala 76:16:@166418.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@166417.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@166421.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@166415.4]
  assign regs_331_clock = clock; // @[:@166424.4]
  assign regs_331_reset = io_reset; // @[:@166425.4 RegFile.scala 76:16:@166432.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@166431.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@166435.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@166429.4]
  assign regs_332_clock = clock; // @[:@166438.4]
  assign regs_332_reset = io_reset; // @[:@166439.4 RegFile.scala 76:16:@166446.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@166445.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@166449.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@166443.4]
  assign regs_333_clock = clock; // @[:@166452.4]
  assign regs_333_reset = io_reset; // @[:@166453.4 RegFile.scala 76:16:@166460.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@166459.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@166463.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@166457.4]
  assign regs_334_clock = clock; // @[:@166466.4]
  assign regs_334_reset = io_reset; // @[:@166467.4 RegFile.scala 76:16:@166474.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@166473.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@166477.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@166471.4]
  assign regs_335_clock = clock; // @[:@166480.4]
  assign regs_335_reset = io_reset; // @[:@166481.4 RegFile.scala 76:16:@166488.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@166487.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@166491.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@166485.4]
  assign regs_336_clock = clock; // @[:@166494.4]
  assign regs_336_reset = io_reset; // @[:@166495.4 RegFile.scala 76:16:@166502.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@166501.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@166505.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@166499.4]
  assign regs_337_clock = clock; // @[:@166508.4]
  assign regs_337_reset = io_reset; // @[:@166509.4 RegFile.scala 76:16:@166516.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@166515.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@166519.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@166513.4]
  assign regs_338_clock = clock; // @[:@166522.4]
  assign regs_338_reset = io_reset; // @[:@166523.4 RegFile.scala 76:16:@166530.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@166529.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@166533.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@166527.4]
  assign regs_339_clock = clock; // @[:@166536.4]
  assign regs_339_reset = io_reset; // @[:@166537.4 RegFile.scala 76:16:@166544.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@166543.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@166547.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@166541.4]
  assign regs_340_clock = clock; // @[:@166550.4]
  assign regs_340_reset = io_reset; // @[:@166551.4 RegFile.scala 76:16:@166558.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@166557.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@166561.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@166555.4]
  assign regs_341_clock = clock; // @[:@166564.4]
  assign regs_341_reset = io_reset; // @[:@166565.4 RegFile.scala 76:16:@166572.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@166571.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@166575.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@166569.4]
  assign regs_342_clock = clock; // @[:@166578.4]
  assign regs_342_reset = io_reset; // @[:@166579.4 RegFile.scala 76:16:@166586.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@166585.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@166589.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@166583.4]
  assign regs_343_clock = clock; // @[:@166592.4]
  assign regs_343_reset = io_reset; // @[:@166593.4 RegFile.scala 76:16:@166600.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@166599.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@166603.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@166597.4]
  assign regs_344_clock = clock; // @[:@166606.4]
  assign regs_344_reset = io_reset; // @[:@166607.4 RegFile.scala 76:16:@166614.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@166613.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@166617.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@166611.4]
  assign regs_345_clock = clock; // @[:@166620.4]
  assign regs_345_reset = io_reset; // @[:@166621.4 RegFile.scala 76:16:@166628.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@166627.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@166631.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@166625.4]
  assign regs_346_clock = clock; // @[:@166634.4]
  assign regs_346_reset = io_reset; // @[:@166635.4 RegFile.scala 76:16:@166642.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@166641.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@166645.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@166639.4]
  assign regs_347_clock = clock; // @[:@166648.4]
  assign regs_347_reset = io_reset; // @[:@166649.4 RegFile.scala 76:16:@166656.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@166655.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@166659.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@166653.4]
  assign regs_348_clock = clock; // @[:@166662.4]
  assign regs_348_reset = io_reset; // @[:@166663.4 RegFile.scala 76:16:@166670.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@166669.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@166673.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@166667.4]
  assign regs_349_clock = clock; // @[:@166676.4]
  assign regs_349_reset = io_reset; // @[:@166677.4 RegFile.scala 76:16:@166684.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@166683.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@166687.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@166681.4]
  assign regs_350_clock = clock; // @[:@166690.4]
  assign regs_350_reset = io_reset; // @[:@166691.4 RegFile.scala 76:16:@166698.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@166697.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@166701.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@166695.4]
  assign regs_351_clock = clock; // @[:@166704.4]
  assign regs_351_reset = io_reset; // @[:@166705.4 RegFile.scala 76:16:@166712.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@166711.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@166715.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@166709.4]
  assign regs_352_clock = clock; // @[:@166718.4]
  assign regs_352_reset = io_reset; // @[:@166719.4 RegFile.scala 76:16:@166726.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@166725.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@166729.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@166723.4]
  assign regs_353_clock = clock; // @[:@166732.4]
  assign regs_353_reset = io_reset; // @[:@166733.4 RegFile.scala 76:16:@166740.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@166739.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@166743.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@166737.4]
  assign regs_354_clock = clock; // @[:@166746.4]
  assign regs_354_reset = io_reset; // @[:@166747.4 RegFile.scala 76:16:@166754.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@166753.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@166757.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@166751.4]
  assign regs_355_clock = clock; // @[:@166760.4]
  assign regs_355_reset = io_reset; // @[:@166761.4 RegFile.scala 76:16:@166768.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@166767.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@166771.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@166765.4]
  assign regs_356_clock = clock; // @[:@166774.4]
  assign regs_356_reset = io_reset; // @[:@166775.4 RegFile.scala 76:16:@166782.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@166781.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@166785.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@166779.4]
  assign regs_357_clock = clock; // @[:@166788.4]
  assign regs_357_reset = io_reset; // @[:@166789.4 RegFile.scala 76:16:@166796.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@166795.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@166799.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@166793.4]
  assign regs_358_clock = clock; // @[:@166802.4]
  assign regs_358_reset = io_reset; // @[:@166803.4 RegFile.scala 76:16:@166810.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@166809.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@166813.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@166807.4]
  assign regs_359_clock = clock; // @[:@166816.4]
  assign regs_359_reset = io_reset; // @[:@166817.4 RegFile.scala 76:16:@166824.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@166823.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@166827.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@166821.4]
  assign regs_360_clock = clock; // @[:@166830.4]
  assign regs_360_reset = io_reset; // @[:@166831.4 RegFile.scala 76:16:@166838.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@166837.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@166841.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@166835.4]
  assign regs_361_clock = clock; // @[:@166844.4]
  assign regs_361_reset = io_reset; // @[:@166845.4 RegFile.scala 76:16:@166852.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@166851.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@166855.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@166849.4]
  assign regs_362_clock = clock; // @[:@166858.4]
  assign regs_362_reset = io_reset; // @[:@166859.4 RegFile.scala 76:16:@166866.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@166865.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@166869.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@166863.4]
  assign regs_363_clock = clock; // @[:@166872.4]
  assign regs_363_reset = io_reset; // @[:@166873.4 RegFile.scala 76:16:@166880.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@166879.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@166883.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@166877.4]
  assign regs_364_clock = clock; // @[:@166886.4]
  assign regs_364_reset = io_reset; // @[:@166887.4 RegFile.scala 76:16:@166894.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@166893.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@166897.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@166891.4]
  assign regs_365_clock = clock; // @[:@166900.4]
  assign regs_365_reset = io_reset; // @[:@166901.4 RegFile.scala 76:16:@166908.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@166907.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@166911.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@166905.4]
  assign regs_366_clock = clock; // @[:@166914.4]
  assign regs_366_reset = io_reset; // @[:@166915.4 RegFile.scala 76:16:@166922.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@166921.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@166925.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@166919.4]
  assign regs_367_clock = clock; // @[:@166928.4]
  assign regs_367_reset = io_reset; // @[:@166929.4 RegFile.scala 76:16:@166936.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@166935.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@166939.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@166933.4]
  assign regs_368_clock = clock; // @[:@166942.4]
  assign regs_368_reset = io_reset; // @[:@166943.4 RegFile.scala 76:16:@166950.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@166949.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@166953.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@166947.4]
  assign regs_369_clock = clock; // @[:@166956.4]
  assign regs_369_reset = io_reset; // @[:@166957.4 RegFile.scala 76:16:@166964.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@166963.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@166967.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@166961.4]
  assign regs_370_clock = clock; // @[:@166970.4]
  assign regs_370_reset = io_reset; // @[:@166971.4 RegFile.scala 76:16:@166978.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@166977.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@166981.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@166975.4]
  assign regs_371_clock = clock; // @[:@166984.4]
  assign regs_371_reset = io_reset; // @[:@166985.4 RegFile.scala 76:16:@166992.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@166991.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@166995.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@166989.4]
  assign regs_372_clock = clock; // @[:@166998.4]
  assign regs_372_reset = io_reset; // @[:@166999.4 RegFile.scala 76:16:@167006.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@167005.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@167009.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@167003.4]
  assign regs_373_clock = clock; // @[:@167012.4]
  assign regs_373_reset = io_reset; // @[:@167013.4 RegFile.scala 76:16:@167020.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@167019.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@167023.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@167017.4]
  assign regs_374_clock = clock; // @[:@167026.4]
  assign regs_374_reset = io_reset; // @[:@167027.4 RegFile.scala 76:16:@167034.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@167033.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@167037.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@167031.4]
  assign regs_375_clock = clock; // @[:@167040.4]
  assign regs_375_reset = io_reset; // @[:@167041.4 RegFile.scala 76:16:@167048.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@167047.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@167051.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@167045.4]
  assign regs_376_clock = clock; // @[:@167054.4]
  assign regs_376_reset = io_reset; // @[:@167055.4 RegFile.scala 76:16:@167062.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@167061.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@167065.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@167059.4]
  assign regs_377_clock = clock; // @[:@167068.4]
  assign regs_377_reset = io_reset; // @[:@167069.4 RegFile.scala 76:16:@167076.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@167075.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@167079.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@167073.4]
  assign regs_378_clock = clock; // @[:@167082.4]
  assign regs_378_reset = io_reset; // @[:@167083.4 RegFile.scala 76:16:@167090.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@167089.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@167093.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@167087.4]
  assign regs_379_clock = clock; // @[:@167096.4]
  assign regs_379_reset = io_reset; // @[:@167097.4 RegFile.scala 76:16:@167104.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@167103.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@167107.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@167101.4]
  assign regs_380_clock = clock; // @[:@167110.4]
  assign regs_380_reset = io_reset; // @[:@167111.4 RegFile.scala 76:16:@167118.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@167117.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@167121.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@167115.4]
  assign regs_381_clock = clock; // @[:@167124.4]
  assign regs_381_reset = io_reset; // @[:@167125.4 RegFile.scala 76:16:@167132.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@167131.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@167135.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@167129.4]
  assign regs_382_clock = clock; // @[:@167138.4]
  assign regs_382_reset = io_reset; // @[:@167139.4 RegFile.scala 76:16:@167146.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@167145.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@167149.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@167143.4]
  assign regs_383_clock = clock; // @[:@167152.4]
  assign regs_383_reset = io_reset; // @[:@167153.4 RegFile.scala 76:16:@167160.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@167159.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@167163.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@167157.4]
  assign regs_384_clock = clock; // @[:@167166.4]
  assign regs_384_reset = io_reset; // @[:@167167.4 RegFile.scala 76:16:@167174.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@167173.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@167177.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@167171.4]
  assign regs_385_clock = clock; // @[:@167180.4]
  assign regs_385_reset = io_reset; // @[:@167181.4 RegFile.scala 76:16:@167188.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@167187.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@167191.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@167185.4]
  assign regs_386_clock = clock; // @[:@167194.4]
  assign regs_386_reset = io_reset; // @[:@167195.4 RegFile.scala 76:16:@167202.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@167201.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@167205.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@167199.4]
  assign regs_387_clock = clock; // @[:@167208.4]
  assign regs_387_reset = io_reset; // @[:@167209.4 RegFile.scala 76:16:@167216.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@167215.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@167219.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@167213.4]
  assign regs_388_clock = clock; // @[:@167222.4]
  assign regs_388_reset = io_reset; // @[:@167223.4 RegFile.scala 76:16:@167230.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@167229.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@167233.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@167227.4]
  assign regs_389_clock = clock; // @[:@167236.4]
  assign regs_389_reset = io_reset; // @[:@167237.4 RegFile.scala 76:16:@167244.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@167243.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@167247.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@167241.4]
  assign regs_390_clock = clock; // @[:@167250.4]
  assign regs_390_reset = io_reset; // @[:@167251.4 RegFile.scala 76:16:@167258.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@167257.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@167261.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@167255.4]
  assign regs_391_clock = clock; // @[:@167264.4]
  assign regs_391_reset = io_reset; // @[:@167265.4 RegFile.scala 76:16:@167272.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@167271.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@167275.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@167269.4]
  assign regs_392_clock = clock; // @[:@167278.4]
  assign regs_392_reset = io_reset; // @[:@167279.4 RegFile.scala 76:16:@167286.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@167285.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@167289.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@167283.4]
  assign regs_393_clock = clock; // @[:@167292.4]
  assign regs_393_reset = io_reset; // @[:@167293.4 RegFile.scala 76:16:@167300.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@167299.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@167303.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@167297.4]
  assign regs_394_clock = clock; // @[:@167306.4]
  assign regs_394_reset = io_reset; // @[:@167307.4 RegFile.scala 76:16:@167314.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@167313.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@167317.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@167311.4]
  assign regs_395_clock = clock; // @[:@167320.4]
  assign regs_395_reset = io_reset; // @[:@167321.4 RegFile.scala 76:16:@167328.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@167327.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@167331.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@167325.4]
  assign regs_396_clock = clock; // @[:@167334.4]
  assign regs_396_reset = io_reset; // @[:@167335.4 RegFile.scala 76:16:@167342.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@167341.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@167345.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@167339.4]
  assign regs_397_clock = clock; // @[:@167348.4]
  assign regs_397_reset = io_reset; // @[:@167349.4 RegFile.scala 76:16:@167356.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@167355.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@167359.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@167353.4]
  assign regs_398_clock = clock; // @[:@167362.4]
  assign regs_398_reset = io_reset; // @[:@167363.4 RegFile.scala 76:16:@167370.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@167369.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@167373.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@167367.4]
  assign regs_399_clock = clock; // @[:@167376.4]
  assign regs_399_reset = io_reset; // @[:@167377.4 RegFile.scala 76:16:@167384.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@167383.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@167387.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@167381.4]
  assign regs_400_clock = clock; // @[:@167390.4]
  assign regs_400_reset = io_reset; // @[:@167391.4 RegFile.scala 76:16:@167398.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@167397.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@167401.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@167395.4]
  assign regs_401_clock = clock; // @[:@167404.4]
  assign regs_401_reset = io_reset; // @[:@167405.4 RegFile.scala 76:16:@167412.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@167411.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@167415.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@167409.4]
  assign regs_402_clock = clock; // @[:@167418.4]
  assign regs_402_reset = io_reset; // @[:@167419.4 RegFile.scala 76:16:@167426.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@167425.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@167429.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@167423.4]
  assign regs_403_clock = clock; // @[:@167432.4]
  assign regs_403_reset = io_reset; // @[:@167433.4 RegFile.scala 76:16:@167440.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@167439.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@167443.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@167437.4]
  assign regs_404_clock = clock; // @[:@167446.4]
  assign regs_404_reset = io_reset; // @[:@167447.4 RegFile.scala 76:16:@167454.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@167453.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@167457.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@167451.4]
  assign regs_405_clock = clock; // @[:@167460.4]
  assign regs_405_reset = io_reset; // @[:@167461.4 RegFile.scala 76:16:@167468.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@167467.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@167471.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@167465.4]
  assign regs_406_clock = clock; // @[:@167474.4]
  assign regs_406_reset = io_reset; // @[:@167475.4 RegFile.scala 76:16:@167482.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@167481.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@167485.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@167479.4]
  assign regs_407_clock = clock; // @[:@167488.4]
  assign regs_407_reset = io_reset; // @[:@167489.4 RegFile.scala 76:16:@167496.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@167495.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@167499.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@167493.4]
  assign regs_408_clock = clock; // @[:@167502.4]
  assign regs_408_reset = io_reset; // @[:@167503.4 RegFile.scala 76:16:@167510.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@167509.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@167513.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@167507.4]
  assign regs_409_clock = clock; // @[:@167516.4]
  assign regs_409_reset = io_reset; // @[:@167517.4 RegFile.scala 76:16:@167524.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@167523.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@167527.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@167521.4]
  assign regs_410_clock = clock; // @[:@167530.4]
  assign regs_410_reset = io_reset; // @[:@167531.4 RegFile.scala 76:16:@167538.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@167537.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@167541.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@167535.4]
  assign regs_411_clock = clock; // @[:@167544.4]
  assign regs_411_reset = io_reset; // @[:@167545.4 RegFile.scala 76:16:@167552.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@167551.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@167555.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@167549.4]
  assign regs_412_clock = clock; // @[:@167558.4]
  assign regs_412_reset = io_reset; // @[:@167559.4 RegFile.scala 76:16:@167566.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@167565.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@167569.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@167563.4]
  assign regs_413_clock = clock; // @[:@167572.4]
  assign regs_413_reset = io_reset; // @[:@167573.4 RegFile.scala 76:16:@167580.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@167579.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@167583.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@167577.4]
  assign regs_414_clock = clock; // @[:@167586.4]
  assign regs_414_reset = io_reset; // @[:@167587.4 RegFile.scala 76:16:@167594.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@167593.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@167597.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@167591.4]
  assign regs_415_clock = clock; // @[:@167600.4]
  assign regs_415_reset = io_reset; // @[:@167601.4 RegFile.scala 76:16:@167608.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@167607.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@167611.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@167605.4]
  assign regs_416_clock = clock; // @[:@167614.4]
  assign regs_416_reset = io_reset; // @[:@167615.4 RegFile.scala 76:16:@167622.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@167621.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@167625.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@167619.4]
  assign regs_417_clock = clock; // @[:@167628.4]
  assign regs_417_reset = io_reset; // @[:@167629.4 RegFile.scala 76:16:@167636.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@167635.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@167639.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@167633.4]
  assign regs_418_clock = clock; // @[:@167642.4]
  assign regs_418_reset = io_reset; // @[:@167643.4 RegFile.scala 76:16:@167650.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@167649.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@167653.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@167647.4]
  assign regs_419_clock = clock; // @[:@167656.4]
  assign regs_419_reset = io_reset; // @[:@167657.4 RegFile.scala 76:16:@167664.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@167663.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@167667.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@167661.4]
  assign regs_420_clock = clock; // @[:@167670.4]
  assign regs_420_reset = io_reset; // @[:@167671.4 RegFile.scala 76:16:@167678.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@167677.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@167681.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@167675.4]
  assign regs_421_clock = clock; // @[:@167684.4]
  assign regs_421_reset = io_reset; // @[:@167685.4 RegFile.scala 76:16:@167692.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@167691.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@167695.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@167689.4]
  assign regs_422_clock = clock; // @[:@167698.4]
  assign regs_422_reset = io_reset; // @[:@167699.4 RegFile.scala 76:16:@167706.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@167705.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@167709.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@167703.4]
  assign regs_423_clock = clock; // @[:@167712.4]
  assign regs_423_reset = io_reset; // @[:@167713.4 RegFile.scala 76:16:@167720.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@167719.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@167723.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@167717.4]
  assign regs_424_clock = clock; // @[:@167726.4]
  assign regs_424_reset = io_reset; // @[:@167727.4 RegFile.scala 76:16:@167734.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@167733.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@167737.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@167731.4]
  assign regs_425_clock = clock; // @[:@167740.4]
  assign regs_425_reset = io_reset; // @[:@167741.4 RegFile.scala 76:16:@167748.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@167747.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@167751.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@167745.4]
  assign regs_426_clock = clock; // @[:@167754.4]
  assign regs_426_reset = io_reset; // @[:@167755.4 RegFile.scala 76:16:@167762.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@167761.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@167765.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@167759.4]
  assign regs_427_clock = clock; // @[:@167768.4]
  assign regs_427_reset = io_reset; // @[:@167769.4 RegFile.scala 76:16:@167776.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@167775.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@167779.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@167773.4]
  assign regs_428_clock = clock; // @[:@167782.4]
  assign regs_428_reset = io_reset; // @[:@167783.4 RegFile.scala 76:16:@167790.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@167789.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@167793.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@167787.4]
  assign regs_429_clock = clock; // @[:@167796.4]
  assign regs_429_reset = io_reset; // @[:@167797.4 RegFile.scala 76:16:@167804.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@167803.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@167807.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@167801.4]
  assign regs_430_clock = clock; // @[:@167810.4]
  assign regs_430_reset = io_reset; // @[:@167811.4 RegFile.scala 76:16:@167818.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@167817.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@167821.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@167815.4]
  assign regs_431_clock = clock; // @[:@167824.4]
  assign regs_431_reset = io_reset; // @[:@167825.4 RegFile.scala 76:16:@167832.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@167831.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@167835.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@167829.4]
  assign regs_432_clock = clock; // @[:@167838.4]
  assign regs_432_reset = io_reset; // @[:@167839.4 RegFile.scala 76:16:@167846.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@167845.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@167849.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@167843.4]
  assign regs_433_clock = clock; // @[:@167852.4]
  assign regs_433_reset = io_reset; // @[:@167853.4 RegFile.scala 76:16:@167860.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@167859.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@167863.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@167857.4]
  assign regs_434_clock = clock; // @[:@167866.4]
  assign regs_434_reset = io_reset; // @[:@167867.4 RegFile.scala 76:16:@167874.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@167873.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@167877.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@167871.4]
  assign regs_435_clock = clock; // @[:@167880.4]
  assign regs_435_reset = io_reset; // @[:@167881.4 RegFile.scala 76:16:@167888.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@167887.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@167891.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@167885.4]
  assign regs_436_clock = clock; // @[:@167894.4]
  assign regs_436_reset = io_reset; // @[:@167895.4 RegFile.scala 76:16:@167902.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@167901.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@167905.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@167899.4]
  assign regs_437_clock = clock; // @[:@167908.4]
  assign regs_437_reset = io_reset; // @[:@167909.4 RegFile.scala 76:16:@167916.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@167915.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@167919.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@167913.4]
  assign regs_438_clock = clock; // @[:@167922.4]
  assign regs_438_reset = io_reset; // @[:@167923.4 RegFile.scala 76:16:@167930.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@167929.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@167933.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@167927.4]
  assign regs_439_clock = clock; // @[:@167936.4]
  assign regs_439_reset = io_reset; // @[:@167937.4 RegFile.scala 76:16:@167944.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@167943.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@167947.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@167941.4]
  assign regs_440_clock = clock; // @[:@167950.4]
  assign regs_440_reset = io_reset; // @[:@167951.4 RegFile.scala 76:16:@167958.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@167957.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@167961.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@167955.4]
  assign regs_441_clock = clock; // @[:@167964.4]
  assign regs_441_reset = io_reset; // @[:@167965.4 RegFile.scala 76:16:@167972.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@167971.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@167975.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@167969.4]
  assign regs_442_clock = clock; // @[:@167978.4]
  assign regs_442_reset = io_reset; // @[:@167979.4 RegFile.scala 76:16:@167986.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@167985.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@167989.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@167983.4]
  assign regs_443_clock = clock; // @[:@167992.4]
  assign regs_443_reset = io_reset; // @[:@167993.4 RegFile.scala 76:16:@168000.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@167999.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@168003.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@167997.4]
  assign regs_444_clock = clock; // @[:@168006.4]
  assign regs_444_reset = io_reset; // @[:@168007.4 RegFile.scala 76:16:@168014.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@168013.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@168017.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@168011.4]
  assign regs_445_clock = clock; // @[:@168020.4]
  assign regs_445_reset = io_reset; // @[:@168021.4 RegFile.scala 76:16:@168028.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@168027.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@168031.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@168025.4]
  assign regs_446_clock = clock; // @[:@168034.4]
  assign regs_446_reset = io_reset; // @[:@168035.4 RegFile.scala 76:16:@168042.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@168041.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@168045.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@168039.4]
  assign regs_447_clock = clock; // @[:@168048.4]
  assign regs_447_reset = io_reset; // @[:@168049.4 RegFile.scala 76:16:@168056.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@168055.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@168059.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@168053.4]
  assign regs_448_clock = clock; // @[:@168062.4]
  assign regs_448_reset = io_reset; // @[:@168063.4 RegFile.scala 76:16:@168070.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@168069.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@168073.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@168067.4]
  assign regs_449_clock = clock; // @[:@168076.4]
  assign regs_449_reset = io_reset; // @[:@168077.4 RegFile.scala 76:16:@168084.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@168083.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@168087.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@168081.4]
  assign regs_450_clock = clock; // @[:@168090.4]
  assign regs_450_reset = io_reset; // @[:@168091.4 RegFile.scala 76:16:@168098.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@168097.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@168101.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@168095.4]
  assign regs_451_clock = clock; // @[:@168104.4]
  assign regs_451_reset = io_reset; // @[:@168105.4 RegFile.scala 76:16:@168112.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@168111.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@168115.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@168109.4]
  assign regs_452_clock = clock; // @[:@168118.4]
  assign regs_452_reset = io_reset; // @[:@168119.4 RegFile.scala 76:16:@168126.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@168125.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@168129.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@168123.4]
  assign regs_453_clock = clock; // @[:@168132.4]
  assign regs_453_reset = io_reset; // @[:@168133.4 RegFile.scala 76:16:@168140.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@168139.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@168143.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@168137.4]
  assign regs_454_clock = clock; // @[:@168146.4]
  assign regs_454_reset = io_reset; // @[:@168147.4 RegFile.scala 76:16:@168154.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@168153.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@168157.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@168151.4]
  assign regs_455_clock = clock; // @[:@168160.4]
  assign regs_455_reset = io_reset; // @[:@168161.4 RegFile.scala 76:16:@168168.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@168167.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@168171.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@168165.4]
  assign regs_456_clock = clock; // @[:@168174.4]
  assign regs_456_reset = io_reset; // @[:@168175.4 RegFile.scala 76:16:@168182.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@168181.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@168185.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@168179.4]
  assign regs_457_clock = clock; // @[:@168188.4]
  assign regs_457_reset = io_reset; // @[:@168189.4 RegFile.scala 76:16:@168196.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@168195.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@168199.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@168193.4]
  assign regs_458_clock = clock; // @[:@168202.4]
  assign regs_458_reset = io_reset; // @[:@168203.4 RegFile.scala 76:16:@168210.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@168209.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@168213.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@168207.4]
  assign regs_459_clock = clock; // @[:@168216.4]
  assign regs_459_reset = io_reset; // @[:@168217.4 RegFile.scala 76:16:@168224.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@168223.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@168227.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@168221.4]
  assign regs_460_clock = clock; // @[:@168230.4]
  assign regs_460_reset = io_reset; // @[:@168231.4 RegFile.scala 76:16:@168238.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@168237.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@168241.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@168235.4]
  assign regs_461_clock = clock; // @[:@168244.4]
  assign regs_461_reset = io_reset; // @[:@168245.4 RegFile.scala 76:16:@168252.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@168251.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@168255.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@168249.4]
  assign regs_462_clock = clock; // @[:@168258.4]
  assign regs_462_reset = io_reset; // @[:@168259.4 RegFile.scala 76:16:@168266.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@168265.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@168269.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@168263.4]
  assign regs_463_clock = clock; // @[:@168272.4]
  assign regs_463_reset = io_reset; // @[:@168273.4 RegFile.scala 76:16:@168280.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@168279.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@168283.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@168277.4]
  assign regs_464_clock = clock; // @[:@168286.4]
  assign regs_464_reset = io_reset; // @[:@168287.4 RegFile.scala 76:16:@168294.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@168293.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@168297.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@168291.4]
  assign regs_465_clock = clock; // @[:@168300.4]
  assign regs_465_reset = io_reset; // @[:@168301.4 RegFile.scala 76:16:@168308.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@168307.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@168311.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@168305.4]
  assign regs_466_clock = clock; // @[:@168314.4]
  assign regs_466_reset = io_reset; // @[:@168315.4 RegFile.scala 76:16:@168322.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@168321.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@168325.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@168319.4]
  assign regs_467_clock = clock; // @[:@168328.4]
  assign regs_467_reset = io_reset; // @[:@168329.4 RegFile.scala 76:16:@168336.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@168335.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@168339.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@168333.4]
  assign regs_468_clock = clock; // @[:@168342.4]
  assign regs_468_reset = io_reset; // @[:@168343.4 RegFile.scala 76:16:@168350.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@168349.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@168353.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@168347.4]
  assign regs_469_clock = clock; // @[:@168356.4]
  assign regs_469_reset = io_reset; // @[:@168357.4 RegFile.scala 76:16:@168364.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@168363.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@168367.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@168361.4]
  assign regs_470_clock = clock; // @[:@168370.4]
  assign regs_470_reset = io_reset; // @[:@168371.4 RegFile.scala 76:16:@168378.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@168377.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@168381.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@168375.4]
  assign regs_471_clock = clock; // @[:@168384.4]
  assign regs_471_reset = io_reset; // @[:@168385.4 RegFile.scala 76:16:@168392.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@168391.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@168395.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@168389.4]
  assign regs_472_clock = clock; // @[:@168398.4]
  assign regs_472_reset = io_reset; // @[:@168399.4 RegFile.scala 76:16:@168406.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@168405.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@168409.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@168403.4]
  assign regs_473_clock = clock; // @[:@168412.4]
  assign regs_473_reset = io_reset; // @[:@168413.4 RegFile.scala 76:16:@168420.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@168419.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@168423.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@168417.4]
  assign regs_474_clock = clock; // @[:@168426.4]
  assign regs_474_reset = io_reset; // @[:@168427.4 RegFile.scala 76:16:@168434.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@168433.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@168437.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@168431.4]
  assign regs_475_clock = clock; // @[:@168440.4]
  assign regs_475_reset = io_reset; // @[:@168441.4 RegFile.scala 76:16:@168448.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@168447.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@168451.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@168445.4]
  assign regs_476_clock = clock; // @[:@168454.4]
  assign regs_476_reset = io_reset; // @[:@168455.4 RegFile.scala 76:16:@168462.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@168461.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@168465.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@168459.4]
  assign regs_477_clock = clock; // @[:@168468.4]
  assign regs_477_reset = io_reset; // @[:@168469.4 RegFile.scala 76:16:@168476.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@168475.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@168479.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@168473.4]
  assign regs_478_clock = clock; // @[:@168482.4]
  assign regs_478_reset = io_reset; // @[:@168483.4 RegFile.scala 76:16:@168490.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@168489.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@168493.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@168487.4]
  assign regs_479_clock = clock; // @[:@168496.4]
  assign regs_479_reset = io_reset; // @[:@168497.4 RegFile.scala 76:16:@168504.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@168503.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@168507.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@168501.4]
  assign regs_480_clock = clock; // @[:@168510.4]
  assign regs_480_reset = io_reset; // @[:@168511.4 RegFile.scala 76:16:@168518.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@168517.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@168521.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@168515.4]
  assign regs_481_clock = clock; // @[:@168524.4]
  assign regs_481_reset = io_reset; // @[:@168525.4 RegFile.scala 76:16:@168532.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@168531.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@168535.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@168529.4]
  assign regs_482_clock = clock; // @[:@168538.4]
  assign regs_482_reset = io_reset; // @[:@168539.4 RegFile.scala 76:16:@168546.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@168545.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@168549.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@168543.4]
  assign regs_483_clock = clock; // @[:@168552.4]
  assign regs_483_reset = io_reset; // @[:@168553.4 RegFile.scala 76:16:@168560.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@168559.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@168563.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@168557.4]
  assign regs_484_clock = clock; // @[:@168566.4]
  assign regs_484_reset = io_reset; // @[:@168567.4 RegFile.scala 76:16:@168574.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@168573.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@168577.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@168571.4]
  assign regs_485_clock = clock; // @[:@168580.4]
  assign regs_485_reset = io_reset; // @[:@168581.4 RegFile.scala 76:16:@168588.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@168587.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@168591.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@168585.4]
  assign regs_486_clock = clock; // @[:@168594.4]
  assign regs_486_reset = io_reset; // @[:@168595.4 RegFile.scala 76:16:@168602.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@168601.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@168605.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@168599.4]
  assign regs_487_clock = clock; // @[:@168608.4]
  assign regs_487_reset = io_reset; // @[:@168609.4 RegFile.scala 76:16:@168616.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@168615.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@168619.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@168613.4]
  assign regs_488_clock = clock; // @[:@168622.4]
  assign regs_488_reset = io_reset; // @[:@168623.4 RegFile.scala 76:16:@168630.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@168629.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@168633.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@168627.4]
  assign regs_489_clock = clock; // @[:@168636.4]
  assign regs_489_reset = io_reset; // @[:@168637.4 RegFile.scala 76:16:@168644.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@168643.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@168647.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@168641.4]
  assign regs_490_clock = clock; // @[:@168650.4]
  assign regs_490_reset = io_reset; // @[:@168651.4 RegFile.scala 76:16:@168658.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@168657.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@168661.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@168655.4]
  assign regs_491_clock = clock; // @[:@168664.4]
  assign regs_491_reset = io_reset; // @[:@168665.4 RegFile.scala 76:16:@168672.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@168671.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@168675.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@168669.4]
  assign regs_492_clock = clock; // @[:@168678.4]
  assign regs_492_reset = io_reset; // @[:@168679.4 RegFile.scala 76:16:@168686.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@168685.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@168689.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@168683.4]
  assign regs_493_clock = clock; // @[:@168692.4]
  assign regs_493_reset = io_reset; // @[:@168693.4 RegFile.scala 76:16:@168700.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@168699.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@168703.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@168697.4]
  assign regs_494_clock = clock; // @[:@168706.4]
  assign regs_494_reset = io_reset; // @[:@168707.4 RegFile.scala 76:16:@168714.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@168713.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@168717.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@168711.4]
  assign regs_495_clock = clock; // @[:@168720.4]
  assign regs_495_reset = io_reset; // @[:@168721.4 RegFile.scala 76:16:@168728.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@168727.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@168731.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@168725.4]
  assign regs_496_clock = clock; // @[:@168734.4]
  assign regs_496_reset = io_reset; // @[:@168735.4 RegFile.scala 76:16:@168742.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@168741.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@168745.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@168739.4]
  assign regs_497_clock = clock; // @[:@168748.4]
  assign regs_497_reset = io_reset; // @[:@168749.4 RegFile.scala 76:16:@168756.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@168755.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@168759.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@168753.4]
  assign regs_498_clock = clock; // @[:@168762.4]
  assign regs_498_reset = io_reset; // @[:@168763.4 RegFile.scala 76:16:@168770.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@168769.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@168773.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@168767.4]
  assign regs_499_clock = clock; // @[:@168776.4]
  assign regs_499_reset = io_reset; // @[:@168777.4 RegFile.scala 76:16:@168784.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@168783.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@168787.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@168781.4]
  assign regs_500_clock = clock; // @[:@168790.4]
  assign regs_500_reset = io_reset; // @[:@168791.4 RegFile.scala 76:16:@168798.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@168797.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@168801.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@168795.4]
  assign regs_501_clock = clock; // @[:@168804.4]
  assign regs_501_reset = io_reset; // @[:@168805.4 RegFile.scala 76:16:@168812.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@168811.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@168815.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@168809.4]
  assign regs_502_clock = clock; // @[:@168818.4]
  assign regs_502_reset = io_reset; // @[:@168819.4 RegFile.scala 76:16:@168826.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@168825.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@168829.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@168823.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@169338.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@169339.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@169340.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@169341.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@169342.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@169343.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@169344.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@169345.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@169346.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@169347.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@169348.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@169349.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@169350.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@169351.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@169352.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@169353.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@169354.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@169355.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@169356.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@169357.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@169358.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@169359.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@169360.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@169361.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@169362.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@169363.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@169364.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@169365.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@169366.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@169367.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@169368.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@169369.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@169370.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@169371.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@169372.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@169373.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@169374.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@169375.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@169376.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@169377.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@169378.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@169379.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@169380.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@169381.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@169382.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@169383.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@169384.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@169385.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@169386.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@169387.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@169388.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@169389.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@169390.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@169391.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@169392.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@169393.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@169394.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@169395.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@169396.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@169397.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@169398.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@169399.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@169400.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@169401.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@169402.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@169403.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@169404.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@169405.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@169406.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@169407.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@169408.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@169409.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@169410.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@169411.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@169412.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@169413.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@169414.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@169415.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@169416.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@169417.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@169418.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@169419.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@169420.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@169421.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@169422.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@169423.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@169424.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@169425.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@169426.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@169427.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@169428.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@169429.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@169430.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@169431.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@169432.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@169433.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@169434.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@169435.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@169436.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@169437.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@169438.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@169439.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@169440.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@169441.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@169442.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@169443.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@169444.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@169445.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@169446.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@169447.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@169448.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@169449.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@169450.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@169451.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@169452.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@169453.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@169454.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@169455.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@169456.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@169457.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@169458.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@169459.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@169460.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@169461.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@169462.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@169463.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@169464.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@169465.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@169466.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@169467.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@169468.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@169469.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@169470.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@169471.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@169472.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@169473.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@169474.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@169475.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@169476.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@169477.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@169478.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@169479.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@169480.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@169481.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@169482.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@169483.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@169484.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@169485.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@169486.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@169487.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@169488.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@169489.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@169490.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@169491.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@169492.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@169493.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@169494.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@169495.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@169496.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@169497.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@169498.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@169499.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@169500.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@169501.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@169502.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@169503.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@169504.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@169505.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@169506.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@169507.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@169508.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@169509.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@169510.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@169511.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@169512.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@169513.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@169514.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@169515.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@169516.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@169517.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@169518.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@169519.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@169520.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@169521.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@169522.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@169523.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@169524.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@169525.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@169526.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@169527.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@169528.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@169529.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@169530.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@169531.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@169532.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@169533.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@169534.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@169535.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@169536.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@169537.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@169538.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@169539.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@169540.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@169541.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@169542.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@169543.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@169544.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@169545.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@169546.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@169547.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@169548.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@169549.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@169550.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@169551.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@169552.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@169553.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@169554.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@169555.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@169556.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@169557.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@169558.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@169559.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@169560.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@169561.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@169562.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@169563.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@169564.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@169565.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@169566.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@169567.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@169568.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@169569.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@169570.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@169571.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@169572.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@169573.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@169574.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@169575.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@169576.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@169577.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@169578.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@169579.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@169580.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@169581.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@169582.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@169583.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@169584.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@169585.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@169586.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@169587.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@169588.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@169589.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@169590.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@169591.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@169592.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@169593.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@169594.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@169595.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@169596.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@169597.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@169598.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@169599.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@169600.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@169601.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@169602.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@169603.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@169604.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@169605.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@169606.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@169607.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@169608.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@169609.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@169610.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@169611.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@169612.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@169613.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@169614.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@169615.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@169616.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@169617.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@169618.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@169619.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@169620.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@169621.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@169622.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@169623.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@169624.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@169625.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@169626.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@169627.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@169628.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@169629.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@169630.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@169631.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@169632.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@169633.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@169634.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@169635.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@169636.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@169637.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@169638.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@169639.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@169640.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@169641.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@169642.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@169643.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@169644.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@169645.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@169646.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@169647.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@169648.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@169649.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@169650.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@169651.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@169652.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@169653.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@169654.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@169655.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@169656.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@169657.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@169658.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@169659.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@169660.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@169661.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@169662.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@169663.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@169664.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@169665.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@169666.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@169667.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@169668.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@169669.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@169670.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@169671.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@169672.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@169673.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@169674.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@169675.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@169676.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@169677.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@169678.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@169679.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@169680.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@169681.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@169682.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@169683.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@169684.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@169685.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@169686.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@169687.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@169688.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@169689.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@169690.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@169691.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@169692.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@169693.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@169694.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@169695.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@169696.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@169697.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@169698.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@169699.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@169700.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@169701.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@169702.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@169703.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@169704.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@169705.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@169706.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@169707.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@169708.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@169709.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@169710.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@169711.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@169712.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@169713.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@169714.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@169715.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@169716.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@169717.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@169718.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@169719.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@169720.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@169721.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@169722.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@169723.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@169724.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@169725.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@169726.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@169727.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@169728.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@169729.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@169730.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@169731.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@169732.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@169733.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@169734.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@169735.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@169736.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@169737.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@169738.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@169739.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@169740.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@169741.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@169742.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@169743.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@169744.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@169745.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@169746.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@169747.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@169748.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@169749.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@169750.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@169751.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@169752.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@169753.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@169754.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@169755.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@169756.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@169757.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@169758.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@169759.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@169760.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@169761.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@169762.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@169763.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@169764.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@169765.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@169766.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@169767.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@169768.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@169769.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@169770.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@169771.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@169772.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@169773.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@169774.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@169775.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@169776.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@169777.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@169778.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@169779.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@169780.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@169781.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@169782.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@169783.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@169784.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@169785.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@169786.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@169787.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@169788.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@169789.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@169790.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@169791.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@169792.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@169793.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@169794.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@169795.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@169796.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@169797.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@169798.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@169799.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@169800.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@169801.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@169802.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@169803.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@169804.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@169805.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@169806.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@169807.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@169808.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@169809.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@169810.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@169811.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@169812.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@169813.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@169814.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@169815.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@169816.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@169817.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@169818.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@169819.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@169820.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@169821.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@169822.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@169823.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@169824.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@169825.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@169826.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@169827.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@169828.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@169829.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@169830.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@169831.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@169832.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@169833.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@169834.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@169835.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@169836.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@169837.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@169838.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@169839.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@169840.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@169841.4]
endmodule
module RetimeWrapper_1222( // @[:@169865.2]
  input         clock, // @[:@169866.4]
  input         reset, // @[:@169867.4]
  input  [39:0] io_in, // @[:@169868.4]
  output [39:0] io_out // @[:@169868.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@169870.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@169870.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@169870.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@169870.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@169870.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@169870.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@169870.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@169883.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@169882.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@169881.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@169880.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@169879.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@169877.4]
endmodule
module FringeFF_503( // @[:@169885.2]
  input         clock, // @[:@169886.4]
  input         reset, // @[:@169887.4]
  input  [39:0] io_in, // @[:@169888.4]
  output [39:0] io_out, // @[:@169888.4]
  input         io_enable // @[:@169888.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@169891.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@169891.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@169891.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@169891.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@169896.4 package.scala 96:25:@169897.4]
  RetimeWrapper_1222 RetimeWrapper ( // @[package.scala 93:22:@169891.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@169896.4 package.scala 96:25:@169897.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@169908.4]
  assign RetimeWrapper_clock = clock; // @[:@169892.4]
  assign RetimeWrapper_reset = reset; // @[:@169893.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@169894.4]
endmodule
module FringeCounter( // @[:@169910.2]
  input   clock, // @[:@169911.4]
  input   reset, // @[:@169912.4]
  input   io_enable, // @[:@169913.4]
  output  io_done // @[:@169913.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@169915.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@169915.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@169915.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@169915.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@169915.4]
  wire [40:0] count; // @[Cat.scala 30:58:@169922.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@169923.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@169924.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@169925.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@169927.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@169915.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@169922.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@169923.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@169924.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@169925.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@169927.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@169938.4]
  assign reg$_clock = clock; // @[:@169916.4]
  assign reg$_reset = reset; // @[:@169917.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@169929.6 FringeCounter.scala 37:15:@169932.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@169920.4]
endmodule
module FringeFF_504( // @[:@169972.2]
  input   clock, // @[:@169973.4]
  input   reset, // @[:@169974.4]
  input   io_in, // @[:@169975.4]
  input   io_reset, // @[:@169975.4]
  output  io_out, // @[:@169975.4]
  input   io_enable // @[:@169975.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@169978.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@169978.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@169978.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@169978.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@169978.4]
  wire  _T_18; // @[package.scala 96:25:@169983.4 package.scala 96:25:@169984.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@169989.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@169978.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@169983.4 package.scala 96:25:@169984.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@169989.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@169995.4]
  assign RetimeWrapper_clock = clock; // @[:@169979.4]
  assign RetimeWrapper_reset = reset; // @[:@169980.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@169982.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@169981.4]
endmodule
module Depulser( // @[:@169997.2]
  input   clock, // @[:@169998.4]
  input   reset, // @[:@169999.4]
  input   io_in, // @[:@170000.4]
  input   io_rst, // @[:@170000.4]
  output  io_out // @[:@170000.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@170002.4]
  wire  r_reset; // @[Depulser.scala 14:17:@170002.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@170002.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@170002.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@170002.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@170002.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@170002.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@170011.4]
  assign r_clock = clock; // @[:@170003.4]
  assign r_reset = reset; // @[:@170004.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@170006.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@170010.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@170009.4]
endmodule
module Fringe( // @[:@170013.2]
  input         clock, // @[:@170014.4]
  input         reset, // @[:@170015.4]
  input  [31:0] io_raddr, // @[:@170016.4]
  input         io_wen, // @[:@170016.4]
  input  [31:0] io_waddr, // @[:@170016.4]
  input  [63:0] io_wdata, // @[:@170016.4]
  output [63:0] io_rdata, // @[:@170016.4]
  output        io_enable, // @[:@170016.4]
  input         io_done, // @[:@170016.4]
  output        io_reset, // @[:@170016.4]
  output [63:0] io_argIns_0, // @[:@170016.4]
  output [63:0] io_argIns_1, // @[:@170016.4]
  input         io_argOuts_0_valid, // @[:@170016.4]
  input  [63:0] io_argOuts_0_bits, // @[:@170016.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@170016.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@170016.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@170016.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@170016.4]
  output        io_memStreams_stores_0_data_ready, // @[:@170016.4]
  input         io_memStreams_stores_0_data_valid, // @[:@170016.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@170016.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@170016.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@170016.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@170016.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@170016.4]
  input         io_dram_0_cmd_ready, // @[:@170016.4]
  output        io_dram_0_cmd_valid, // @[:@170016.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@170016.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@170016.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@170016.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@170016.4]
  input         io_dram_0_wdata_ready, // @[:@170016.4]
  output        io_dram_0_wdata_valid, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@170016.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@170016.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@170016.4]
  output        io_dram_0_rresp_ready, // @[:@170016.4]
  output        io_dram_0_wresp_ready, // @[:@170016.4]
  input         io_dram_0_wresp_valid, // @[:@170016.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@170016.4]
  input         io_dram_1_cmd_ready, // @[:@170016.4]
  output        io_dram_1_cmd_valid, // @[:@170016.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@170016.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@170016.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@170016.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@170016.4]
  input         io_dram_1_wdata_ready, // @[:@170016.4]
  output        io_dram_1_wdata_valid, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@170016.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@170016.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@170016.4]
  output        io_dram_1_rresp_ready, // @[:@170016.4]
  output        io_dram_1_wresp_ready, // @[:@170016.4]
  input         io_dram_1_wresp_valid, // @[:@170016.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@170016.4]
  input         io_dram_2_cmd_ready, // @[:@170016.4]
  output        io_dram_2_cmd_valid, // @[:@170016.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@170016.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@170016.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@170016.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@170016.4]
  input         io_dram_2_wdata_ready, // @[:@170016.4]
  output        io_dram_2_wdata_valid, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@170016.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@170016.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@170016.4]
  output        io_dram_2_rresp_ready, // @[:@170016.4]
  output        io_dram_2_wresp_ready, // @[:@170016.4]
  input         io_dram_2_wresp_valid, // @[:@170016.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@170016.4]
  input         io_dram_3_cmd_ready, // @[:@170016.4]
  output        io_dram_3_cmd_valid, // @[:@170016.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@170016.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@170016.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@170016.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@170016.4]
  input         io_dram_3_wdata_ready, // @[:@170016.4]
  output        io_dram_3_wdata_valid, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@170016.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@170016.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@170016.4]
  output        io_dram_3_rresp_ready, // @[:@170016.4]
  output        io_dram_3_wresp_ready, // @[:@170016.4]
  input         io_dram_3_wresp_valid, // @[:@170016.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@170016.4]
  input         io_heap_0_req_valid, // @[:@170016.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@170016.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@170016.4]
  output        io_heap_0_resp_valid, // @[:@170016.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@170016.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@170016.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@170022.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@170022.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@170022.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@170022.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@171015.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@171015.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@171015.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@171975.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@171975.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@171975.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@172935.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@172935.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@172935.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@172935.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@173895.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@173895.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@173895.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@173895.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@173895.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@173895.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@173895.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@173895.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@173895.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@173895.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@173895.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@173895.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@173904.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@173904.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@173904.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@173904.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@173904.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@173904.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@173904.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@173904.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@173904.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@173904.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@173904.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@173904.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@173904.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@173904.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@173904.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@173904.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@175954.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@175954.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@175954.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@175954.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@175973.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@175973.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@175973.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@175973.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@175973.4]
  wire [63:0] _T_1020; // @[:@175931.4 :@175932.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@175933.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@175935.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@175937.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@175939.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@175941.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@175943.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@175945.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@175981.4]
  reg  _T_1047; // @[package.scala 152:20:@175984.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@175986.4]
  wire  _T_1049; // @[package.scala 153:8:@175987.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@175991.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@175992.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@175995.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@175996.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@175998.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@175999.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@176001.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@176004.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@175983.4 Fringe.scala 163:24:@176002.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@175983.4 Fringe.scala 162:28:@176000.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@176005.4]
  wire  alloc; // @[Fringe.scala 202:38:@177635.4]
  wire  dealloc; // @[Fringe.scala 203:40:@177636.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@177637.4]
  reg  _T_1572; // @[package.scala 152:20:@177638.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@177640.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@170022.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@171015.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@171975.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@172935.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@173895.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@173904.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@175954.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@175973.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@175931.4 :@175932.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@175933.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@175935.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@175937.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@175939.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@175941.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@175943.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@175945.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@175981.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@175986.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@175987.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@175991.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@175992.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@175995.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@175996.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@175998.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@175999.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@176001.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@176004.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@175983.4 Fringe.scala 163:24:@176002.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@175983.4 Fringe.scala 162:28:@176000.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@176005.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@177635.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@177636.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@177637.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@177640.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@175929.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@175949.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@175950.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@175971.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@175972.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@170941.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@170937.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@170932.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@170931.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@177133.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@177132.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@177131.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@177129.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@177128.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@177126.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@177110.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@177111.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@177112.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@177113.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@177114.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@177115.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@177116.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@177117.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@177118.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@177119.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@177120.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@177121.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@177122.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@177123.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@177124.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@177125.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@177046.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@177047.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@177048.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@177049.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@177050.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@177051.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@177052.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@177053.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@177054.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@177055.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@177056.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@177057.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@177058.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@177059.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@177060.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@177061.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@177062.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@177063.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@177064.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@177065.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@177066.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@177067.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@177068.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@177069.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@177070.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@177071.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@177072.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@177073.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@177074.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@177075.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@177076.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@177077.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@177078.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@177079.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@177080.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@177081.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@177082.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@177083.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@177084.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@177085.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@177086.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@177087.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@177088.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@177089.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@177090.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@177091.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@177092.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@177093.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@177094.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@177095.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@177096.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@177097.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@177098.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@177099.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@177100.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@177101.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@177102.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@177103.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@177104.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@177105.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@177106.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@177107.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@177108.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@177109.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@177045.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@177044.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@177025.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@177245.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@177244.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@177243.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@177241.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@177240.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@177238.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@177222.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@177223.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@177224.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@177225.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@177226.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@177227.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@177228.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@177229.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@177230.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@177231.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@177232.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@177233.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@177234.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@177235.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@177236.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@177237.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@177158.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@177159.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@177160.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@177161.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@177162.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@177163.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@177164.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@177165.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@177166.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@177167.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@177168.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@177169.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@177170.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@177171.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@177172.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@177173.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@177174.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@177175.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@177176.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@177177.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@177178.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@177179.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@177180.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@177181.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@177182.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@177183.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@177184.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@177185.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@177186.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@177187.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@177188.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@177189.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@177190.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@177191.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@177192.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@177193.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@177194.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@177195.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@177196.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@177197.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@177198.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@177199.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@177200.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@177201.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@177202.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@177203.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@177204.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@177205.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@177206.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@177207.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@177208.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@177209.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@177210.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@177211.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@177212.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@177213.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@177214.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@177215.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@177216.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@177217.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@177218.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@177219.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@177220.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@177221.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@177157.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@177156.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@177137.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@177357.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@177356.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@177355.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@177353.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@177352.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@177350.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@177334.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@177335.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@177336.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@177337.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@177338.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@177339.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@177340.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@177341.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@177342.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@177343.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@177344.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@177345.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@177346.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@177347.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@177348.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@177349.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@177270.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@177271.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@177272.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@177273.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@177274.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@177275.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@177276.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@177277.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@177278.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@177279.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@177280.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@177281.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@177282.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@177283.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@177284.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@177285.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@177286.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@177287.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@177288.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@177289.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@177290.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@177291.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@177292.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@177293.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@177294.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@177295.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@177296.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@177297.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@177298.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@177299.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@177300.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@177301.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@177302.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@177303.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@177304.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@177305.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@177306.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@177307.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@177308.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@177309.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@177310.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@177311.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@177312.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@177313.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@177314.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@177315.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@177316.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@177317.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@177318.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@177319.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@177320.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@177321.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@177322.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@177323.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@177324.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@177325.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@177326.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@177327.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@177328.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@177329.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@177330.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@177331.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@177332.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@177333.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@177269.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@177268.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@177249.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@177469.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@177468.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@177467.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@177465.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@177464.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@177462.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@177446.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@177447.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@177448.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@177449.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@177450.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@177451.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@177452.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@177453.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@177454.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@177455.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@177456.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@177457.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@177458.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@177459.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@177460.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@177461.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@177382.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@177383.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@177384.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@177385.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@177386.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@177387.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@177388.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@177389.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@177390.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@177391.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@177392.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@177393.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@177394.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@177395.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@177396.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@177397.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@177398.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@177399.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@177400.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@177401.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@177402.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@177403.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@177404.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@177405.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@177406.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@177407.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@177408.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@177409.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@177410.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@177411.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@177412.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@177413.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@177414.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@177415.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@177416.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@177417.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@177418.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@177419.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@177420.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@177421.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@177422.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@177423.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@177424.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@177425.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@177426.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@177427.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@177428.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@177429.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@177430.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@177431.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@177432.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@177433.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@177434.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@177435.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@177436.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@177437.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@177438.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@177439.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@177440.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@177441.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@177442.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@177443.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@177444.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@177445.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@177381.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@177380.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@177361.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@173900.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@173899.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@173898.4]
  assign dramArbs_0_clock = clock; // @[:@170023.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@170024.4 Fringe.scala 187:30:@177015.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@177019.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@170940.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@170939.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@170938.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@170936.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@170935.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@170934.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@170933.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@177134.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@177127.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@177024.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@177023.4]
  assign dramArbs_1_clock = clock; // @[:@171016.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@171017.4 Fringe.scala 187:30:@177016.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@177020.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@177246.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@177239.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@177136.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@177135.4]
  assign dramArbs_2_clock = clock; // @[:@171976.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@171977.4 Fringe.scala 187:30:@177017.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@177021.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@177358.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@177351.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@177248.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@177247.4]
  assign dramArbs_3_clock = clock; // @[:@172936.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@172937.4 Fringe.scala 187:30:@177018.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@177022.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@177470.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@177463.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@177360.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@177359.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@173903.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@173902.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@173901.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@177642.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@177643.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@177644.4]
  assign regs_clock = clock; // @[:@173905.4]
  assign regs_reset = reset; // @[:@173906.4 Fringe.scala 139:14:@175953.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@175925.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@175927.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@175926.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@175928.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@175951.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@176003.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@176007.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@176010.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@176009.4]
  assign timeoutCtr_clock = clock; // @[:@175955.4]
  assign timeoutCtr_reset = reset; // @[:@175956.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@175970.4]
  assign depulser_clock = clock; // @[:@175974.4]
  assign depulser_reset = reset; // @[:@175975.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@175980.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@175982.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@177659.2]
  input         clock, // @[:@177660.4]
  input         reset, // @[:@177661.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@177662.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@177662.4]
  input         io_S_AXI_AWVALID, // @[:@177662.4]
  output        io_S_AXI_AWREADY, // @[:@177662.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@177662.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@177662.4]
  input         io_S_AXI_ARVALID, // @[:@177662.4]
  output        io_S_AXI_ARREADY, // @[:@177662.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@177662.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@177662.4]
  input         io_S_AXI_WVALID, // @[:@177662.4]
  output        io_S_AXI_WREADY, // @[:@177662.4]
  output [31:0] io_S_AXI_RDATA, // @[:@177662.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@177662.4]
  output        io_S_AXI_RVALID, // @[:@177662.4]
  input         io_S_AXI_RREADY, // @[:@177662.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@177662.4]
  output        io_S_AXI_BVALID, // @[:@177662.4]
  input         io_S_AXI_BREADY, // @[:@177662.4]
  output [31:0] io_raddr, // @[:@177662.4]
  output        io_wen, // @[:@177662.4]
  output [31:0] io_waddr, // @[:@177662.4]
  output [31:0] io_wdata, // @[:@177662.4]
  input  [31:0] io_rdata // @[:@177662.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@177664.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@177688.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@177684.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@177680.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@177679.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@177678.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@177677.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@177675.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@177674.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@177696.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@177699.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@177697.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@177698.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@177700.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@177695.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@177692.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@177691.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@177690.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@177689.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@177687.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@177686.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@177685.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@177683.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@177682.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@177681.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@177676.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@177673.4]
endmodule
module MAGToAXI4Bridge( // @[:@177702.2]
  output         io_in_cmd_ready, // @[:@177705.4]
  input          io_in_cmd_valid, // @[:@177705.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@177705.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@177705.4]
  input          io_in_cmd_bits_isWr, // @[:@177705.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@177705.4]
  output         io_in_wdata_ready, // @[:@177705.4]
  input          io_in_wdata_valid, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@177705.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@177705.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@177705.4]
  input          io_in_wdata_bits_wlast, // @[:@177705.4]
  input          io_in_rresp_ready, // @[:@177705.4]
  input          io_in_wresp_ready, // @[:@177705.4]
  output         io_in_wresp_valid, // @[:@177705.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@177705.4]
  output [31:0]  io_M_AXI_AWID, // @[:@177705.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@177705.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@177705.4]
  output         io_M_AXI_AWVALID, // @[:@177705.4]
  input          io_M_AXI_AWREADY, // @[:@177705.4]
  output [31:0]  io_M_AXI_ARID, // @[:@177705.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@177705.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@177705.4]
  output         io_M_AXI_ARVALID, // @[:@177705.4]
  input          io_M_AXI_ARREADY, // @[:@177705.4]
  output [511:0] io_M_AXI_WDATA, // @[:@177705.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@177705.4]
  output         io_M_AXI_WLAST, // @[:@177705.4]
  output         io_M_AXI_WVALID, // @[:@177705.4]
  input          io_M_AXI_WREADY, // @[:@177705.4]
  output         io_M_AXI_RREADY, // @[:@177705.4]
  input  [31:0]  io_M_AXI_BID, // @[:@177705.4]
  input          io_M_AXI_BVALID, // @[:@177705.4]
  output         io_M_AXI_BREADY // @[:@177705.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@177862.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@177863.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@177864.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@177872.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@177899.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@177904.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@177915.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@177924.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@177933.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@177942.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@177951.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@177960.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@177968.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@177862.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@177863.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@177864.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@177872.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@177899.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@177904.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@177915.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@177924.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@177933.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@177942.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@177951.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@177960.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@177968.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@177876.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@177973.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@178026.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@178028.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@177877.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@177878.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@177882.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@177890.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@177860.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@177861.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@177865.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@177874.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@177906.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@177970.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@177971.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@177972.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@178023.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@178024.4]
endmodule
module FringeZynq( // @[:@179014.2]
  input          clock, // @[:@179015.4]
  input          reset, // @[:@179016.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@179017.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@179017.4]
  input          io_S_AXI_AWVALID, // @[:@179017.4]
  output         io_S_AXI_AWREADY, // @[:@179017.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@179017.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@179017.4]
  input          io_S_AXI_ARVALID, // @[:@179017.4]
  output         io_S_AXI_ARREADY, // @[:@179017.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@179017.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@179017.4]
  input          io_S_AXI_WVALID, // @[:@179017.4]
  output         io_S_AXI_WREADY, // @[:@179017.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@179017.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@179017.4]
  output         io_S_AXI_RVALID, // @[:@179017.4]
  input          io_S_AXI_RREADY, // @[:@179017.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@179017.4]
  output         io_S_AXI_BVALID, // @[:@179017.4]
  input          io_S_AXI_BREADY, // @[:@179017.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@179017.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@179017.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@179017.4]
  output         io_M_AXI_0_AWVALID, // @[:@179017.4]
  input          io_M_AXI_0_AWREADY, // @[:@179017.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@179017.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@179017.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@179017.4]
  output         io_M_AXI_0_ARVALID, // @[:@179017.4]
  input          io_M_AXI_0_ARREADY, // @[:@179017.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@179017.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@179017.4]
  output         io_M_AXI_0_WLAST, // @[:@179017.4]
  output         io_M_AXI_0_WVALID, // @[:@179017.4]
  input          io_M_AXI_0_WREADY, // @[:@179017.4]
  output         io_M_AXI_0_RREADY, // @[:@179017.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@179017.4]
  input          io_M_AXI_0_BVALID, // @[:@179017.4]
  output         io_M_AXI_0_BREADY, // @[:@179017.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@179017.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@179017.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@179017.4]
  output         io_M_AXI_1_AWVALID, // @[:@179017.4]
  input          io_M_AXI_1_AWREADY, // @[:@179017.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@179017.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@179017.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@179017.4]
  output         io_M_AXI_1_ARVALID, // @[:@179017.4]
  input          io_M_AXI_1_ARREADY, // @[:@179017.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@179017.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@179017.4]
  output         io_M_AXI_1_WLAST, // @[:@179017.4]
  output         io_M_AXI_1_WVALID, // @[:@179017.4]
  input          io_M_AXI_1_WREADY, // @[:@179017.4]
  output         io_M_AXI_1_RREADY, // @[:@179017.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@179017.4]
  input          io_M_AXI_1_BVALID, // @[:@179017.4]
  output         io_M_AXI_1_BREADY, // @[:@179017.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@179017.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@179017.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@179017.4]
  output         io_M_AXI_2_AWVALID, // @[:@179017.4]
  input          io_M_AXI_2_AWREADY, // @[:@179017.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@179017.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@179017.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@179017.4]
  output         io_M_AXI_2_ARVALID, // @[:@179017.4]
  input          io_M_AXI_2_ARREADY, // @[:@179017.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@179017.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@179017.4]
  output         io_M_AXI_2_WLAST, // @[:@179017.4]
  output         io_M_AXI_2_WVALID, // @[:@179017.4]
  input          io_M_AXI_2_WREADY, // @[:@179017.4]
  output         io_M_AXI_2_RREADY, // @[:@179017.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@179017.4]
  input          io_M_AXI_2_BVALID, // @[:@179017.4]
  output         io_M_AXI_2_BREADY, // @[:@179017.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@179017.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@179017.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@179017.4]
  output         io_M_AXI_3_AWVALID, // @[:@179017.4]
  input          io_M_AXI_3_AWREADY, // @[:@179017.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@179017.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@179017.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@179017.4]
  output         io_M_AXI_3_ARVALID, // @[:@179017.4]
  input          io_M_AXI_3_ARREADY, // @[:@179017.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@179017.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@179017.4]
  output         io_M_AXI_3_WLAST, // @[:@179017.4]
  output         io_M_AXI_3_WVALID, // @[:@179017.4]
  input          io_M_AXI_3_WREADY, // @[:@179017.4]
  output         io_M_AXI_3_RREADY, // @[:@179017.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@179017.4]
  input          io_M_AXI_3_BVALID, // @[:@179017.4]
  output         io_M_AXI_3_BREADY, // @[:@179017.4]
  output         io_enable, // @[:@179017.4]
  input          io_done, // @[:@179017.4]
  output         io_reset, // @[:@179017.4]
  output [63:0]  io_argIns_0, // @[:@179017.4]
  output [63:0]  io_argIns_1, // @[:@179017.4]
  input          io_argOuts_0_valid, // @[:@179017.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@179017.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@179017.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@179017.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@179017.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@179017.4]
  output         io_memStreams_stores_0_data_ready, // @[:@179017.4]
  input          io_memStreams_stores_0_data_valid, // @[:@179017.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@179017.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@179017.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@179017.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@179017.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@179017.4]
  input          io_heap_0_req_valid, // @[:@179017.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@179017.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@179017.4]
  output         io_heap_0_resp_valid, // @[:@179017.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@179017.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@179017.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@179488.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@179488.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@179488.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@180394.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@180394.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@180394.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@180394.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@180394.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@180394.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@180394.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@180394.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@180394.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@180394.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@180394.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@180394.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@180394.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@180394.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@180394.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@180544.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@180544.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@180544.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@180544.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@180544.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@180544.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@180544.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@180700.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@180700.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@180700.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@180700.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@180700.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@180700.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@180700.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@180856.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@180856.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@180856.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@180856.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@180856.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@180856.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@180856.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@181012.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@181012.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@181012.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@181012.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@181012.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@181012.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@181012.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@181012.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@179488.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@180394.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@180544.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@180700.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@180856.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@181012.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@180412.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@180408.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@180404.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@180403.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@180402.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@180401.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@180399.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@180398.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@180699.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@180697.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@180696.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@180689.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@180687.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@180685.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@180684.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@180677.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@180675.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@180674.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@180673.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@180672.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@180664.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@180659.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@180855.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@180853.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@180852.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@180845.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@180843.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@180841.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@180840.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@180833.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@180831.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@180830.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@180829.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@180828.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@180820.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@180815.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@181011.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@181009.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@181008.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@181001.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@180999.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@180997.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@180996.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@180989.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@180987.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@180986.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@180985.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@180984.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@180976.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@180971.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@181167.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@181165.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@181164.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@181157.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@181155.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@181153.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@181152.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@181145.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@181143.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@181142.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@181141.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@181140.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@181132.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@181127.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@180422.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@180426.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@180427.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@180428.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@180515.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@180511.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@180506.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@180505.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@180540.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@180539.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@180538.4]
  assign fringeCommon_clock = clock; // @[:@179489.4]
  assign fringeCommon_reset = reset; // @[:@179490.4 FringeZynq.scala 117:22:@180425.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@180416.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@180417.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@180418.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@180419.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@180423.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@180430.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@180429.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@180514.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@180513.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@180512.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@180510.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@180509.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@180508.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@180507.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@180658.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@180651.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@180548.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@180547.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@180814.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@180807.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@180704.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@180703.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@180970.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@180963.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@180860.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@180859.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@181126.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@181119.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@181016.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@181015.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@180543.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@180542.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@180541.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@180395.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@180396.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@180415.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@180414.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@180413.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@180411.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@180410.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@180409.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@180407.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@180406.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@180405.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@180400.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@180397.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@180420.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@180657.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@180656.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@180655.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@180653.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@180652.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@180650.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@180634.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@180635.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@180636.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@180637.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@180638.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@180639.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@180640.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@180641.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@180642.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@180643.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@180644.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@180645.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@180646.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@180647.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@180648.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@180649.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@180570.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@180571.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@180572.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@180573.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@180574.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@180575.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@180576.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@180577.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@180578.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@180579.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@180580.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@180581.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@180582.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@180583.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@180584.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@180585.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@180586.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@180587.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@180588.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@180589.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@180590.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@180591.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@180592.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@180593.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@180594.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@180595.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@180596.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@180597.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@180598.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@180599.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@180600.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@180601.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@180602.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@180603.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@180604.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@180605.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@180606.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@180607.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@180608.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@180609.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@180610.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@180611.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@180612.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@180613.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@180614.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@180615.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@180616.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@180617.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@180618.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@180619.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@180620.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@180621.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@180622.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@180623.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@180624.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@180625.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@180626.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@180627.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@180628.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@180629.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@180630.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@180631.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@180632.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@180633.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@180569.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@180568.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@180549.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@180688.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@180676.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@180671.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@180663.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@180660.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@180813.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@180812.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@180811.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@180809.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@180808.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@180806.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@180790.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@180791.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@180792.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@180793.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@180794.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@180795.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@180796.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@180797.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@180798.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@180799.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@180800.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@180801.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@180802.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@180803.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@180804.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@180805.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@180726.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@180727.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@180728.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@180729.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@180730.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@180731.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@180732.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@180733.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@180734.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@180735.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@180736.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@180737.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@180738.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@180739.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@180740.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@180741.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@180742.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@180743.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@180744.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@180745.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@180746.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@180747.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@180748.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@180749.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@180750.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@180751.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@180752.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@180753.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@180754.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@180755.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@180756.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@180757.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@180758.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@180759.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@180760.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@180761.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@180762.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@180763.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@180764.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@180765.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@180766.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@180767.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@180768.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@180769.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@180770.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@180771.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@180772.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@180773.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@180774.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@180775.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@180776.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@180777.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@180778.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@180779.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@180780.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@180781.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@180782.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@180783.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@180784.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@180785.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@180786.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@180787.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@180788.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@180789.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@180725.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@180724.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@180705.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@180844.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@180832.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@180827.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@180819.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@180816.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@180969.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@180968.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@180967.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@180965.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@180964.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@180962.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@180946.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@180947.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@180948.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@180949.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@180950.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@180951.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@180952.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@180953.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@180954.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@180955.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@180956.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@180957.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@180958.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@180959.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@180960.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@180961.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@180882.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@180883.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@180884.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@180885.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@180886.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@180887.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@180888.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@180889.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@180890.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@180891.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@180892.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@180893.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@180894.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@180895.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@180896.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@180897.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@180898.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@180899.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@180900.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@180901.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@180902.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@180903.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@180904.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@180905.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@180906.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@180907.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@180908.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@180909.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@180910.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@180911.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@180912.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@180913.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@180914.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@180915.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@180916.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@180917.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@180918.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@180919.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@180920.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@180921.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@180922.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@180923.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@180924.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@180925.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@180926.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@180927.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@180928.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@180929.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@180930.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@180931.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@180932.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@180933.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@180934.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@180935.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@180936.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@180937.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@180938.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@180939.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@180940.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@180941.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@180942.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@180943.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@180944.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@180945.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@180881.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@180880.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@180861.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@181000.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@180988.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@180983.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@180975.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@180972.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@181125.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@181124.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@181123.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@181121.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@181120.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@181118.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@181102.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@181103.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@181104.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@181105.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@181106.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@181107.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@181108.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@181109.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@181110.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@181111.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@181112.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@181113.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@181114.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@181115.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@181116.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@181117.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@181038.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@181039.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@181040.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@181041.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@181042.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@181043.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@181044.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@181045.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@181046.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@181047.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@181048.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@181049.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@181050.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@181051.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@181052.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@181053.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@181054.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@181055.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@181056.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@181057.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@181058.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@181059.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@181060.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@181061.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@181062.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@181063.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@181064.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@181065.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@181066.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@181067.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@181068.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@181069.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@181070.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@181071.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@181072.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@181073.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@181074.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@181075.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@181076.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@181077.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@181078.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@181079.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@181080.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@181081.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@181082.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@181083.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@181084.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@181085.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@181086.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@181087.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@181088.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@181089.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@181090.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@181091.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@181092.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@181093.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@181094.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@181095.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@181096.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@181097.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@181098.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@181099.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@181100.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@181101.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@181037.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@181036.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@181017.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@181156.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@181144.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@181139.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@181131.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@181128.4]
endmodule
module SpatialIP( // @[:@181169.2]
  input          clock, // @[:@181170.4]
  input          reset, // @[:@181171.4]
  input          io_raddr, // @[:@181172.4]
  input          io_wen, // @[:@181172.4]
  input          io_waddr, // @[:@181172.4]
  input          io_wdata, // @[:@181172.4]
  output         io_rdata, // @[:@181172.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@181172.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@181172.4]
  input          io_S_AXI_AWVALID, // @[:@181172.4]
  output         io_S_AXI_AWREADY, // @[:@181172.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@181172.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@181172.4]
  input          io_S_AXI_ARVALID, // @[:@181172.4]
  output         io_S_AXI_ARREADY, // @[:@181172.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@181172.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@181172.4]
  input          io_S_AXI_WVALID, // @[:@181172.4]
  output         io_S_AXI_WREADY, // @[:@181172.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@181172.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@181172.4]
  output         io_S_AXI_RVALID, // @[:@181172.4]
  input          io_S_AXI_RREADY, // @[:@181172.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@181172.4]
  output         io_S_AXI_BVALID, // @[:@181172.4]
  input          io_S_AXI_BREADY, // @[:@181172.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@181172.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@181172.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@181172.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@181172.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@181172.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@181172.4]
  output         io_M_AXI_0_AWLOCK, // @[:@181172.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@181172.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@181172.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@181172.4]
  output         io_M_AXI_0_AWVALID, // @[:@181172.4]
  input          io_M_AXI_0_AWREADY, // @[:@181172.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@181172.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@181172.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@181172.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@181172.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@181172.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@181172.4]
  output         io_M_AXI_0_ARLOCK, // @[:@181172.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@181172.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@181172.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@181172.4]
  output         io_M_AXI_0_ARVALID, // @[:@181172.4]
  input          io_M_AXI_0_ARREADY, // @[:@181172.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@181172.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@181172.4]
  output         io_M_AXI_0_WLAST, // @[:@181172.4]
  output         io_M_AXI_0_WVALID, // @[:@181172.4]
  input          io_M_AXI_0_WREADY, // @[:@181172.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@181172.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@181172.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@181172.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@181172.4]
  input          io_M_AXI_0_RLAST, // @[:@181172.4]
  input          io_M_AXI_0_RVALID, // @[:@181172.4]
  output         io_M_AXI_0_RREADY, // @[:@181172.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@181172.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@181172.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@181172.4]
  input          io_M_AXI_0_BVALID, // @[:@181172.4]
  output         io_M_AXI_0_BREADY, // @[:@181172.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@181172.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@181172.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@181172.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@181172.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@181172.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@181172.4]
  output         io_M_AXI_1_AWLOCK, // @[:@181172.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@181172.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@181172.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@181172.4]
  output         io_M_AXI_1_AWVALID, // @[:@181172.4]
  input          io_M_AXI_1_AWREADY, // @[:@181172.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@181172.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@181172.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@181172.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@181172.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@181172.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@181172.4]
  output         io_M_AXI_1_ARLOCK, // @[:@181172.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@181172.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@181172.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@181172.4]
  output         io_M_AXI_1_ARVALID, // @[:@181172.4]
  input          io_M_AXI_1_ARREADY, // @[:@181172.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@181172.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@181172.4]
  output         io_M_AXI_1_WLAST, // @[:@181172.4]
  output         io_M_AXI_1_WVALID, // @[:@181172.4]
  input          io_M_AXI_1_WREADY, // @[:@181172.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@181172.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@181172.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@181172.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@181172.4]
  input          io_M_AXI_1_RLAST, // @[:@181172.4]
  input          io_M_AXI_1_RVALID, // @[:@181172.4]
  output         io_M_AXI_1_RREADY, // @[:@181172.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@181172.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@181172.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@181172.4]
  input          io_M_AXI_1_BVALID, // @[:@181172.4]
  output         io_M_AXI_1_BREADY, // @[:@181172.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@181172.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@181172.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@181172.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@181172.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@181172.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@181172.4]
  output         io_M_AXI_2_AWLOCK, // @[:@181172.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@181172.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@181172.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@181172.4]
  output         io_M_AXI_2_AWVALID, // @[:@181172.4]
  input          io_M_AXI_2_AWREADY, // @[:@181172.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@181172.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@181172.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@181172.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@181172.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@181172.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@181172.4]
  output         io_M_AXI_2_ARLOCK, // @[:@181172.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@181172.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@181172.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@181172.4]
  output         io_M_AXI_2_ARVALID, // @[:@181172.4]
  input          io_M_AXI_2_ARREADY, // @[:@181172.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@181172.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@181172.4]
  output         io_M_AXI_2_WLAST, // @[:@181172.4]
  output         io_M_AXI_2_WVALID, // @[:@181172.4]
  input          io_M_AXI_2_WREADY, // @[:@181172.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@181172.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@181172.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@181172.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@181172.4]
  input          io_M_AXI_2_RLAST, // @[:@181172.4]
  input          io_M_AXI_2_RVALID, // @[:@181172.4]
  output         io_M_AXI_2_RREADY, // @[:@181172.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@181172.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@181172.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@181172.4]
  input          io_M_AXI_2_BVALID, // @[:@181172.4]
  output         io_M_AXI_2_BREADY, // @[:@181172.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@181172.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@181172.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@181172.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@181172.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@181172.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@181172.4]
  output         io_M_AXI_3_AWLOCK, // @[:@181172.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@181172.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@181172.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@181172.4]
  output         io_M_AXI_3_AWVALID, // @[:@181172.4]
  input          io_M_AXI_3_AWREADY, // @[:@181172.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@181172.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@181172.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@181172.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@181172.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@181172.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@181172.4]
  output         io_M_AXI_3_ARLOCK, // @[:@181172.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@181172.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@181172.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@181172.4]
  output         io_M_AXI_3_ARVALID, // @[:@181172.4]
  input          io_M_AXI_3_ARREADY, // @[:@181172.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@181172.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@181172.4]
  output         io_M_AXI_3_WLAST, // @[:@181172.4]
  output         io_M_AXI_3_WVALID, // @[:@181172.4]
  input          io_M_AXI_3_WREADY, // @[:@181172.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@181172.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@181172.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@181172.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@181172.4]
  input          io_M_AXI_3_RLAST, // @[:@181172.4]
  input          io_M_AXI_3_RVALID, // @[:@181172.4]
  output         io_M_AXI_3_RREADY, // @[:@181172.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@181172.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@181172.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@181172.4]
  input          io_M_AXI_3_BVALID, // @[:@181172.4]
  output         io_M_AXI_3_BREADY, // @[:@181172.4]
  input          io_TOP_AXI_AWID, // @[:@181172.4]
  input          io_TOP_AXI_AWUSER, // @[:@181172.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@181172.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@181172.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@181172.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@181172.4]
  input          io_TOP_AXI_AWLOCK, // @[:@181172.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@181172.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@181172.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@181172.4]
  input          io_TOP_AXI_AWVALID, // @[:@181172.4]
  input          io_TOP_AXI_AWREADY, // @[:@181172.4]
  input          io_TOP_AXI_ARID, // @[:@181172.4]
  input          io_TOP_AXI_ARUSER, // @[:@181172.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@181172.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@181172.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@181172.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@181172.4]
  input          io_TOP_AXI_ARLOCK, // @[:@181172.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@181172.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@181172.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@181172.4]
  input          io_TOP_AXI_ARVALID, // @[:@181172.4]
  input          io_TOP_AXI_ARREADY, // @[:@181172.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@181172.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@181172.4]
  input          io_TOP_AXI_WLAST, // @[:@181172.4]
  input          io_TOP_AXI_WVALID, // @[:@181172.4]
  input          io_TOP_AXI_WREADY, // @[:@181172.4]
  input          io_TOP_AXI_RID, // @[:@181172.4]
  input          io_TOP_AXI_RUSER, // @[:@181172.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@181172.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@181172.4]
  input          io_TOP_AXI_RLAST, // @[:@181172.4]
  input          io_TOP_AXI_RVALID, // @[:@181172.4]
  input          io_TOP_AXI_RREADY, // @[:@181172.4]
  input          io_TOP_AXI_BID, // @[:@181172.4]
  input          io_TOP_AXI_BUSER, // @[:@181172.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@181172.4]
  input          io_TOP_AXI_BVALID, // @[:@181172.4]
  input          io_TOP_AXI_BREADY, // @[:@181172.4]
  input          io_DWIDTH_AXI_AWID, // @[:@181172.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@181172.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@181172.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@181172.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@181172.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@181172.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@181172.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@181172.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@181172.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@181172.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@181172.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@181172.4]
  input          io_DWIDTH_AXI_ARID, // @[:@181172.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@181172.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@181172.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@181172.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@181172.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@181172.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@181172.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@181172.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@181172.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@181172.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@181172.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@181172.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@181172.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@181172.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@181172.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@181172.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@181172.4]
  input          io_DWIDTH_AXI_RID, // @[:@181172.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@181172.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@181172.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@181172.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@181172.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@181172.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@181172.4]
  input          io_DWIDTH_AXI_BID, // @[:@181172.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@181172.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@181172.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@181172.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@181172.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@181172.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@181172.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@181172.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@181172.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@181172.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@181172.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@181172.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@181172.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@181172.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@181172.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@181172.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@181172.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@181172.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@181172.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@181172.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@181172.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@181172.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@181172.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@181172.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@181172.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@181172.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@181172.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@181172.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@181172.4]
  input          io_PROTOCOL_AXI_RID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@181172.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@181172.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@181172.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@181172.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@181172.4]
  input          io_PROTOCOL_AXI_BID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@181172.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@181172.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@181172.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@181172.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@181172.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@181172.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@181172.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@181172.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@181172.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@181172.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@181172.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@181172.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@181172.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@181172.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@181172.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@181172.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@181172.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@181172.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@181172.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@181172.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@181172.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@181172.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@181172.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@181172.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@181174.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@181174.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@181174.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@181174.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@181174.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@181174.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@181174.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@181174.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@181174.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@181174.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@181316.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@181316.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@181316.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@181316.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@181316.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@181316.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@181316.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@181174.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@181316.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@181334.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@181330.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@181326.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@181325.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@181324.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@181323.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@181321.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@181320.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@181378.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@181377.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@181376.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@181375.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@181374.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@181373.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@181372.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@181371.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@181370.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@181369.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@181368.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@181366.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@181365.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@181364.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@181363.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@181362.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@181361.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@181360.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@181359.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@181358.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@181357.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@181356.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@181354.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@181353.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@181352.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@181351.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@181343.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@181338.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@181419.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@181418.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@181417.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@181416.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@181415.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@181414.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@181413.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@181412.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@181411.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@181410.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@181409.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@181407.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@181406.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@181405.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@181404.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@181403.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@181402.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@181401.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@181400.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@181399.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@181398.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@181397.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@181395.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@181394.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@181393.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@181392.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@181384.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@181379.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@181460.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@181459.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@181458.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@181457.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@181456.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@181455.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@181454.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@181453.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@181452.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@181451.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@181450.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@181448.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@181447.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@181446.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@181445.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@181444.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@181443.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@181442.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@181441.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@181440.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@181439.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@181438.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@181436.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@181435.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@181434.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@181433.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@181425.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@181420.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@181501.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@181500.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@181499.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@181498.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@181497.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@181496.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@181495.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@181494.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@181493.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@181492.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@181491.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@181489.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@181488.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@181487.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@181486.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@181485.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@181484.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@181483.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@181482.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@181481.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@181480.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@181479.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@181477.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@181476.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@181475.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@181474.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@181466.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@181461.4]
  assign accel_clock = clock; // @[:@181175.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@181176.4 Zynq.scala 54:17:@181790.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@181785.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@181778.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@181773.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@181757.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@181758.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@181759.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@181760.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@181761.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@181762.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@181763.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@181764.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@181765.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@181766.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@181767.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@181768.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@181769.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@181770.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@181771.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@181772.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@181756.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@181752.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@181747.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@181746.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@181745.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@181726.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@181710.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@181711.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@181712.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@181713.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@181714.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@181715.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@181716.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@181717.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@181718.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@181719.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@181720.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@181721.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@181722.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@181723.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@181724.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@181725.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@181709.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@181674.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@181673.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@181781.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@181780.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@181779.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@181667.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@181668.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@181671.4]
  assign FringeZynq_clock = clock; // @[:@181317.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@181318.4 Zynq.scala 53:18:@181789.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@181337.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@181336.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@181335.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@181333.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@181332.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@181331.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@181329.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@181328.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@181327.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@181322.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@181319.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@181367.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@181355.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@181350.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@181342.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@181339.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@181408.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@181396.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@181391.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@181383.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@181380.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@181449.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@181437.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@181432.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@181424.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@181421.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@181490.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@181478.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@181473.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@181465.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@181462.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@181786.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@181670.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@181669.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@181755.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@181754.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@181753.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@181751.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@181750.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@181749.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@181748.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@181784.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@181783.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@181782.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




