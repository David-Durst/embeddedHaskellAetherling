module FIFO(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  reg [7:0] _T__0; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_0;
  reg [7:0] _T__1; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_1;
  reg [7:0] _T__2; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_2;
  reg [7:0] _T__3; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_3;
  reg [7:0] _T__4; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_4;
  reg [7:0] _T__5; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_5;
  reg [7:0] _T__6; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_6;
  reg [7:0] _T__7; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_7;
  reg [7:0] _T__8; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_8;
  reg [7:0] _T__9; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_9;
  reg [7:0] _T__10; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_10;
  reg [7:0] _T__11; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_11;
  reg [7:0] _T__12; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_12;
  reg [7:0] _T__13; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_13;
  reg [7:0] _T__14; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_14;
  reg [7:0] _T__15; // @[FIFO.scala 13:26]
  reg [31:0] _RAND_15;
  reg  _T_1; // @[FIFO.scala 15:27]
  reg [31:0] _RAND_16;
  assign valid_down = _T_1; // @[FIFO.scala 16:16]
  assign O_0 = _T__0; // @[FIFO.scala 14:7]
  assign O_1 = _T__1; // @[FIFO.scala 14:7]
  assign O_2 = _T__2; // @[FIFO.scala 14:7]
  assign O_3 = _T__3; // @[FIFO.scala 14:7]
  assign O_4 = _T__4; // @[FIFO.scala 14:7]
  assign O_5 = _T__5; // @[FIFO.scala 14:7]
  assign O_6 = _T__6; // @[FIFO.scala 14:7]
  assign O_7 = _T__7; // @[FIFO.scala 14:7]
  assign O_8 = _T__8; // @[FIFO.scala 14:7]
  assign O_9 = _T__9; // @[FIFO.scala 14:7]
  assign O_10 = _T__10; // @[FIFO.scala 14:7]
  assign O_11 = _T__11; // @[FIFO.scala 14:7]
  assign O_12 = _T__12; // @[FIFO.scala 14:7]
  assign O_13 = _T__13; // @[FIFO.scala 14:7]
  assign O_14 = _T__14; // @[FIFO.scala 14:7]
  assign O_15 = _T__15; // @[FIFO.scala 14:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T__0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T__1 = _RAND_1[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T__2 = _RAND_2[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T__3 = _RAND_3[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T__4 = _RAND_4[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T__5 = _RAND_5[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T__6 = _RAND_6[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T__7 = _RAND_7[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T__8 = _RAND_8[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T__9 = _RAND_9[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T__10 = _RAND_10[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T__11 = _RAND_11[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T__12 = _RAND_12[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T__13 = _RAND_13[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T__14 = _RAND_14[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  _T__15 = _RAND_15[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  _T_1 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T__0 <= I_0;
    _T__1 <= I_1;
    _T__2 <= I_2;
    _T__3 <= I_3;
    _T__4 <= I_4;
    _T__5 <= I_5;
    _T__6 <= I_6;
    _T__7 <= I_7;
    _T__8 <= I_8;
    _T__9 <= I_9;
    _T__10 <= I_10;
    _T__11 <= I_11;
    _T__12 <= I_12;
    _T__13 <= I_13;
    _T__14 <= I_14;
    _T__15 <= I_15;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module NestedCounters(
  input   CE,
  output  valid
);
  assign valid = CE; // @[NestedCounters.scala 65:13]
endmodule
module NestedCountersWithNumValid(
  input   CE,
  output  valid
);
  wire  NestedCounters_CE; // @[NestedCounters.scala 20:44]
  wire  NestedCounters_valid; // @[NestedCounters.scala 20:44]
  NestedCounters NestedCounters ( // @[NestedCounters.scala 20:44]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign valid = NestedCounters_valid; // @[NestedCounters.scala 22:9]
  assign NestedCounters_CE = CE; // @[NestedCounters.scala 21:27]
endmodule
module RAM_ST(
  input        clock,
  input        RE,
  input  [6:0] RADDR,
  output [7:0] RDATA,
  input        WE,
  input  [6:0] WADDR,
  input  [7:0] WDATA
);
  wire  write_elem_counter_CE; // @[RAM_ST.scala 20:34]
  wire  write_elem_counter_valid; // @[RAM_ST.scala 20:34]
  wire  read_elem_counter_CE; // @[RAM_ST.scala 21:33]
  wire  read_elem_counter_valid; // @[RAM_ST.scala 21:33]
  reg [7:0] ram [0:119]; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_0;
  wire [7:0] ram__T_8_data; // @[RAM_ST.scala 29:24]
  wire [6:0] ram__T_8_addr; // @[RAM_ST.scala 29:24]
  reg [31:0] _RAND_1;
  wire [7:0] ram__T_2_data; // @[RAM_ST.scala 29:24]
  wire [6:0] ram__T_2_addr; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_mask; // @[RAM_ST.scala 29:24]
  wire  ram__T_2_en; // @[RAM_ST.scala 29:24]
  reg  ram__T_8_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [6:0] ram__T_8_addr_pipe_0;
  reg [31:0] _RAND_3;
  wire [6:0] _GEN_1; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_2; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_3; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_4; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_5; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_6; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_7; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_8; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_9; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_10; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_11; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_12; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_13; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_14; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_15; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_16; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_17; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_18; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_19; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_20; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_21; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_22; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_23; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_24; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_25; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_26; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_27; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_28; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_29; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_30; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_31; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_32; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_33; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_34; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_35; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_36; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_37; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_38; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_39; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_40; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_41; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_42; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_43; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_44; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_45; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_46; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_47; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_48; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_49; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_50; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_51; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_52; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_53; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_54; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_55; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_56; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_57; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_58; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_59; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_60; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_61; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_62; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_63; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_64; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_65; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_66; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_67; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_68; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_69; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_70; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_71; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_72; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_73; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_74; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_75; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_76; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_77; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_78; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_79; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_80; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_81; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_82; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_83; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_84; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_85; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_86; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_87; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_88; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_89; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_90; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_91; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_92; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_93; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_94; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_95; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_96; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_97; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_98; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_99; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_100; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_101; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_102; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_103; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_104; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_105; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_106; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_107; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_108; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_109; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_110; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_111; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_112; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_113; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_114; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_115; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_116; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_117; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_118; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_119; // @[RAM_ST.scala 31:71]
  wire [7:0] _T; // @[RAM_ST.scala 31:71]
  wire [6:0] _GEN_126; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_127; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_128; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_129; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_130; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_131; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_132; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_133; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_134; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_135; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_136; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_137; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_138; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_139; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_140; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_141; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_142; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_143; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_144; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_145; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_146; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_147; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_148; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_149; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_150; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_151; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_152; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_153; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_154; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_155; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_156; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_157; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_158; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_159; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_160; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_161; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_162; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_163; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_164; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_165; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_166; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_167; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_168; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_169; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_170; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_171; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_172; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_173; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_174; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_175; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_176; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_177; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_178; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_179; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_180; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_181; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_182; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_183; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_184; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_185; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_186; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_187; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_188; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_189; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_190; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_191; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_192; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_193; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_194; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_195; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_196; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_197; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_198; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_199; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_200; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_201; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_202; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_203; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_204; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_205; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_206; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_207; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_208; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_209; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_210; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_211; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_212; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_213; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_214; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_215; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_216; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_217; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_218; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_219; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_220; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_221; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_222; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_223; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_224; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_225; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_226; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_227; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_228; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_229; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_230; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_231; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_232; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_233; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_234; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_235; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_236; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_237; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_238; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_239; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_240; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_241; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_242; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_243; // @[RAM_ST.scala 32:46]
  wire [6:0] _GEN_244; // @[RAM_ST.scala 32:46]
  wire [7:0] _T_3; // @[RAM_ST.scala 32:46]
  NestedCountersWithNumValid write_elem_counter ( // @[RAM_ST.scala 20:34]
    .CE(write_elem_counter_CE),
    .valid(write_elem_counter_valid)
  );
  NestedCountersWithNumValid read_elem_counter ( // @[RAM_ST.scala 21:33]
    .CE(read_elem_counter_CE),
    .valid(read_elem_counter_valid)
  );
  assign ram__T_8_addr = ram__T_8_addr_pipe_0;
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_8_data = ram[ram__T_8_addr]; // @[RAM_ST.scala 29:24]
  `else
  assign ram__T_8_data = ram__T_8_addr >= 7'h78 ? _RAND_1[7:0] : ram[ram__T_8_addr]; // @[RAM_ST.scala 29:24]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign ram__T_2_data = WDATA;
  assign ram__T_2_addr = _T[6:0];
  assign ram__T_2_mask = 1'h1;
  assign ram__T_2_en = write_elem_counter_valid;
  assign _GEN_1 = 7'h1 == WADDR ? 7'h1 : 7'h0; // @[RAM_ST.scala 31:71]
  assign _GEN_2 = 7'h2 == WADDR ? 7'h2 : _GEN_1; // @[RAM_ST.scala 31:71]
  assign _GEN_3 = 7'h3 == WADDR ? 7'h3 : _GEN_2; // @[RAM_ST.scala 31:71]
  assign _GEN_4 = 7'h4 == WADDR ? 7'h4 : _GEN_3; // @[RAM_ST.scala 31:71]
  assign _GEN_5 = 7'h5 == WADDR ? 7'h5 : _GEN_4; // @[RAM_ST.scala 31:71]
  assign _GEN_6 = 7'h6 == WADDR ? 7'h6 : _GEN_5; // @[RAM_ST.scala 31:71]
  assign _GEN_7 = 7'h7 == WADDR ? 7'h7 : _GEN_6; // @[RAM_ST.scala 31:71]
  assign _GEN_8 = 7'h8 == WADDR ? 7'h8 : _GEN_7; // @[RAM_ST.scala 31:71]
  assign _GEN_9 = 7'h9 == WADDR ? 7'h9 : _GEN_8; // @[RAM_ST.scala 31:71]
  assign _GEN_10 = 7'ha == WADDR ? 7'ha : _GEN_9; // @[RAM_ST.scala 31:71]
  assign _GEN_11 = 7'hb == WADDR ? 7'hb : _GEN_10; // @[RAM_ST.scala 31:71]
  assign _GEN_12 = 7'hc == WADDR ? 7'hc : _GEN_11; // @[RAM_ST.scala 31:71]
  assign _GEN_13 = 7'hd == WADDR ? 7'hd : _GEN_12; // @[RAM_ST.scala 31:71]
  assign _GEN_14 = 7'he == WADDR ? 7'he : _GEN_13; // @[RAM_ST.scala 31:71]
  assign _GEN_15 = 7'hf == WADDR ? 7'hf : _GEN_14; // @[RAM_ST.scala 31:71]
  assign _GEN_16 = 7'h10 == WADDR ? 7'h10 : _GEN_15; // @[RAM_ST.scala 31:71]
  assign _GEN_17 = 7'h11 == WADDR ? 7'h11 : _GEN_16; // @[RAM_ST.scala 31:71]
  assign _GEN_18 = 7'h12 == WADDR ? 7'h12 : _GEN_17; // @[RAM_ST.scala 31:71]
  assign _GEN_19 = 7'h13 == WADDR ? 7'h13 : _GEN_18; // @[RAM_ST.scala 31:71]
  assign _GEN_20 = 7'h14 == WADDR ? 7'h14 : _GEN_19; // @[RAM_ST.scala 31:71]
  assign _GEN_21 = 7'h15 == WADDR ? 7'h15 : _GEN_20; // @[RAM_ST.scala 31:71]
  assign _GEN_22 = 7'h16 == WADDR ? 7'h16 : _GEN_21; // @[RAM_ST.scala 31:71]
  assign _GEN_23 = 7'h17 == WADDR ? 7'h17 : _GEN_22; // @[RAM_ST.scala 31:71]
  assign _GEN_24 = 7'h18 == WADDR ? 7'h18 : _GEN_23; // @[RAM_ST.scala 31:71]
  assign _GEN_25 = 7'h19 == WADDR ? 7'h19 : _GEN_24; // @[RAM_ST.scala 31:71]
  assign _GEN_26 = 7'h1a == WADDR ? 7'h1a : _GEN_25; // @[RAM_ST.scala 31:71]
  assign _GEN_27 = 7'h1b == WADDR ? 7'h1b : _GEN_26; // @[RAM_ST.scala 31:71]
  assign _GEN_28 = 7'h1c == WADDR ? 7'h1c : _GEN_27; // @[RAM_ST.scala 31:71]
  assign _GEN_29 = 7'h1d == WADDR ? 7'h1d : _GEN_28; // @[RAM_ST.scala 31:71]
  assign _GEN_30 = 7'h1e == WADDR ? 7'h1e : _GEN_29; // @[RAM_ST.scala 31:71]
  assign _GEN_31 = 7'h1f == WADDR ? 7'h1f : _GEN_30; // @[RAM_ST.scala 31:71]
  assign _GEN_32 = 7'h20 == WADDR ? 7'h20 : _GEN_31; // @[RAM_ST.scala 31:71]
  assign _GEN_33 = 7'h21 == WADDR ? 7'h21 : _GEN_32; // @[RAM_ST.scala 31:71]
  assign _GEN_34 = 7'h22 == WADDR ? 7'h22 : _GEN_33; // @[RAM_ST.scala 31:71]
  assign _GEN_35 = 7'h23 == WADDR ? 7'h23 : _GEN_34; // @[RAM_ST.scala 31:71]
  assign _GEN_36 = 7'h24 == WADDR ? 7'h24 : _GEN_35; // @[RAM_ST.scala 31:71]
  assign _GEN_37 = 7'h25 == WADDR ? 7'h25 : _GEN_36; // @[RAM_ST.scala 31:71]
  assign _GEN_38 = 7'h26 == WADDR ? 7'h26 : _GEN_37; // @[RAM_ST.scala 31:71]
  assign _GEN_39 = 7'h27 == WADDR ? 7'h27 : _GEN_38; // @[RAM_ST.scala 31:71]
  assign _GEN_40 = 7'h28 == WADDR ? 7'h28 : _GEN_39; // @[RAM_ST.scala 31:71]
  assign _GEN_41 = 7'h29 == WADDR ? 7'h29 : _GEN_40; // @[RAM_ST.scala 31:71]
  assign _GEN_42 = 7'h2a == WADDR ? 7'h2a : _GEN_41; // @[RAM_ST.scala 31:71]
  assign _GEN_43 = 7'h2b == WADDR ? 7'h2b : _GEN_42; // @[RAM_ST.scala 31:71]
  assign _GEN_44 = 7'h2c == WADDR ? 7'h2c : _GEN_43; // @[RAM_ST.scala 31:71]
  assign _GEN_45 = 7'h2d == WADDR ? 7'h2d : _GEN_44; // @[RAM_ST.scala 31:71]
  assign _GEN_46 = 7'h2e == WADDR ? 7'h2e : _GEN_45; // @[RAM_ST.scala 31:71]
  assign _GEN_47 = 7'h2f == WADDR ? 7'h2f : _GEN_46; // @[RAM_ST.scala 31:71]
  assign _GEN_48 = 7'h30 == WADDR ? 7'h30 : _GEN_47; // @[RAM_ST.scala 31:71]
  assign _GEN_49 = 7'h31 == WADDR ? 7'h31 : _GEN_48; // @[RAM_ST.scala 31:71]
  assign _GEN_50 = 7'h32 == WADDR ? 7'h32 : _GEN_49; // @[RAM_ST.scala 31:71]
  assign _GEN_51 = 7'h33 == WADDR ? 7'h33 : _GEN_50; // @[RAM_ST.scala 31:71]
  assign _GEN_52 = 7'h34 == WADDR ? 7'h34 : _GEN_51; // @[RAM_ST.scala 31:71]
  assign _GEN_53 = 7'h35 == WADDR ? 7'h35 : _GEN_52; // @[RAM_ST.scala 31:71]
  assign _GEN_54 = 7'h36 == WADDR ? 7'h36 : _GEN_53; // @[RAM_ST.scala 31:71]
  assign _GEN_55 = 7'h37 == WADDR ? 7'h37 : _GEN_54; // @[RAM_ST.scala 31:71]
  assign _GEN_56 = 7'h38 == WADDR ? 7'h38 : _GEN_55; // @[RAM_ST.scala 31:71]
  assign _GEN_57 = 7'h39 == WADDR ? 7'h39 : _GEN_56; // @[RAM_ST.scala 31:71]
  assign _GEN_58 = 7'h3a == WADDR ? 7'h3a : _GEN_57; // @[RAM_ST.scala 31:71]
  assign _GEN_59 = 7'h3b == WADDR ? 7'h3b : _GEN_58; // @[RAM_ST.scala 31:71]
  assign _GEN_60 = 7'h3c == WADDR ? 7'h3c : _GEN_59; // @[RAM_ST.scala 31:71]
  assign _GEN_61 = 7'h3d == WADDR ? 7'h3d : _GEN_60; // @[RAM_ST.scala 31:71]
  assign _GEN_62 = 7'h3e == WADDR ? 7'h3e : _GEN_61; // @[RAM_ST.scala 31:71]
  assign _GEN_63 = 7'h3f == WADDR ? 7'h3f : _GEN_62; // @[RAM_ST.scala 31:71]
  assign _GEN_64 = 7'h40 == WADDR ? 7'h40 : _GEN_63; // @[RAM_ST.scala 31:71]
  assign _GEN_65 = 7'h41 == WADDR ? 7'h41 : _GEN_64; // @[RAM_ST.scala 31:71]
  assign _GEN_66 = 7'h42 == WADDR ? 7'h42 : _GEN_65; // @[RAM_ST.scala 31:71]
  assign _GEN_67 = 7'h43 == WADDR ? 7'h43 : _GEN_66; // @[RAM_ST.scala 31:71]
  assign _GEN_68 = 7'h44 == WADDR ? 7'h44 : _GEN_67; // @[RAM_ST.scala 31:71]
  assign _GEN_69 = 7'h45 == WADDR ? 7'h45 : _GEN_68; // @[RAM_ST.scala 31:71]
  assign _GEN_70 = 7'h46 == WADDR ? 7'h46 : _GEN_69; // @[RAM_ST.scala 31:71]
  assign _GEN_71 = 7'h47 == WADDR ? 7'h47 : _GEN_70; // @[RAM_ST.scala 31:71]
  assign _GEN_72 = 7'h48 == WADDR ? 7'h48 : _GEN_71; // @[RAM_ST.scala 31:71]
  assign _GEN_73 = 7'h49 == WADDR ? 7'h49 : _GEN_72; // @[RAM_ST.scala 31:71]
  assign _GEN_74 = 7'h4a == WADDR ? 7'h4a : _GEN_73; // @[RAM_ST.scala 31:71]
  assign _GEN_75 = 7'h4b == WADDR ? 7'h4b : _GEN_74; // @[RAM_ST.scala 31:71]
  assign _GEN_76 = 7'h4c == WADDR ? 7'h4c : _GEN_75; // @[RAM_ST.scala 31:71]
  assign _GEN_77 = 7'h4d == WADDR ? 7'h4d : _GEN_76; // @[RAM_ST.scala 31:71]
  assign _GEN_78 = 7'h4e == WADDR ? 7'h4e : _GEN_77; // @[RAM_ST.scala 31:71]
  assign _GEN_79 = 7'h4f == WADDR ? 7'h4f : _GEN_78; // @[RAM_ST.scala 31:71]
  assign _GEN_80 = 7'h50 == WADDR ? 7'h50 : _GEN_79; // @[RAM_ST.scala 31:71]
  assign _GEN_81 = 7'h51 == WADDR ? 7'h51 : _GEN_80; // @[RAM_ST.scala 31:71]
  assign _GEN_82 = 7'h52 == WADDR ? 7'h52 : _GEN_81; // @[RAM_ST.scala 31:71]
  assign _GEN_83 = 7'h53 == WADDR ? 7'h53 : _GEN_82; // @[RAM_ST.scala 31:71]
  assign _GEN_84 = 7'h54 == WADDR ? 7'h54 : _GEN_83; // @[RAM_ST.scala 31:71]
  assign _GEN_85 = 7'h55 == WADDR ? 7'h55 : _GEN_84; // @[RAM_ST.scala 31:71]
  assign _GEN_86 = 7'h56 == WADDR ? 7'h56 : _GEN_85; // @[RAM_ST.scala 31:71]
  assign _GEN_87 = 7'h57 == WADDR ? 7'h57 : _GEN_86; // @[RAM_ST.scala 31:71]
  assign _GEN_88 = 7'h58 == WADDR ? 7'h58 : _GEN_87; // @[RAM_ST.scala 31:71]
  assign _GEN_89 = 7'h59 == WADDR ? 7'h59 : _GEN_88; // @[RAM_ST.scala 31:71]
  assign _GEN_90 = 7'h5a == WADDR ? 7'h5a : _GEN_89; // @[RAM_ST.scala 31:71]
  assign _GEN_91 = 7'h5b == WADDR ? 7'h5b : _GEN_90; // @[RAM_ST.scala 31:71]
  assign _GEN_92 = 7'h5c == WADDR ? 7'h5c : _GEN_91; // @[RAM_ST.scala 31:71]
  assign _GEN_93 = 7'h5d == WADDR ? 7'h5d : _GEN_92; // @[RAM_ST.scala 31:71]
  assign _GEN_94 = 7'h5e == WADDR ? 7'h5e : _GEN_93; // @[RAM_ST.scala 31:71]
  assign _GEN_95 = 7'h5f == WADDR ? 7'h5f : _GEN_94; // @[RAM_ST.scala 31:71]
  assign _GEN_96 = 7'h60 == WADDR ? 7'h60 : _GEN_95; // @[RAM_ST.scala 31:71]
  assign _GEN_97 = 7'h61 == WADDR ? 7'h61 : _GEN_96; // @[RAM_ST.scala 31:71]
  assign _GEN_98 = 7'h62 == WADDR ? 7'h62 : _GEN_97; // @[RAM_ST.scala 31:71]
  assign _GEN_99 = 7'h63 == WADDR ? 7'h63 : _GEN_98; // @[RAM_ST.scala 31:71]
  assign _GEN_100 = 7'h64 == WADDR ? 7'h64 : _GEN_99; // @[RAM_ST.scala 31:71]
  assign _GEN_101 = 7'h65 == WADDR ? 7'h65 : _GEN_100; // @[RAM_ST.scala 31:71]
  assign _GEN_102 = 7'h66 == WADDR ? 7'h66 : _GEN_101; // @[RAM_ST.scala 31:71]
  assign _GEN_103 = 7'h67 == WADDR ? 7'h67 : _GEN_102; // @[RAM_ST.scala 31:71]
  assign _GEN_104 = 7'h68 == WADDR ? 7'h68 : _GEN_103; // @[RAM_ST.scala 31:71]
  assign _GEN_105 = 7'h69 == WADDR ? 7'h69 : _GEN_104; // @[RAM_ST.scala 31:71]
  assign _GEN_106 = 7'h6a == WADDR ? 7'h6a : _GEN_105; // @[RAM_ST.scala 31:71]
  assign _GEN_107 = 7'h6b == WADDR ? 7'h6b : _GEN_106; // @[RAM_ST.scala 31:71]
  assign _GEN_108 = 7'h6c == WADDR ? 7'h6c : _GEN_107; // @[RAM_ST.scala 31:71]
  assign _GEN_109 = 7'h6d == WADDR ? 7'h6d : _GEN_108; // @[RAM_ST.scala 31:71]
  assign _GEN_110 = 7'h6e == WADDR ? 7'h6e : _GEN_109; // @[RAM_ST.scala 31:71]
  assign _GEN_111 = 7'h6f == WADDR ? 7'h6f : _GEN_110; // @[RAM_ST.scala 31:71]
  assign _GEN_112 = 7'h70 == WADDR ? 7'h70 : _GEN_111; // @[RAM_ST.scala 31:71]
  assign _GEN_113 = 7'h71 == WADDR ? 7'h71 : _GEN_112; // @[RAM_ST.scala 31:71]
  assign _GEN_114 = 7'h72 == WADDR ? 7'h72 : _GEN_113; // @[RAM_ST.scala 31:71]
  assign _GEN_115 = 7'h73 == WADDR ? 7'h73 : _GEN_114; // @[RAM_ST.scala 31:71]
  assign _GEN_116 = 7'h74 == WADDR ? 7'h74 : _GEN_115; // @[RAM_ST.scala 31:71]
  assign _GEN_117 = 7'h75 == WADDR ? 7'h75 : _GEN_116; // @[RAM_ST.scala 31:71]
  assign _GEN_118 = 7'h76 == WADDR ? 7'h76 : _GEN_117; // @[RAM_ST.scala 31:71]
  assign _GEN_119 = 7'h77 == WADDR ? 7'h77 : _GEN_118; // @[RAM_ST.scala 31:71]
  assign _T = {{1'd0}, _GEN_119}; // @[RAM_ST.scala 31:71]
  assign _GEN_126 = 7'h1 == RADDR ? 7'h1 : 7'h0; // @[RAM_ST.scala 32:46]
  assign _GEN_127 = 7'h2 == RADDR ? 7'h2 : _GEN_126; // @[RAM_ST.scala 32:46]
  assign _GEN_128 = 7'h3 == RADDR ? 7'h3 : _GEN_127; // @[RAM_ST.scala 32:46]
  assign _GEN_129 = 7'h4 == RADDR ? 7'h4 : _GEN_128; // @[RAM_ST.scala 32:46]
  assign _GEN_130 = 7'h5 == RADDR ? 7'h5 : _GEN_129; // @[RAM_ST.scala 32:46]
  assign _GEN_131 = 7'h6 == RADDR ? 7'h6 : _GEN_130; // @[RAM_ST.scala 32:46]
  assign _GEN_132 = 7'h7 == RADDR ? 7'h7 : _GEN_131; // @[RAM_ST.scala 32:46]
  assign _GEN_133 = 7'h8 == RADDR ? 7'h8 : _GEN_132; // @[RAM_ST.scala 32:46]
  assign _GEN_134 = 7'h9 == RADDR ? 7'h9 : _GEN_133; // @[RAM_ST.scala 32:46]
  assign _GEN_135 = 7'ha == RADDR ? 7'ha : _GEN_134; // @[RAM_ST.scala 32:46]
  assign _GEN_136 = 7'hb == RADDR ? 7'hb : _GEN_135; // @[RAM_ST.scala 32:46]
  assign _GEN_137 = 7'hc == RADDR ? 7'hc : _GEN_136; // @[RAM_ST.scala 32:46]
  assign _GEN_138 = 7'hd == RADDR ? 7'hd : _GEN_137; // @[RAM_ST.scala 32:46]
  assign _GEN_139 = 7'he == RADDR ? 7'he : _GEN_138; // @[RAM_ST.scala 32:46]
  assign _GEN_140 = 7'hf == RADDR ? 7'hf : _GEN_139; // @[RAM_ST.scala 32:46]
  assign _GEN_141 = 7'h10 == RADDR ? 7'h10 : _GEN_140; // @[RAM_ST.scala 32:46]
  assign _GEN_142 = 7'h11 == RADDR ? 7'h11 : _GEN_141; // @[RAM_ST.scala 32:46]
  assign _GEN_143 = 7'h12 == RADDR ? 7'h12 : _GEN_142; // @[RAM_ST.scala 32:46]
  assign _GEN_144 = 7'h13 == RADDR ? 7'h13 : _GEN_143; // @[RAM_ST.scala 32:46]
  assign _GEN_145 = 7'h14 == RADDR ? 7'h14 : _GEN_144; // @[RAM_ST.scala 32:46]
  assign _GEN_146 = 7'h15 == RADDR ? 7'h15 : _GEN_145; // @[RAM_ST.scala 32:46]
  assign _GEN_147 = 7'h16 == RADDR ? 7'h16 : _GEN_146; // @[RAM_ST.scala 32:46]
  assign _GEN_148 = 7'h17 == RADDR ? 7'h17 : _GEN_147; // @[RAM_ST.scala 32:46]
  assign _GEN_149 = 7'h18 == RADDR ? 7'h18 : _GEN_148; // @[RAM_ST.scala 32:46]
  assign _GEN_150 = 7'h19 == RADDR ? 7'h19 : _GEN_149; // @[RAM_ST.scala 32:46]
  assign _GEN_151 = 7'h1a == RADDR ? 7'h1a : _GEN_150; // @[RAM_ST.scala 32:46]
  assign _GEN_152 = 7'h1b == RADDR ? 7'h1b : _GEN_151; // @[RAM_ST.scala 32:46]
  assign _GEN_153 = 7'h1c == RADDR ? 7'h1c : _GEN_152; // @[RAM_ST.scala 32:46]
  assign _GEN_154 = 7'h1d == RADDR ? 7'h1d : _GEN_153; // @[RAM_ST.scala 32:46]
  assign _GEN_155 = 7'h1e == RADDR ? 7'h1e : _GEN_154; // @[RAM_ST.scala 32:46]
  assign _GEN_156 = 7'h1f == RADDR ? 7'h1f : _GEN_155; // @[RAM_ST.scala 32:46]
  assign _GEN_157 = 7'h20 == RADDR ? 7'h20 : _GEN_156; // @[RAM_ST.scala 32:46]
  assign _GEN_158 = 7'h21 == RADDR ? 7'h21 : _GEN_157; // @[RAM_ST.scala 32:46]
  assign _GEN_159 = 7'h22 == RADDR ? 7'h22 : _GEN_158; // @[RAM_ST.scala 32:46]
  assign _GEN_160 = 7'h23 == RADDR ? 7'h23 : _GEN_159; // @[RAM_ST.scala 32:46]
  assign _GEN_161 = 7'h24 == RADDR ? 7'h24 : _GEN_160; // @[RAM_ST.scala 32:46]
  assign _GEN_162 = 7'h25 == RADDR ? 7'h25 : _GEN_161; // @[RAM_ST.scala 32:46]
  assign _GEN_163 = 7'h26 == RADDR ? 7'h26 : _GEN_162; // @[RAM_ST.scala 32:46]
  assign _GEN_164 = 7'h27 == RADDR ? 7'h27 : _GEN_163; // @[RAM_ST.scala 32:46]
  assign _GEN_165 = 7'h28 == RADDR ? 7'h28 : _GEN_164; // @[RAM_ST.scala 32:46]
  assign _GEN_166 = 7'h29 == RADDR ? 7'h29 : _GEN_165; // @[RAM_ST.scala 32:46]
  assign _GEN_167 = 7'h2a == RADDR ? 7'h2a : _GEN_166; // @[RAM_ST.scala 32:46]
  assign _GEN_168 = 7'h2b == RADDR ? 7'h2b : _GEN_167; // @[RAM_ST.scala 32:46]
  assign _GEN_169 = 7'h2c == RADDR ? 7'h2c : _GEN_168; // @[RAM_ST.scala 32:46]
  assign _GEN_170 = 7'h2d == RADDR ? 7'h2d : _GEN_169; // @[RAM_ST.scala 32:46]
  assign _GEN_171 = 7'h2e == RADDR ? 7'h2e : _GEN_170; // @[RAM_ST.scala 32:46]
  assign _GEN_172 = 7'h2f == RADDR ? 7'h2f : _GEN_171; // @[RAM_ST.scala 32:46]
  assign _GEN_173 = 7'h30 == RADDR ? 7'h30 : _GEN_172; // @[RAM_ST.scala 32:46]
  assign _GEN_174 = 7'h31 == RADDR ? 7'h31 : _GEN_173; // @[RAM_ST.scala 32:46]
  assign _GEN_175 = 7'h32 == RADDR ? 7'h32 : _GEN_174; // @[RAM_ST.scala 32:46]
  assign _GEN_176 = 7'h33 == RADDR ? 7'h33 : _GEN_175; // @[RAM_ST.scala 32:46]
  assign _GEN_177 = 7'h34 == RADDR ? 7'h34 : _GEN_176; // @[RAM_ST.scala 32:46]
  assign _GEN_178 = 7'h35 == RADDR ? 7'h35 : _GEN_177; // @[RAM_ST.scala 32:46]
  assign _GEN_179 = 7'h36 == RADDR ? 7'h36 : _GEN_178; // @[RAM_ST.scala 32:46]
  assign _GEN_180 = 7'h37 == RADDR ? 7'h37 : _GEN_179; // @[RAM_ST.scala 32:46]
  assign _GEN_181 = 7'h38 == RADDR ? 7'h38 : _GEN_180; // @[RAM_ST.scala 32:46]
  assign _GEN_182 = 7'h39 == RADDR ? 7'h39 : _GEN_181; // @[RAM_ST.scala 32:46]
  assign _GEN_183 = 7'h3a == RADDR ? 7'h3a : _GEN_182; // @[RAM_ST.scala 32:46]
  assign _GEN_184 = 7'h3b == RADDR ? 7'h3b : _GEN_183; // @[RAM_ST.scala 32:46]
  assign _GEN_185 = 7'h3c == RADDR ? 7'h3c : _GEN_184; // @[RAM_ST.scala 32:46]
  assign _GEN_186 = 7'h3d == RADDR ? 7'h3d : _GEN_185; // @[RAM_ST.scala 32:46]
  assign _GEN_187 = 7'h3e == RADDR ? 7'h3e : _GEN_186; // @[RAM_ST.scala 32:46]
  assign _GEN_188 = 7'h3f == RADDR ? 7'h3f : _GEN_187; // @[RAM_ST.scala 32:46]
  assign _GEN_189 = 7'h40 == RADDR ? 7'h40 : _GEN_188; // @[RAM_ST.scala 32:46]
  assign _GEN_190 = 7'h41 == RADDR ? 7'h41 : _GEN_189; // @[RAM_ST.scala 32:46]
  assign _GEN_191 = 7'h42 == RADDR ? 7'h42 : _GEN_190; // @[RAM_ST.scala 32:46]
  assign _GEN_192 = 7'h43 == RADDR ? 7'h43 : _GEN_191; // @[RAM_ST.scala 32:46]
  assign _GEN_193 = 7'h44 == RADDR ? 7'h44 : _GEN_192; // @[RAM_ST.scala 32:46]
  assign _GEN_194 = 7'h45 == RADDR ? 7'h45 : _GEN_193; // @[RAM_ST.scala 32:46]
  assign _GEN_195 = 7'h46 == RADDR ? 7'h46 : _GEN_194; // @[RAM_ST.scala 32:46]
  assign _GEN_196 = 7'h47 == RADDR ? 7'h47 : _GEN_195; // @[RAM_ST.scala 32:46]
  assign _GEN_197 = 7'h48 == RADDR ? 7'h48 : _GEN_196; // @[RAM_ST.scala 32:46]
  assign _GEN_198 = 7'h49 == RADDR ? 7'h49 : _GEN_197; // @[RAM_ST.scala 32:46]
  assign _GEN_199 = 7'h4a == RADDR ? 7'h4a : _GEN_198; // @[RAM_ST.scala 32:46]
  assign _GEN_200 = 7'h4b == RADDR ? 7'h4b : _GEN_199; // @[RAM_ST.scala 32:46]
  assign _GEN_201 = 7'h4c == RADDR ? 7'h4c : _GEN_200; // @[RAM_ST.scala 32:46]
  assign _GEN_202 = 7'h4d == RADDR ? 7'h4d : _GEN_201; // @[RAM_ST.scala 32:46]
  assign _GEN_203 = 7'h4e == RADDR ? 7'h4e : _GEN_202; // @[RAM_ST.scala 32:46]
  assign _GEN_204 = 7'h4f == RADDR ? 7'h4f : _GEN_203; // @[RAM_ST.scala 32:46]
  assign _GEN_205 = 7'h50 == RADDR ? 7'h50 : _GEN_204; // @[RAM_ST.scala 32:46]
  assign _GEN_206 = 7'h51 == RADDR ? 7'h51 : _GEN_205; // @[RAM_ST.scala 32:46]
  assign _GEN_207 = 7'h52 == RADDR ? 7'h52 : _GEN_206; // @[RAM_ST.scala 32:46]
  assign _GEN_208 = 7'h53 == RADDR ? 7'h53 : _GEN_207; // @[RAM_ST.scala 32:46]
  assign _GEN_209 = 7'h54 == RADDR ? 7'h54 : _GEN_208; // @[RAM_ST.scala 32:46]
  assign _GEN_210 = 7'h55 == RADDR ? 7'h55 : _GEN_209; // @[RAM_ST.scala 32:46]
  assign _GEN_211 = 7'h56 == RADDR ? 7'h56 : _GEN_210; // @[RAM_ST.scala 32:46]
  assign _GEN_212 = 7'h57 == RADDR ? 7'h57 : _GEN_211; // @[RAM_ST.scala 32:46]
  assign _GEN_213 = 7'h58 == RADDR ? 7'h58 : _GEN_212; // @[RAM_ST.scala 32:46]
  assign _GEN_214 = 7'h59 == RADDR ? 7'h59 : _GEN_213; // @[RAM_ST.scala 32:46]
  assign _GEN_215 = 7'h5a == RADDR ? 7'h5a : _GEN_214; // @[RAM_ST.scala 32:46]
  assign _GEN_216 = 7'h5b == RADDR ? 7'h5b : _GEN_215; // @[RAM_ST.scala 32:46]
  assign _GEN_217 = 7'h5c == RADDR ? 7'h5c : _GEN_216; // @[RAM_ST.scala 32:46]
  assign _GEN_218 = 7'h5d == RADDR ? 7'h5d : _GEN_217; // @[RAM_ST.scala 32:46]
  assign _GEN_219 = 7'h5e == RADDR ? 7'h5e : _GEN_218; // @[RAM_ST.scala 32:46]
  assign _GEN_220 = 7'h5f == RADDR ? 7'h5f : _GEN_219; // @[RAM_ST.scala 32:46]
  assign _GEN_221 = 7'h60 == RADDR ? 7'h60 : _GEN_220; // @[RAM_ST.scala 32:46]
  assign _GEN_222 = 7'h61 == RADDR ? 7'h61 : _GEN_221; // @[RAM_ST.scala 32:46]
  assign _GEN_223 = 7'h62 == RADDR ? 7'h62 : _GEN_222; // @[RAM_ST.scala 32:46]
  assign _GEN_224 = 7'h63 == RADDR ? 7'h63 : _GEN_223; // @[RAM_ST.scala 32:46]
  assign _GEN_225 = 7'h64 == RADDR ? 7'h64 : _GEN_224; // @[RAM_ST.scala 32:46]
  assign _GEN_226 = 7'h65 == RADDR ? 7'h65 : _GEN_225; // @[RAM_ST.scala 32:46]
  assign _GEN_227 = 7'h66 == RADDR ? 7'h66 : _GEN_226; // @[RAM_ST.scala 32:46]
  assign _GEN_228 = 7'h67 == RADDR ? 7'h67 : _GEN_227; // @[RAM_ST.scala 32:46]
  assign _GEN_229 = 7'h68 == RADDR ? 7'h68 : _GEN_228; // @[RAM_ST.scala 32:46]
  assign _GEN_230 = 7'h69 == RADDR ? 7'h69 : _GEN_229; // @[RAM_ST.scala 32:46]
  assign _GEN_231 = 7'h6a == RADDR ? 7'h6a : _GEN_230; // @[RAM_ST.scala 32:46]
  assign _GEN_232 = 7'h6b == RADDR ? 7'h6b : _GEN_231; // @[RAM_ST.scala 32:46]
  assign _GEN_233 = 7'h6c == RADDR ? 7'h6c : _GEN_232; // @[RAM_ST.scala 32:46]
  assign _GEN_234 = 7'h6d == RADDR ? 7'h6d : _GEN_233; // @[RAM_ST.scala 32:46]
  assign _GEN_235 = 7'h6e == RADDR ? 7'h6e : _GEN_234; // @[RAM_ST.scala 32:46]
  assign _GEN_236 = 7'h6f == RADDR ? 7'h6f : _GEN_235; // @[RAM_ST.scala 32:46]
  assign _GEN_237 = 7'h70 == RADDR ? 7'h70 : _GEN_236; // @[RAM_ST.scala 32:46]
  assign _GEN_238 = 7'h71 == RADDR ? 7'h71 : _GEN_237; // @[RAM_ST.scala 32:46]
  assign _GEN_239 = 7'h72 == RADDR ? 7'h72 : _GEN_238; // @[RAM_ST.scala 32:46]
  assign _GEN_240 = 7'h73 == RADDR ? 7'h73 : _GEN_239; // @[RAM_ST.scala 32:46]
  assign _GEN_241 = 7'h74 == RADDR ? 7'h74 : _GEN_240; // @[RAM_ST.scala 32:46]
  assign _GEN_242 = 7'h75 == RADDR ? 7'h75 : _GEN_241; // @[RAM_ST.scala 32:46]
  assign _GEN_243 = 7'h76 == RADDR ? 7'h76 : _GEN_242; // @[RAM_ST.scala 32:46]
  assign _GEN_244 = 7'h77 == RADDR ? 7'h77 : _GEN_243; // @[RAM_ST.scala 32:46]
  assign _T_3 = {{1'd0}, _GEN_244}; // @[RAM_ST.scala 32:46]
  assign RDATA = ram__T_8_data; // @[RAM_ST.scala 32:9]
  assign write_elem_counter_CE = WE; // @[RAM_ST.scala 23:25]
  assign read_elem_counter_CE = RE; // @[RAM_ST.scala 24:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 120; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ram__T_8_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ram__T_8_addr_pipe_0 = _RAND_3[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram__T_2_en & ram__T_2_mask) begin
      ram[ram__T_2_addr] <= ram__T_2_data; // @[RAM_ST.scala 29:24]
    end
    ram__T_8_en_pipe_0 <= read_elem_counter_valid;
    if (read_elem_counter_valid) begin
      ram__T_8_addr_pipe_0 <= _T_3[6:0];
    end
  end
endmodule
module ShiftT(
  input        clock,
  input        reset,
  input        valid_up,
  input  [7:0] I,
  output [7:0] O
);
  wire  RAM_ST_clock; // @[ShiftT.scala 39:29]
  wire  RAM_ST_RE; // @[ShiftT.scala 39:29]
  wire [6:0] RAM_ST_RADDR; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_RDATA; // @[ShiftT.scala 39:29]
  wire  RAM_ST_WE; // @[ShiftT.scala 39:29]
  wire [6:0] RAM_ST_WADDR; // @[ShiftT.scala 39:29]
  wire [7:0] RAM_ST_WDATA; // @[ShiftT.scala 39:29]
  wire  NestedCounters_CE; // @[ShiftT.scala 41:31]
  wire  NestedCounters_valid; // @[ShiftT.scala 41:31]
  reg [6:0] value; // @[Counter.scala 29:33]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[Counter.scala 37:24]
  wire [6:0] _T_3; // @[Counter.scala 38:22]
  RAM_ST RAM_ST ( // @[ShiftT.scala 39:29]
    .clock(RAM_ST_clock),
    .RE(RAM_ST_RE),
    .RADDR(RAM_ST_RADDR),
    .RDATA(RAM_ST_RDATA),
    .WE(RAM_ST_WE),
    .WADDR(RAM_ST_WADDR),
    .WDATA(RAM_ST_WDATA)
  );
  NestedCounters NestedCounters ( // @[ShiftT.scala 41:31]
    .CE(NestedCounters_CE),
    .valid(NestedCounters_valid)
  );
  assign _T_1 = value == 7'h77; // @[Counter.scala 37:24]
  assign _T_3 = value + 7'h1; // @[Counter.scala 38:22]
  assign O = RAM_ST_RDATA; // @[ShiftT.scala 51:7]
  assign RAM_ST_clock = clock;
  assign RAM_ST_RE = valid_up; // @[ShiftT.scala 49:20]
  assign RAM_ST_RADDR = _T_1 ? 7'h0 : _T_3; // @[ShiftT.scala 46:76 ShiftT.scala 47:38]
  assign RAM_ST_WE = valid_up; // @[ShiftT.scala 48:20]
  assign RAM_ST_WADDR = value; // @[ShiftT.scala 45:23]
  assign RAM_ST_WDATA = I; // @[ShiftT.scala 50:23]
  assign NestedCounters_CE = valid_up; // @[ShiftT.scala 42:22]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[6:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 7'h0;
    end else if (valid_up) begin
      if (_T_1) begin
        value <= 7'h0;
      end else begin
        value <= _T_3;
      end
    end
  end
endmodule
module ShiftTS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_1_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_1_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_1_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_2_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_2_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_2_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_3_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_3_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_3_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_4_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_4_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_4_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_5_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_5_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_5_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_6_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_6_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_6_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_7_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_7_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_7_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_8_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_8_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_8_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_9_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_9_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_9_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_10_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_10_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_10_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_11_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_11_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_11_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_12_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_12_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_12_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_13_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_13_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_13_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_14_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_14_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_14_O; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_clock; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_reset; // @[ShiftTS.scala 32:34]
  wire  ShiftT_15_valid_up; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_15_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_15_O; // @[ShiftTS.scala 32:34]
  ShiftT ShiftT ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_clock),
    .reset(ShiftT_reset),
    .valid_up(ShiftT_valid_up),
    .I(ShiftT_I),
    .O(ShiftT_O)
  );
  ShiftT ShiftT_1 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_1_clock),
    .reset(ShiftT_1_reset),
    .valid_up(ShiftT_1_valid_up),
    .I(ShiftT_1_I),
    .O(ShiftT_1_O)
  );
  ShiftT ShiftT_2 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_2_clock),
    .reset(ShiftT_2_reset),
    .valid_up(ShiftT_2_valid_up),
    .I(ShiftT_2_I),
    .O(ShiftT_2_O)
  );
  ShiftT ShiftT_3 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_3_clock),
    .reset(ShiftT_3_reset),
    .valid_up(ShiftT_3_valid_up),
    .I(ShiftT_3_I),
    .O(ShiftT_3_O)
  );
  ShiftT ShiftT_4 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_4_clock),
    .reset(ShiftT_4_reset),
    .valid_up(ShiftT_4_valid_up),
    .I(ShiftT_4_I),
    .O(ShiftT_4_O)
  );
  ShiftT ShiftT_5 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_5_clock),
    .reset(ShiftT_5_reset),
    .valid_up(ShiftT_5_valid_up),
    .I(ShiftT_5_I),
    .O(ShiftT_5_O)
  );
  ShiftT ShiftT_6 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_6_clock),
    .reset(ShiftT_6_reset),
    .valid_up(ShiftT_6_valid_up),
    .I(ShiftT_6_I),
    .O(ShiftT_6_O)
  );
  ShiftT ShiftT_7 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_7_clock),
    .reset(ShiftT_7_reset),
    .valid_up(ShiftT_7_valid_up),
    .I(ShiftT_7_I),
    .O(ShiftT_7_O)
  );
  ShiftT ShiftT_8 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_8_clock),
    .reset(ShiftT_8_reset),
    .valid_up(ShiftT_8_valid_up),
    .I(ShiftT_8_I),
    .O(ShiftT_8_O)
  );
  ShiftT ShiftT_9 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_9_clock),
    .reset(ShiftT_9_reset),
    .valid_up(ShiftT_9_valid_up),
    .I(ShiftT_9_I),
    .O(ShiftT_9_O)
  );
  ShiftT ShiftT_10 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_10_clock),
    .reset(ShiftT_10_reset),
    .valid_up(ShiftT_10_valid_up),
    .I(ShiftT_10_I),
    .O(ShiftT_10_O)
  );
  ShiftT ShiftT_11 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_11_clock),
    .reset(ShiftT_11_reset),
    .valid_up(ShiftT_11_valid_up),
    .I(ShiftT_11_I),
    .O(ShiftT_11_O)
  );
  ShiftT ShiftT_12 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_12_clock),
    .reset(ShiftT_12_reset),
    .valid_up(ShiftT_12_valid_up),
    .I(ShiftT_12_I),
    .O(ShiftT_12_O)
  );
  ShiftT ShiftT_13 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_13_clock),
    .reset(ShiftT_13_reset),
    .valid_up(ShiftT_13_valid_up),
    .I(ShiftT_13_I),
    .O(ShiftT_13_O)
  );
  ShiftT ShiftT_14 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_14_clock),
    .reset(ShiftT_14_reset),
    .valid_up(ShiftT_14_valid_up),
    .I(ShiftT_14_I),
    .O(ShiftT_14_O)
  );
  ShiftT ShiftT_15 ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_15_clock),
    .reset(ShiftT_15_reset),
    .valid_up(ShiftT_15_valid_up),
    .I(ShiftT_15_I),
    .O(ShiftT_15_O)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 39:14]
  assign O_0 = ShiftT_O; // @[ShiftTS.scala 34:36]
  assign O_1 = ShiftT_1_O; // @[ShiftTS.scala 34:36]
  assign O_2 = ShiftT_2_O; // @[ShiftTS.scala 34:36]
  assign O_3 = ShiftT_3_O; // @[ShiftTS.scala 34:36]
  assign O_4 = ShiftT_4_O; // @[ShiftTS.scala 34:36]
  assign O_5 = ShiftT_5_O; // @[ShiftTS.scala 34:36]
  assign O_6 = ShiftT_6_O; // @[ShiftTS.scala 34:36]
  assign O_7 = ShiftT_7_O; // @[ShiftTS.scala 34:36]
  assign O_8 = ShiftT_8_O; // @[ShiftTS.scala 34:36]
  assign O_9 = ShiftT_9_O; // @[ShiftTS.scala 34:36]
  assign O_10 = ShiftT_10_O; // @[ShiftTS.scala 34:36]
  assign O_11 = ShiftT_11_O; // @[ShiftTS.scala 34:36]
  assign O_12 = ShiftT_12_O; // @[ShiftTS.scala 34:36]
  assign O_13 = ShiftT_13_O; // @[ShiftTS.scala 34:36]
  assign O_14 = ShiftT_14_O; // @[ShiftTS.scala 34:36]
  assign O_15 = ShiftT_15_O; // @[ShiftTS.scala 34:36]
  assign ShiftT_clock = clock;
  assign ShiftT_reset = reset;
  assign ShiftT_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_I = I_0; // @[ShiftTS.scala 33:24]
  assign ShiftT_1_clock = clock;
  assign ShiftT_1_reset = reset;
  assign ShiftT_1_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_1_I = I_1; // @[ShiftTS.scala 33:24]
  assign ShiftT_2_clock = clock;
  assign ShiftT_2_reset = reset;
  assign ShiftT_2_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_2_I = I_2; // @[ShiftTS.scala 33:24]
  assign ShiftT_3_clock = clock;
  assign ShiftT_3_reset = reset;
  assign ShiftT_3_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_3_I = I_3; // @[ShiftTS.scala 33:24]
  assign ShiftT_4_clock = clock;
  assign ShiftT_4_reset = reset;
  assign ShiftT_4_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_4_I = I_4; // @[ShiftTS.scala 33:24]
  assign ShiftT_5_clock = clock;
  assign ShiftT_5_reset = reset;
  assign ShiftT_5_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_5_I = I_5; // @[ShiftTS.scala 33:24]
  assign ShiftT_6_clock = clock;
  assign ShiftT_6_reset = reset;
  assign ShiftT_6_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_6_I = I_6; // @[ShiftTS.scala 33:24]
  assign ShiftT_7_clock = clock;
  assign ShiftT_7_reset = reset;
  assign ShiftT_7_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_7_I = I_7; // @[ShiftTS.scala 33:24]
  assign ShiftT_8_clock = clock;
  assign ShiftT_8_reset = reset;
  assign ShiftT_8_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_8_I = I_8; // @[ShiftTS.scala 33:24]
  assign ShiftT_9_clock = clock;
  assign ShiftT_9_reset = reset;
  assign ShiftT_9_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_9_I = I_9; // @[ShiftTS.scala 33:24]
  assign ShiftT_10_clock = clock;
  assign ShiftT_10_reset = reset;
  assign ShiftT_10_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_10_I = I_10; // @[ShiftTS.scala 33:24]
  assign ShiftT_11_clock = clock;
  assign ShiftT_11_reset = reset;
  assign ShiftT_11_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_11_I = I_11; // @[ShiftTS.scala 33:24]
  assign ShiftT_12_clock = clock;
  assign ShiftT_12_reset = reset;
  assign ShiftT_12_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_12_I = I_12; // @[ShiftTS.scala 33:24]
  assign ShiftT_13_clock = clock;
  assign ShiftT_13_reset = reset;
  assign ShiftT_13_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_13_I = I_13; // @[ShiftTS.scala 33:24]
  assign ShiftT_14_clock = clock;
  assign ShiftT_14_reset = reset;
  assign ShiftT_14_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_14_I = I_14; // @[ShiftTS.scala 33:24]
  assign ShiftT_15_clock = clock;
  assign ShiftT_15_reset = reset;
  assign ShiftT_15_valid_up = valid_up; // @[ShiftTS.scala 35:31]
  assign ShiftT_15_I = I_15; // @[ShiftTS.scala 33:24]
endmodule
module ShiftT_32(
  input        clock,
  input  [7:0] I,
  output [7:0] O
);
  reg [7:0] _T; // @[ShiftT.scala 24:82]
  reg [31:0] _RAND_0;
  assign O = _T; // @[ShiftT.scala 24:7]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= I;
  end
endmodule
module ShiftTS_2(
  input        clock,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  wire  ShiftT_clock; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_I; // @[ShiftTS.scala 32:34]
  wire [7:0] ShiftT_O; // @[ShiftTS.scala 32:34]
  ShiftT_32 ShiftT ( // @[ShiftTS.scala 32:34]
    .clock(ShiftT_clock),
    .I(ShiftT_I),
    .O(ShiftT_O)
  );
  assign valid_down = valid_up; // @[ShiftTS.scala 39:14]
  assign O_0 = ShiftT_O; // @[ShiftTS.scala 34:36]
  assign O_1 = I_0; // @[ShiftTS.scala 29:36]
  assign O_2 = I_1; // @[ShiftTS.scala 29:36]
  assign O_3 = I_2; // @[ShiftTS.scala 29:36]
  assign O_4 = I_3; // @[ShiftTS.scala 29:36]
  assign O_5 = I_4; // @[ShiftTS.scala 29:36]
  assign O_6 = I_5; // @[ShiftTS.scala 29:36]
  assign O_7 = I_6; // @[ShiftTS.scala 29:36]
  assign O_8 = I_7; // @[ShiftTS.scala 29:36]
  assign O_9 = I_8; // @[ShiftTS.scala 29:36]
  assign O_10 = I_9; // @[ShiftTS.scala 29:36]
  assign O_11 = I_10; // @[ShiftTS.scala 29:36]
  assign O_12 = I_11; // @[ShiftTS.scala 29:36]
  assign O_13 = I_12; // @[ShiftTS.scala 29:36]
  assign O_14 = I_13; // @[ShiftTS.scala 29:36]
  assign O_15 = I_14; // @[ShiftTS.scala 29:36]
  assign ShiftT_clock = clock;
  assign ShiftT_I = I_15; // @[ShiftTS.scala 33:24]
endmodule
module SSeqTupleCreator(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0 = I0; // @[Tuple.scala 12:32]
  assign O_1 = I1; // @[Tuple.scala 13:32]
endmodule
module Map2S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I0_3,
  input  [7:0] I0_4,
  input  [7:0] I0_5,
  input  [7:0] I0_6,
  input  [7:0] I0_7,
  input  [7:0] I0_8,
  input  [7:0] I0_9,
  input  [7:0] I0_10,
  input  [7:0] I0_11,
  input  [7:0] I0_12,
  input  [7:0] I0_13,
  input  [7:0] I0_14,
  input  [7:0] I0_15,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  input  [7:0] I1_3,
  input  [7:0] I1_4,
  input  [7:0] I1_5,
  input  [7:0] I1_6,
  input  [7:0] I1_7,
  input  [7:0] I1_8,
  input  [7:0] I1_9,
  input  [7:0] I1_10,
  input  [7:0] I1_11,
  input  [7:0] I1_12,
  input  [7:0] I1_13,
  input  [7:0] I1_14,
  input  [7:0] I1_15,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_15_0,
  output [7:0] O_15_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  SSeqTupleCreator other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  SSeqTupleCreator other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  SSeqTupleCreator other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0(other_ops_2_I0),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  SSeqTupleCreator other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0(other_ops_3_I0),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1)
  );
  SSeqTupleCreator other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0(other_ops_4_I0),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1)
  );
  SSeqTupleCreator other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0(other_ops_5_I0),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1)
  );
  SSeqTupleCreator other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0(other_ops_6_I0),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1)
  );
  SSeqTupleCreator other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0(other_ops_7_I0),
    .I1(other_ops_7_I1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1)
  );
  SSeqTupleCreator other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0(other_ops_8_I0),
    .I1(other_ops_8_I1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1)
  );
  SSeqTupleCreator other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0(other_ops_9_I0),
    .I1(other_ops_9_I1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1)
  );
  SSeqTupleCreator other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0(other_ops_10_I0),
    .I1(other_ops_10_I1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1)
  );
  SSeqTupleCreator other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0(other_ops_11_I0),
    .I1(other_ops_11_I1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1)
  );
  SSeqTupleCreator other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0(other_ops_12_I0),
    .I1(other_ops_12_I1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1)
  );
  SSeqTupleCreator other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0(other_ops_13_I0),
    .I1(other_ops_13_I1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1)
  );
  SSeqTupleCreator other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0(other_ops_14_I0),
    .I1(other_ops_14_I1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_8_0 = other_ops_7_O_0; // @[Map2S.scala 24:12]
  assign O_8_1 = other_ops_7_O_1; // @[Map2S.scala 24:12]
  assign O_9_0 = other_ops_8_O_0; // @[Map2S.scala 24:12]
  assign O_9_1 = other_ops_8_O_1; // @[Map2S.scala 24:12]
  assign O_10_0 = other_ops_9_O_0; // @[Map2S.scala 24:12]
  assign O_10_1 = other_ops_9_O_1; // @[Map2S.scala 24:12]
  assign O_11_0 = other_ops_10_O_0; // @[Map2S.scala 24:12]
  assign O_11_1 = other_ops_10_O_1; // @[Map2S.scala 24:12]
  assign O_12_0 = other_ops_11_O_0; // @[Map2S.scala 24:12]
  assign O_12_1 = other_ops_11_O_1; // @[Map2S.scala 24:12]
  assign O_13_0 = other_ops_12_O_0; // @[Map2S.scala 24:12]
  assign O_13_1 = other_ops_12_O_1; // @[Map2S.scala 24:12]
  assign O_14_0 = other_ops_13_O_0; // @[Map2S.scala 24:12]
  assign O_14_1 = other_ops_13_O_1; // @[Map2S.scala 24:12]
  assign O_15_0 = other_ops_14_O_0; // @[Map2S.scala 24:12]
  assign O_15_1 = other_ops_14_O_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0 = I0_3; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0 = I0_4; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0 = I0_5; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0 = I0_6; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0 = I0_7; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0 = I0_8; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0 = I0_9; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0 = I0_10; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0 = I0_11; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0 = I0_12; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0 = I0_13; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0 = I0_14; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0 = I0_15; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module Map2T(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I0_3,
  input  [7:0] I0_4,
  input  [7:0] I0_5,
  input  [7:0] I0_6,
  input  [7:0] I0_7,
  input  [7:0] I0_8,
  input  [7:0] I0_9,
  input  [7:0] I0_10,
  input  [7:0] I0_11,
  input  [7:0] I0_12,
  input  [7:0] I0_13,
  input  [7:0] I0_14,
  input  [7:0] I0_15,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  input  [7:0] I1_3,
  input  [7:0] I1_4,
  input  [7:0] I1_5,
  input  [7:0] I1_6,
  input  [7:0] I1_7,
  input  [7:0] I1_8,
  input  [7:0] I1_9,
  input  [7:0] I1_10,
  input  [7:0] I1_11,
  input  [7:0] I1_12,
  input  [7:0] I1_13,
  input  [7:0] I1_14,
  input  [7:0] I1_15,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_15_0,
  output [7:0] O_15_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1; // @[Map2T.scala 8:20]
  Map2S op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0(op_I0_0),
    .I0_1(op_I0_1),
    .I0_2(op_I0_2),
    .I0_3(op_I0_3),
    .I0_4(op_I0_4),
    .I0_5(op_I0_5),
    .I0_6(op_I0_6),
    .I0_7(op_I0_7),
    .I0_8(op_I0_8),
    .I0_9(op_I0_9),
    .I0_10(op_I0_10),
    .I0_11(op_I0_11),
    .I0_12(op_I0_12),
    .I0_13(op_I0_13),
    .I0_14(op_I0_14),
    .I0_15(op_I0_15),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .I1_8(op_I1_8),
    .I1_9(op_I1_9),
    .I1_10(op_I1_10),
    .I1_11(op_I1_11),
    .I1_12(op_I1_12),
    .I1_13(op_I1_13),
    .I1_14(op_I1_14),
    .I1_15(op_I1_15),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign O_8_0 = op_O_8_0; // @[Map2T.scala 17:7]
  assign O_8_1 = op_O_8_1; // @[Map2T.scala 17:7]
  assign O_9_0 = op_O_9_0; // @[Map2T.scala 17:7]
  assign O_9_1 = op_O_9_1; // @[Map2T.scala 17:7]
  assign O_10_0 = op_O_10_0; // @[Map2T.scala 17:7]
  assign O_10_1 = op_O_10_1; // @[Map2T.scala 17:7]
  assign O_11_0 = op_O_11_0; // @[Map2T.scala 17:7]
  assign O_11_1 = op_O_11_1; // @[Map2T.scala 17:7]
  assign O_12_0 = op_O_12_0; // @[Map2T.scala 17:7]
  assign O_12_1 = op_O_12_1; // @[Map2T.scala 17:7]
  assign O_13_0 = op_O_13_0; // @[Map2T.scala 17:7]
  assign O_13_1 = op_O_13_1; // @[Map2T.scala 17:7]
  assign O_14_0 = op_O_14_0; // @[Map2T.scala 17:7]
  assign O_14_1 = op_O_14_1; // @[Map2T.scala 17:7]
  assign O_15_0 = op_O_15_0; // @[Map2T.scala 17:7]
  assign O_15_1 = op_O_15_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0 = I0_0; // @[Map2T.scala 15:11]
  assign op_I0_1 = I0_1; // @[Map2T.scala 15:11]
  assign op_I0_2 = I0_2; // @[Map2T.scala 15:11]
  assign op_I0_3 = I0_3; // @[Map2T.scala 15:11]
  assign op_I0_4 = I0_4; // @[Map2T.scala 15:11]
  assign op_I0_5 = I0_5; // @[Map2T.scala 15:11]
  assign op_I0_6 = I0_6; // @[Map2T.scala 15:11]
  assign op_I0_7 = I0_7; // @[Map2T.scala 15:11]
  assign op_I0_8 = I0_8; // @[Map2T.scala 15:11]
  assign op_I0_9 = I0_9; // @[Map2T.scala 15:11]
  assign op_I0_10 = I0_10; // @[Map2T.scala 15:11]
  assign op_I0_11 = I0_11; // @[Map2T.scala 15:11]
  assign op_I0_12 = I0_12; // @[Map2T.scala 15:11]
  assign op_I0_13 = I0_13; // @[Map2T.scala 15:11]
  assign op_I0_14 = I0_14; // @[Map2T.scala 15:11]
  assign op_I0_15 = I0_15; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
  assign op_I1_8 = I1_8; // @[Map2T.scala 16:11]
  assign op_I1_9 = I1_9; // @[Map2T.scala 16:11]
  assign op_I1_10 = I1_10; // @[Map2T.scala 16:11]
  assign op_I1_11 = I1_11; // @[Map2T.scala 16:11]
  assign op_I1_12 = I1_12; // @[Map2T.scala 16:11]
  assign op_I1_13 = I1_13; // @[Map2T.scala 16:11]
  assign op_I1_14 = I1_14; // @[Map2T.scala 16:11]
  assign op_I1_15 = I1_15; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0 = I0_0; // @[Tuple.scala 24:34]
  assign O_1 = I0_1; // @[Tuple.scala 24:34]
  assign O_2 = I1; // @[Tuple.scala 26:32]
endmodule
module Map2S_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_3_0,
  input  [7:0] I0_3_1,
  input  [7:0] I0_4_0,
  input  [7:0] I0_4_1,
  input  [7:0] I0_5_0,
  input  [7:0] I0_5_1,
  input  [7:0] I0_6_0,
  input  [7:0] I0_6_1,
  input  [7:0] I0_7_0,
  input  [7:0] I0_7_1,
  input  [7:0] I0_8_0,
  input  [7:0] I0_8_1,
  input  [7:0] I0_9_0,
  input  [7:0] I0_9_1,
  input  [7:0] I0_10_0,
  input  [7:0] I0_10_1,
  input  [7:0] I0_11_0,
  input  [7:0] I0_11_1,
  input  [7:0] I0_12_0,
  input  [7:0] I0_12_1,
  input  [7:0] I0_13_0,
  input  [7:0] I0_13_1,
  input  [7:0] I0_14_0,
  input  [7:0] I0_14_1,
  input  [7:0] I0_15_0,
  input  [7:0] I0_15_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  input  [7:0] I1_3,
  input  [7:0] I1_4,
  input  [7:0] I1_5,
  input  [7:0] I1_6,
  input  [7:0] I1_7,
  input  [7:0] I1_8,
  input  [7:0] I1_9,
  input  [7:0] I1_10,
  input  [7:0] I1_11,
  input  [7:0] I1_12,
  input  [7:0] I1_13,
  input  [7:0] I1_14,
  input  [7:0] I1_15,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_3_2,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_4_2,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_5_2,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_6_2,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_7_2,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_8_2,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_9_2,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_10_2,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_11_2,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_12_2,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_13_2,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_14_2,
  output [7:0] O_15_0,
  output [7:0] O_15_1,
  output [7:0] O_15_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleAppender fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1(fst_op_I1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  SSeqTupleAppender other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1(other_ops_0_I1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  SSeqTupleAppender other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1(other_ops_1_I1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  SSeqTupleAppender other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1(other_ops_2_I1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  SSeqTupleAppender other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I1(other_ops_3_I1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  SSeqTupleAppender other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I1(other_ops_4_I1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  SSeqTupleAppender other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I1(other_ops_5_I1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  SSeqTupleAppender other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I1(other_ops_6_I1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  SSeqTupleAppender other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I1(other_ops_7_I1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1),
    .O_2(other_ops_7_O_2)
  );
  SSeqTupleAppender other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I1(other_ops_8_I1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1),
    .O_2(other_ops_8_O_2)
  );
  SSeqTupleAppender other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I1(other_ops_9_I1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1),
    .O_2(other_ops_9_O_2)
  );
  SSeqTupleAppender other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I1(other_ops_10_I1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1),
    .O_2(other_ops_10_O_2)
  );
  SSeqTupleAppender other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I1(other_ops_11_I1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1),
    .O_2(other_ops_11_O_2)
  );
  SSeqTupleAppender other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I1(other_ops_12_I1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1),
    .O_2(other_ops_12_O_2)
  );
  SSeqTupleAppender other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I1(other_ops_13_I1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1),
    .O_2(other_ops_13_O_2)
  );
  SSeqTupleAppender other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I1(other_ops_14_I1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1),
    .O_2(other_ops_14_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0 = fst_op_O_0; // @[Map2S.scala 19:8]
  assign O_0_1 = fst_op_O_1; // @[Map2S.scala 19:8]
  assign O_0_2 = fst_op_O_2; // @[Map2S.scala 19:8]
  assign O_1_0 = other_ops_0_O_0; // @[Map2S.scala 24:12]
  assign O_1_1 = other_ops_0_O_1; // @[Map2S.scala 24:12]
  assign O_1_2 = other_ops_0_O_2; // @[Map2S.scala 24:12]
  assign O_2_0 = other_ops_1_O_0; // @[Map2S.scala 24:12]
  assign O_2_1 = other_ops_1_O_1; // @[Map2S.scala 24:12]
  assign O_2_2 = other_ops_1_O_2; // @[Map2S.scala 24:12]
  assign O_3_0 = other_ops_2_O_0; // @[Map2S.scala 24:12]
  assign O_3_1 = other_ops_2_O_1; // @[Map2S.scala 24:12]
  assign O_3_2 = other_ops_2_O_2; // @[Map2S.scala 24:12]
  assign O_4_0 = other_ops_3_O_0; // @[Map2S.scala 24:12]
  assign O_4_1 = other_ops_3_O_1; // @[Map2S.scala 24:12]
  assign O_4_2 = other_ops_3_O_2; // @[Map2S.scala 24:12]
  assign O_5_0 = other_ops_4_O_0; // @[Map2S.scala 24:12]
  assign O_5_1 = other_ops_4_O_1; // @[Map2S.scala 24:12]
  assign O_5_2 = other_ops_4_O_2; // @[Map2S.scala 24:12]
  assign O_6_0 = other_ops_5_O_0; // @[Map2S.scala 24:12]
  assign O_6_1 = other_ops_5_O_1; // @[Map2S.scala 24:12]
  assign O_6_2 = other_ops_5_O_2; // @[Map2S.scala 24:12]
  assign O_7_0 = other_ops_6_O_0; // @[Map2S.scala 24:12]
  assign O_7_1 = other_ops_6_O_1; // @[Map2S.scala 24:12]
  assign O_7_2 = other_ops_6_O_2; // @[Map2S.scala 24:12]
  assign O_8_0 = other_ops_7_O_0; // @[Map2S.scala 24:12]
  assign O_8_1 = other_ops_7_O_1; // @[Map2S.scala 24:12]
  assign O_8_2 = other_ops_7_O_2; // @[Map2S.scala 24:12]
  assign O_9_0 = other_ops_8_O_0; // @[Map2S.scala 24:12]
  assign O_9_1 = other_ops_8_O_1; // @[Map2S.scala 24:12]
  assign O_9_2 = other_ops_8_O_2; // @[Map2S.scala 24:12]
  assign O_10_0 = other_ops_9_O_0; // @[Map2S.scala 24:12]
  assign O_10_1 = other_ops_9_O_1; // @[Map2S.scala 24:12]
  assign O_10_2 = other_ops_9_O_2; // @[Map2S.scala 24:12]
  assign O_11_0 = other_ops_10_O_0; // @[Map2S.scala 24:12]
  assign O_11_1 = other_ops_10_O_1; // @[Map2S.scala 24:12]
  assign O_11_2 = other_ops_10_O_2; // @[Map2S.scala 24:12]
  assign O_12_0 = other_ops_11_O_0; // @[Map2S.scala 24:12]
  assign O_12_1 = other_ops_11_O_1; // @[Map2S.scala 24:12]
  assign O_12_2 = other_ops_11_O_2; // @[Map2S.scala 24:12]
  assign O_13_0 = other_ops_12_O_0; // @[Map2S.scala 24:12]
  assign O_13_1 = other_ops_12_O_1; // @[Map2S.scala 24:12]
  assign O_13_2 = other_ops_12_O_2; // @[Map2S.scala 24:12]
  assign O_14_0 = other_ops_13_O_0; // @[Map2S.scala 24:12]
  assign O_14_1 = other_ops_13_O_1; // @[Map2S.scala 24:12]
  assign O_14_2 = other_ops_13_O_2; // @[Map2S.scala 24:12]
  assign O_15_0 = other_ops_14_O_0; // @[Map2S.scala 24:12]
  assign O_15_1 = other_ops_14_O_1; // @[Map2S.scala 24:12]
  assign O_15_2 = other_ops_14_O_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1 = I1_3; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1 = I1_4; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1 = I1_5; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1 = I1_6; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1 = I1_7; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I1 = I1_8; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I1 = I1_9; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I1 = I1_10; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I1 = I1_11; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I1 = I1_12; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I1 = I1_13; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I1 = I1_14; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I1 = I1_15; // @[Map2S.scala 23:43]
endmodule
module Map2T_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_3_0,
  input  [7:0] I0_3_1,
  input  [7:0] I0_4_0,
  input  [7:0] I0_4_1,
  input  [7:0] I0_5_0,
  input  [7:0] I0_5_1,
  input  [7:0] I0_6_0,
  input  [7:0] I0_6_1,
  input  [7:0] I0_7_0,
  input  [7:0] I0_7_1,
  input  [7:0] I0_8_0,
  input  [7:0] I0_8_1,
  input  [7:0] I0_9_0,
  input  [7:0] I0_9_1,
  input  [7:0] I0_10_0,
  input  [7:0] I0_10_1,
  input  [7:0] I0_11_0,
  input  [7:0] I0_11_1,
  input  [7:0] I0_12_0,
  input  [7:0] I0_12_1,
  input  [7:0] I0_13_0,
  input  [7:0] I0_13_1,
  input  [7:0] I0_14_0,
  input  [7:0] I0_14_1,
  input  [7:0] I0_15_0,
  input  [7:0] I0_15_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  input  [7:0] I1_3,
  input  [7:0] I1_4,
  input  [7:0] I1_5,
  input  [7:0] I1_6,
  input  [7:0] I1_7,
  input  [7:0] I1_8,
  input  [7:0] I1_9,
  input  [7:0] I1_10,
  input  [7:0] I1_11,
  input  [7:0] I1_12,
  input  [7:0] I1_13,
  input  [7:0] I1_14,
  input  [7:0] I1_15,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_3_2,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_4_2,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_5_2,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_6_2,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_7_2,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_8_2,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_9_2,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_10_2,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_11_2,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_12_2,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_13_2,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_14_2,
  output [7:0] O_15_0,
  output [7:0] O_15_1,
  output [7:0] O_15_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_2; // @[Map2T.scala 8:20]
  Map2S_1 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_8_0(op_I0_8_0),
    .I0_8_1(op_I0_8_1),
    .I0_9_0(op_I0_9_0),
    .I0_9_1(op_I0_9_1),
    .I0_10_0(op_I0_10_0),
    .I0_10_1(op_I0_10_1),
    .I0_11_0(op_I0_11_0),
    .I0_11_1(op_I0_11_1),
    .I0_12_0(op_I0_12_0),
    .I0_12_1(op_I0_12_1),
    .I0_13_0(op_I0_13_0),
    .I0_13_1(op_I0_13_1),
    .I0_14_0(op_I0_14_0),
    .I0_14_1(op_I0_14_1),
    .I0_15_0(op_I0_15_0),
    .I0_15_1(op_I0_15_1),
    .I1_0(op_I1_0),
    .I1_1(op_I1_1),
    .I1_2(op_I1_2),
    .I1_3(op_I1_3),
    .I1_4(op_I1_4),
    .I1_5(op_I1_5),
    .I1_6(op_I1_6),
    .I1_7(op_I1_7),
    .I1_8(op_I1_8),
    .I1_9(op_I1_9),
    .I1_10(op_I1_10),
    .I1_11(op_I1_11),
    .I1_12(op_I1_12),
    .I1_13(op_I1_13),
    .I1_14(op_I1_14),
    .I1_15(op_I1_15),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_8_2(op_O_8_2),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_9_2(op_O_9_2),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_10_2(op_O_10_2),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_11_2(op_O_11_2),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_12_2(op_O_12_2),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_13_2(op_O_13_2),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_14_2(op_O_14_2),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1),
    .O_15_2(op_O_15_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0 = op_O_0_0; // @[Map2T.scala 17:7]
  assign O_0_1 = op_O_0_1; // @[Map2T.scala 17:7]
  assign O_0_2 = op_O_0_2; // @[Map2T.scala 17:7]
  assign O_1_0 = op_O_1_0; // @[Map2T.scala 17:7]
  assign O_1_1 = op_O_1_1; // @[Map2T.scala 17:7]
  assign O_1_2 = op_O_1_2; // @[Map2T.scala 17:7]
  assign O_2_0 = op_O_2_0; // @[Map2T.scala 17:7]
  assign O_2_1 = op_O_2_1; // @[Map2T.scala 17:7]
  assign O_2_2 = op_O_2_2; // @[Map2T.scala 17:7]
  assign O_3_0 = op_O_3_0; // @[Map2T.scala 17:7]
  assign O_3_1 = op_O_3_1; // @[Map2T.scala 17:7]
  assign O_3_2 = op_O_3_2; // @[Map2T.scala 17:7]
  assign O_4_0 = op_O_4_0; // @[Map2T.scala 17:7]
  assign O_4_1 = op_O_4_1; // @[Map2T.scala 17:7]
  assign O_4_2 = op_O_4_2; // @[Map2T.scala 17:7]
  assign O_5_0 = op_O_5_0; // @[Map2T.scala 17:7]
  assign O_5_1 = op_O_5_1; // @[Map2T.scala 17:7]
  assign O_5_2 = op_O_5_2; // @[Map2T.scala 17:7]
  assign O_6_0 = op_O_6_0; // @[Map2T.scala 17:7]
  assign O_6_1 = op_O_6_1; // @[Map2T.scala 17:7]
  assign O_6_2 = op_O_6_2; // @[Map2T.scala 17:7]
  assign O_7_0 = op_O_7_0; // @[Map2T.scala 17:7]
  assign O_7_1 = op_O_7_1; // @[Map2T.scala 17:7]
  assign O_7_2 = op_O_7_2; // @[Map2T.scala 17:7]
  assign O_8_0 = op_O_8_0; // @[Map2T.scala 17:7]
  assign O_8_1 = op_O_8_1; // @[Map2T.scala 17:7]
  assign O_8_2 = op_O_8_2; // @[Map2T.scala 17:7]
  assign O_9_0 = op_O_9_0; // @[Map2T.scala 17:7]
  assign O_9_1 = op_O_9_1; // @[Map2T.scala 17:7]
  assign O_9_2 = op_O_9_2; // @[Map2T.scala 17:7]
  assign O_10_0 = op_O_10_0; // @[Map2T.scala 17:7]
  assign O_10_1 = op_O_10_1; // @[Map2T.scala 17:7]
  assign O_10_2 = op_O_10_2; // @[Map2T.scala 17:7]
  assign O_11_0 = op_O_11_0; // @[Map2T.scala 17:7]
  assign O_11_1 = op_O_11_1; // @[Map2T.scala 17:7]
  assign O_11_2 = op_O_11_2; // @[Map2T.scala 17:7]
  assign O_12_0 = op_O_12_0; // @[Map2T.scala 17:7]
  assign O_12_1 = op_O_12_1; // @[Map2T.scala 17:7]
  assign O_12_2 = op_O_12_2; // @[Map2T.scala 17:7]
  assign O_13_0 = op_O_13_0; // @[Map2T.scala 17:7]
  assign O_13_1 = op_O_13_1; // @[Map2T.scala 17:7]
  assign O_13_2 = op_O_13_2; // @[Map2T.scala 17:7]
  assign O_14_0 = op_O_14_0; // @[Map2T.scala 17:7]
  assign O_14_1 = op_O_14_1; // @[Map2T.scala 17:7]
  assign O_14_2 = op_O_14_2; // @[Map2T.scala 17:7]
  assign O_15_0 = op_O_15_0; // @[Map2T.scala 17:7]
  assign O_15_1 = op_O_15_1; // @[Map2T.scala 17:7]
  assign O_15_2 = op_O_15_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0 = I0_8_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1 = I0_8_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0 = I0_9_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1 = I0_9_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0 = I0_10_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1 = I0_10_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0 = I0_11_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1 = I0_11_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0 = I0_12_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1 = I0_12_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0 = I0_13_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1 = I0_13_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0 = I0_14_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1 = I0_14_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0 = I0_15_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1 = I0_15_1; // @[Map2T.scala 15:11]
  assign op_I1_0 = I1_0; // @[Map2T.scala 16:11]
  assign op_I1_1 = I1_1; // @[Map2T.scala 16:11]
  assign op_I1_2 = I1_2; // @[Map2T.scala 16:11]
  assign op_I1_3 = I1_3; // @[Map2T.scala 16:11]
  assign op_I1_4 = I1_4; // @[Map2T.scala 16:11]
  assign op_I1_5 = I1_5; // @[Map2T.scala 16:11]
  assign op_I1_6 = I1_6; // @[Map2T.scala 16:11]
  assign op_I1_7 = I1_7; // @[Map2T.scala 16:11]
  assign op_I1_8 = I1_8; // @[Map2T.scala 16:11]
  assign op_I1_9 = I1_9; // @[Map2T.scala 16:11]
  assign op_I1_10 = I1_10; // @[Map2T.scala 16:11]
  assign op_I1_11 = I1_11; // @[Map2T.scala 16:11]
  assign op_I1_12 = I1_12; // @[Map2T.scala 16:11]
  assign op_I1_13 = I1_13; // @[Map2T.scala 16:11]
  assign op_I1_14 = I1_14; // @[Map2T.scala 16:11]
  assign op_I1_15 = I1_15; // @[Map2T.scala 16:11]
endmodule
module PartitionS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  input  [7:0] I_3_0,
  input  [7:0] I_3_1,
  input  [7:0] I_3_2,
  input  [7:0] I_4_0,
  input  [7:0] I_4_1,
  input  [7:0] I_4_2,
  input  [7:0] I_5_0,
  input  [7:0] I_5_1,
  input  [7:0] I_5_2,
  input  [7:0] I_6_0,
  input  [7:0] I_6_1,
  input  [7:0] I_6_2,
  input  [7:0] I_7_0,
  input  [7:0] I_7_1,
  input  [7:0] I_7_2,
  input  [7:0] I_8_0,
  input  [7:0] I_8_1,
  input  [7:0] I_8_2,
  input  [7:0] I_9_0,
  input  [7:0] I_9_1,
  input  [7:0] I_9_2,
  input  [7:0] I_10_0,
  input  [7:0] I_10_1,
  input  [7:0] I_10_2,
  input  [7:0] I_11_0,
  input  [7:0] I_11_1,
  input  [7:0] I_11_2,
  input  [7:0] I_12_0,
  input  [7:0] I_12_1,
  input  [7:0] I_12_2,
  input  [7:0] I_13_0,
  input  [7:0] I_13_1,
  input  [7:0] I_13_2,
  input  [7:0] I_14_0,
  input  [7:0] I_14_1,
  input  [7:0] I_14_2,
  input  [7:0] I_15_0,
  input  [7:0] I_15_1,
  input  [7:0] I_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_0_0_2 = I_0_2; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_1_0_2 = I_1_2; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2 = I_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
  assign O_3_0_2 = I_3_2; // @[Partition.scala 15:39]
  assign O_4_0_0 = I_4_0; // @[Partition.scala 15:39]
  assign O_4_0_1 = I_4_1; // @[Partition.scala 15:39]
  assign O_4_0_2 = I_4_2; // @[Partition.scala 15:39]
  assign O_5_0_0 = I_5_0; // @[Partition.scala 15:39]
  assign O_5_0_1 = I_5_1; // @[Partition.scala 15:39]
  assign O_5_0_2 = I_5_2; // @[Partition.scala 15:39]
  assign O_6_0_0 = I_6_0; // @[Partition.scala 15:39]
  assign O_6_0_1 = I_6_1; // @[Partition.scala 15:39]
  assign O_6_0_2 = I_6_2; // @[Partition.scala 15:39]
  assign O_7_0_0 = I_7_0; // @[Partition.scala 15:39]
  assign O_7_0_1 = I_7_1; // @[Partition.scala 15:39]
  assign O_7_0_2 = I_7_2; // @[Partition.scala 15:39]
  assign O_8_0_0 = I_8_0; // @[Partition.scala 15:39]
  assign O_8_0_1 = I_8_1; // @[Partition.scala 15:39]
  assign O_8_0_2 = I_8_2; // @[Partition.scala 15:39]
  assign O_9_0_0 = I_9_0; // @[Partition.scala 15:39]
  assign O_9_0_1 = I_9_1; // @[Partition.scala 15:39]
  assign O_9_0_2 = I_9_2; // @[Partition.scala 15:39]
  assign O_10_0_0 = I_10_0; // @[Partition.scala 15:39]
  assign O_10_0_1 = I_10_1; // @[Partition.scala 15:39]
  assign O_10_0_2 = I_10_2; // @[Partition.scala 15:39]
  assign O_11_0_0 = I_11_0; // @[Partition.scala 15:39]
  assign O_11_0_1 = I_11_1; // @[Partition.scala 15:39]
  assign O_11_0_2 = I_11_2; // @[Partition.scala 15:39]
  assign O_12_0_0 = I_12_0; // @[Partition.scala 15:39]
  assign O_12_0_1 = I_12_1; // @[Partition.scala 15:39]
  assign O_12_0_2 = I_12_2; // @[Partition.scala 15:39]
  assign O_13_0_0 = I_13_0; // @[Partition.scala 15:39]
  assign O_13_0_1 = I_13_1; // @[Partition.scala 15:39]
  assign O_13_0_2 = I_13_2; // @[Partition.scala 15:39]
  assign O_14_0_0 = I_14_0; // @[Partition.scala 15:39]
  assign O_14_0_1 = I_14_1; // @[Partition.scala 15:39]
  assign O_14_0_2 = I_14_2; // @[Partition.scala 15:39]
  assign O_15_0_0 = I_15_0; // @[Partition.scala 15:39]
  assign O_15_0_1 = I_15_1; // @[Partition.scala 15:39]
  assign O_15_0_2 = I_15_2; // @[Partition.scala 15:39]
endmodule
module MapT(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  input  [7:0] I_3_0,
  input  [7:0] I_3_1,
  input  [7:0] I_3_2,
  input  [7:0] I_4_0,
  input  [7:0] I_4_1,
  input  [7:0] I_4_2,
  input  [7:0] I_5_0,
  input  [7:0] I_5_1,
  input  [7:0] I_5_2,
  input  [7:0] I_6_0,
  input  [7:0] I_6_1,
  input  [7:0] I_6_2,
  input  [7:0] I_7_0,
  input  [7:0] I_7_1,
  input  [7:0] I_7_2,
  input  [7:0] I_8_0,
  input  [7:0] I_8_1,
  input  [7:0] I_8_2,
  input  [7:0] I_9_0,
  input  [7:0] I_9_1,
  input  [7:0] I_9_2,
  input  [7:0] I_10_0,
  input  [7:0] I_10_1,
  input  [7:0] I_10_2,
  input  [7:0] I_11_0,
  input  [7:0] I_11_1,
  input  [7:0] I_11_2,
  input  [7:0] I_12_0,
  input  [7:0] I_12_1,
  input  [7:0] I_12_2,
  input  [7:0] I_13_0,
  input  [7:0] I_13_1,
  input  [7:0] I_13_2,
  input  [7:0] I_14_0,
  input  [7:0] I_14_1,
  input  [7:0] I_14_2,
  input  [7:0] I_15_0,
  input  [7:0] I_15_1,
  input  [7:0] I_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_2; // @[MapT.scala 8:20]
  PartitionS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_0_2(op_I_0_2),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_1_2(op_I_1_2),
    .I_2_0(op_I_2_0),
    .I_2_1(op_I_2_1),
    .I_2_2(op_I_2_2),
    .I_3_0(op_I_3_0),
    .I_3_1(op_I_3_1),
    .I_3_2(op_I_3_2),
    .I_4_0(op_I_4_0),
    .I_4_1(op_I_4_1),
    .I_4_2(op_I_4_2),
    .I_5_0(op_I_5_0),
    .I_5_1(op_I_5_1),
    .I_5_2(op_I_5_2),
    .I_6_0(op_I_6_0),
    .I_6_1(op_I_6_1),
    .I_6_2(op_I_6_2),
    .I_7_0(op_I_7_0),
    .I_7_1(op_I_7_1),
    .I_7_2(op_I_7_2),
    .I_8_0(op_I_8_0),
    .I_8_1(op_I_8_1),
    .I_8_2(op_I_8_2),
    .I_9_0(op_I_9_0),
    .I_9_1(op_I_9_1),
    .I_9_2(op_I_9_2),
    .I_10_0(op_I_10_0),
    .I_10_1(op_I_10_1),
    .I_10_2(op_I_10_2),
    .I_11_0(op_I_11_0),
    .I_11_1(op_I_11_1),
    .I_11_2(op_I_11_2),
    .I_12_0(op_I_12_0),
    .I_12_1(op_I_12_1),
    .I_12_2(op_I_12_2),
    .I_13_0(op_I_13_0),
    .I_13_1(op_I_13_1),
    .I_13_2(op_I_13_2),
    .I_14_0(op_I_14_0),
    .I_14_1(op_I_14_1),
    .I_14_2(op_I_14_2),
    .I_15_0(op_I_15_0),
    .I_15_1(op_I_15_1),
    .I_15_2(op_I_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_0_2 = op_O_8_0_2; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_0_2 = op_O_9_0_2; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_0_2 = op_O_10_0_2; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_0_2 = op_O_11_0_2; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_0_2 = op_O_12_0_2; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_0_2 = op_O_13_0_2; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_0_2 = op_O_14_0_2; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_0_2 = op_O_15_0_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_0_2 = I_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_1_2 = I_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0 = I_2_0; // @[MapT.scala 14:10]
  assign op_I_2_1 = I_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2 = I_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0 = I_3_0; // @[MapT.scala 14:10]
  assign op_I_3_1 = I_3_1; // @[MapT.scala 14:10]
  assign op_I_3_2 = I_3_2; // @[MapT.scala 14:10]
  assign op_I_4_0 = I_4_0; // @[MapT.scala 14:10]
  assign op_I_4_1 = I_4_1; // @[MapT.scala 14:10]
  assign op_I_4_2 = I_4_2; // @[MapT.scala 14:10]
  assign op_I_5_0 = I_5_0; // @[MapT.scala 14:10]
  assign op_I_5_1 = I_5_1; // @[MapT.scala 14:10]
  assign op_I_5_2 = I_5_2; // @[MapT.scala 14:10]
  assign op_I_6_0 = I_6_0; // @[MapT.scala 14:10]
  assign op_I_6_1 = I_6_1; // @[MapT.scala 14:10]
  assign op_I_6_2 = I_6_2; // @[MapT.scala 14:10]
  assign op_I_7_0 = I_7_0; // @[MapT.scala 14:10]
  assign op_I_7_1 = I_7_1; // @[MapT.scala 14:10]
  assign op_I_7_2 = I_7_2; // @[MapT.scala 14:10]
  assign op_I_8_0 = I_8_0; // @[MapT.scala 14:10]
  assign op_I_8_1 = I_8_1; // @[MapT.scala 14:10]
  assign op_I_8_2 = I_8_2; // @[MapT.scala 14:10]
  assign op_I_9_0 = I_9_0; // @[MapT.scala 14:10]
  assign op_I_9_1 = I_9_1; // @[MapT.scala 14:10]
  assign op_I_9_2 = I_9_2; // @[MapT.scala 14:10]
  assign op_I_10_0 = I_10_0; // @[MapT.scala 14:10]
  assign op_I_10_1 = I_10_1; // @[MapT.scala 14:10]
  assign op_I_10_2 = I_10_2; // @[MapT.scala 14:10]
  assign op_I_11_0 = I_11_0; // @[MapT.scala 14:10]
  assign op_I_11_1 = I_11_1; // @[MapT.scala 14:10]
  assign op_I_11_2 = I_11_2; // @[MapT.scala 14:10]
  assign op_I_12_0 = I_12_0; // @[MapT.scala 14:10]
  assign op_I_12_1 = I_12_1; // @[MapT.scala 14:10]
  assign op_I_12_2 = I_12_2; // @[MapT.scala 14:10]
  assign op_I_13_0 = I_13_0; // @[MapT.scala 14:10]
  assign op_I_13_1 = I_13_1; // @[MapT.scala 14:10]
  assign op_I_13_2 = I_13_2; // @[MapT.scala 14:10]
  assign op_I_14_0 = I_14_0; // @[MapT.scala 14:10]
  assign op_I_14_1 = I_14_1; // @[MapT.scala 14:10]
  assign op_I_14_2 = I_14_2; // @[MapT.scala 14:10]
  assign op_I_15_0 = I_15_0; // @[MapT.scala 14:10]
  assign op_I_15_1 = I_15_1; // @[MapT.scala 14:10]
  assign op_I_15_2 = I_15_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
  assign O_2 = I_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .I_2(op_inst_I_2),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1),
    .O_2(op_inst_O_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign O_2 = op_inst_O_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2 = I_0_2; // @[Remove1S.scala 13:13]
endmodule
module MapS(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_3_2,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_4_2,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_5_2,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_6_2,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_7_2,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_8_2,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_9_2,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_10_2,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_11_2,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_12_2,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_13_2,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_14_2,
  output [7:0] O_15_0,
  output [7:0] O_15_1,
  output [7:0] O_15_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  Remove1S other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  Remove1S other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  Remove1S other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1),
    .O_2(other_ops_2_O_2)
  );
  Remove1S other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1),
    .O_2(other_ops_3_O_2)
  );
  Remove1S other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1),
    .O_2(other_ops_4_O_2)
  );
  Remove1S other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1),
    .O_2(other_ops_5_O_2)
  );
  Remove1S other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1),
    .O_2(other_ops_6_O_2)
  );
  Remove1S other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_0_2(other_ops_7_I_0_2),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1),
    .O_2(other_ops_7_O_2)
  );
  Remove1S other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_0_2(other_ops_8_I_0_2),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1),
    .O_2(other_ops_8_O_2)
  );
  Remove1S other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_0_2(other_ops_9_I_0_2),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1),
    .O_2(other_ops_9_O_2)
  );
  Remove1S other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_0_2(other_ops_10_I_0_2),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1),
    .O_2(other_ops_10_O_2)
  );
  Remove1S other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_0_2(other_ops_11_I_0_2),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1),
    .O_2(other_ops_11_O_2)
  );
  Remove1S other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_0_2(other_ops_12_I_0_2),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1),
    .O_2(other_ops_12_O_2)
  );
  Remove1S other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_0_2(other_ops_13_I_0_2),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1),
    .O_2(other_ops_13_O_2)
  );
  Remove1S other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_0_2(other_ops_14_I_0_2),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1),
    .O_2(other_ops_14_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign O_3_2 = other_ops_2_O_2; // @[MapS.scala 21:12]
  assign O_4_0 = other_ops_3_O_0; // @[MapS.scala 21:12]
  assign O_4_1 = other_ops_3_O_1; // @[MapS.scala 21:12]
  assign O_4_2 = other_ops_3_O_2; // @[MapS.scala 21:12]
  assign O_5_0 = other_ops_4_O_0; // @[MapS.scala 21:12]
  assign O_5_1 = other_ops_4_O_1; // @[MapS.scala 21:12]
  assign O_5_2 = other_ops_4_O_2; // @[MapS.scala 21:12]
  assign O_6_0 = other_ops_5_O_0; // @[MapS.scala 21:12]
  assign O_6_1 = other_ops_5_O_1; // @[MapS.scala 21:12]
  assign O_6_2 = other_ops_5_O_2; // @[MapS.scala 21:12]
  assign O_7_0 = other_ops_6_O_0; // @[MapS.scala 21:12]
  assign O_7_1 = other_ops_6_O_1; // @[MapS.scala 21:12]
  assign O_7_2 = other_ops_6_O_2; // @[MapS.scala 21:12]
  assign O_8_0 = other_ops_7_O_0; // @[MapS.scala 21:12]
  assign O_8_1 = other_ops_7_O_1; // @[MapS.scala 21:12]
  assign O_8_2 = other_ops_7_O_2; // @[MapS.scala 21:12]
  assign O_9_0 = other_ops_8_O_0; // @[MapS.scala 21:12]
  assign O_9_1 = other_ops_8_O_1; // @[MapS.scala 21:12]
  assign O_9_2 = other_ops_8_O_2; // @[MapS.scala 21:12]
  assign O_10_0 = other_ops_9_O_0; // @[MapS.scala 21:12]
  assign O_10_1 = other_ops_9_O_1; // @[MapS.scala 21:12]
  assign O_10_2 = other_ops_9_O_2; // @[MapS.scala 21:12]
  assign O_11_0 = other_ops_10_O_0; // @[MapS.scala 21:12]
  assign O_11_1 = other_ops_10_O_1; // @[MapS.scala 21:12]
  assign O_11_2 = other_ops_10_O_2; // @[MapS.scala 21:12]
  assign O_12_0 = other_ops_11_O_0; // @[MapS.scala 21:12]
  assign O_12_1 = other_ops_11_O_1; // @[MapS.scala 21:12]
  assign O_12_2 = other_ops_11_O_2; // @[MapS.scala 21:12]
  assign O_13_0 = other_ops_12_O_0; // @[MapS.scala 21:12]
  assign O_13_1 = other_ops_12_O_1; // @[MapS.scala 21:12]
  assign O_13_2 = other_ops_12_O_2; // @[MapS.scala 21:12]
  assign O_14_0 = other_ops_13_O_0; // @[MapS.scala 21:12]
  assign O_14_1 = other_ops_13_O_1; // @[MapS.scala 21:12]
  assign O_14_2 = other_ops_13_O_2; // @[MapS.scala 21:12]
  assign O_15_0 = other_ops_14_O_0; // @[MapS.scala 21:12]
  assign O_15_1 = other_ops_14_O_1; // @[MapS.scala 21:12]
  assign O_15_2 = other_ops_14_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2 = I_8_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2 = I_9_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2 = I_10_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2 = I_11_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2 = I_12_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2 = I_13_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2 = I_14_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2 = I_15_0_2; // @[MapS.scala 20:41]
endmodule
module MapT_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_3_2,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_4_2,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_5_2,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_6_2,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_7_2,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_8_2,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_9_2,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_10_2,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_11_2,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_12_2,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_13_2,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_14_2,
  output [7:0] O_15_0,
  output [7:0] O_15_1,
  output [7:0] O_15_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_2; // @[MapT.scala 8:20]
  MapS op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_0_2(op_O_0_2),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_1_2(op_O_1_2),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_2_2(op_O_2_2),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_3_2(op_O_3_2),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_4_2(op_O_4_2),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_5_2(op_O_5_2),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_6_2(op_O_6_2),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_7_2(op_O_7_2),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_8_2(op_O_8_2),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_9_2(op_O_9_2),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_10_2(op_O_10_2),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_11_2(op_O_11_2),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_12_2(op_O_12_2),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_13_2(op_O_13_2),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_14_2(op_O_14_2),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1),
    .O_15_2(op_O_15_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_0_2 = op_O_0_2; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_1_2 = op_O_1_2; // @[MapT.scala 15:7]
  assign O_2_0 = op_O_2_0; // @[MapT.scala 15:7]
  assign O_2_1 = op_O_2_1; // @[MapT.scala 15:7]
  assign O_2_2 = op_O_2_2; // @[MapT.scala 15:7]
  assign O_3_0 = op_O_3_0; // @[MapT.scala 15:7]
  assign O_3_1 = op_O_3_1; // @[MapT.scala 15:7]
  assign O_3_2 = op_O_3_2; // @[MapT.scala 15:7]
  assign O_4_0 = op_O_4_0; // @[MapT.scala 15:7]
  assign O_4_1 = op_O_4_1; // @[MapT.scala 15:7]
  assign O_4_2 = op_O_4_2; // @[MapT.scala 15:7]
  assign O_5_0 = op_O_5_0; // @[MapT.scala 15:7]
  assign O_5_1 = op_O_5_1; // @[MapT.scala 15:7]
  assign O_5_2 = op_O_5_2; // @[MapT.scala 15:7]
  assign O_6_0 = op_O_6_0; // @[MapT.scala 15:7]
  assign O_6_1 = op_O_6_1; // @[MapT.scala 15:7]
  assign O_6_2 = op_O_6_2; // @[MapT.scala 15:7]
  assign O_7_0 = op_O_7_0; // @[MapT.scala 15:7]
  assign O_7_1 = op_O_7_1; // @[MapT.scala 15:7]
  assign O_7_2 = op_O_7_2; // @[MapT.scala 15:7]
  assign O_8_0 = op_O_8_0; // @[MapT.scala 15:7]
  assign O_8_1 = op_O_8_1; // @[MapT.scala 15:7]
  assign O_8_2 = op_O_8_2; // @[MapT.scala 15:7]
  assign O_9_0 = op_O_9_0; // @[MapT.scala 15:7]
  assign O_9_1 = op_O_9_1; // @[MapT.scala 15:7]
  assign O_9_2 = op_O_9_2; // @[MapT.scala 15:7]
  assign O_10_0 = op_O_10_0; // @[MapT.scala 15:7]
  assign O_10_1 = op_O_10_1; // @[MapT.scala 15:7]
  assign O_10_2 = op_O_10_2; // @[MapT.scala 15:7]
  assign O_11_0 = op_O_11_0; // @[MapT.scala 15:7]
  assign O_11_1 = op_O_11_1; // @[MapT.scala 15:7]
  assign O_11_2 = op_O_11_2; // @[MapT.scala 15:7]
  assign O_12_0 = op_O_12_0; // @[MapT.scala 15:7]
  assign O_12_1 = op_O_12_1; // @[MapT.scala 15:7]
  assign O_12_2 = op_O_12_2; // @[MapT.scala 15:7]
  assign O_13_0 = op_O_13_0; // @[MapT.scala 15:7]
  assign O_13_1 = op_O_13_1; // @[MapT.scala 15:7]
  assign O_13_2 = op_O_13_2; // @[MapT.scala 15:7]
  assign O_14_0 = op_O_14_0; // @[MapT.scala 15:7]
  assign O_14_1 = op_O_14_1; // @[MapT.scala 15:7]
  assign O_14_2 = op_O_14_2; // @[MapT.scala 15:7]
  assign O_15_0 = op_O_15_0; // @[MapT.scala 15:7]
  assign O_15_1 = op_O_15_1; // @[MapT.scala 15:7]
  assign O_15_2 = op_O_15_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_2(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_0_2 = I0_2; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
  assign O_1_2 = I1_2; // @[Tuple.scala 13:32]
endmodule
module Map2S_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_2_2,
  input  [7:0] I0_3_0,
  input  [7:0] I0_3_1,
  input  [7:0] I0_3_2,
  input  [7:0] I0_4_0,
  input  [7:0] I0_4_1,
  input  [7:0] I0_4_2,
  input  [7:0] I0_5_0,
  input  [7:0] I0_5_1,
  input  [7:0] I0_5_2,
  input  [7:0] I0_6_0,
  input  [7:0] I0_6_1,
  input  [7:0] I0_6_2,
  input  [7:0] I0_7_0,
  input  [7:0] I0_7_1,
  input  [7:0] I0_7_2,
  input  [7:0] I0_8_0,
  input  [7:0] I0_8_1,
  input  [7:0] I0_8_2,
  input  [7:0] I0_9_0,
  input  [7:0] I0_9_1,
  input  [7:0] I0_9_2,
  input  [7:0] I0_10_0,
  input  [7:0] I0_10_1,
  input  [7:0] I0_10_2,
  input  [7:0] I0_11_0,
  input  [7:0] I0_11_1,
  input  [7:0] I0_11_2,
  input  [7:0] I0_12_0,
  input  [7:0] I0_12_1,
  input  [7:0] I0_12_2,
  input  [7:0] I0_13_0,
  input  [7:0] I0_13_1,
  input  [7:0] I0_13_2,
  input  [7:0] I0_14_0,
  input  [7:0] I0_14_1,
  input  [7:0] I0_14_2,
  input  [7:0] I0_15_0,
  input  [7:0] I0_15_1,
  input  [7:0] I0_15_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  input  [7:0] I1_2_0,
  input  [7:0] I1_2_1,
  input  [7:0] I1_2_2,
  input  [7:0] I1_3_0,
  input  [7:0] I1_3_1,
  input  [7:0] I1_3_2,
  input  [7:0] I1_4_0,
  input  [7:0] I1_4_1,
  input  [7:0] I1_4_2,
  input  [7:0] I1_5_0,
  input  [7:0] I1_5_1,
  input  [7:0] I1_5_2,
  input  [7:0] I1_6_0,
  input  [7:0] I1_6_1,
  input  [7:0] I1_6_2,
  input  [7:0] I1_7_0,
  input  [7:0] I1_7_1,
  input  [7:0] I1_7_2,
  input  [7:0] I1_8_0,
  input  [7:0] I1_8_1,
  input  [7:0] I1_8_2,
  input  [7:0] I1_9_0,
  input  [7:0] I1_9_1,
  input  [7:0] I1_9_2,
  input  [7:0] I1_10_0,
  input  [7:0] I1_10_1,
  input  [7:0] I1_10_2,
  input  [7:0] I1_11_0,
  input  [7:0] I1_11_1,
  input  [7:0] I1_11_2,
  input  [7:0] I1_12_0,
  input  [7:0] I1_12_1,
  input  [7:0] I1_12_2,
  input  [7:0] I1_13_0,
  input  [7:0] I1_13_1,
  input  [7:0] I1_13_2,
  input  [7:0] I1_14_0,
  input  [7:0] I1_14_1,
  input  [7:0] I1_14_2,
  input  [7:0] I1_15_0,
  input  [7:0] I1_15_1,
  input  [7:0] I1_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator_2 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I0_2(other_ops_2_I0_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I0_2(other_ops_3_I0_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I0_2(other_ops_4_I0_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I0_2(other_ops_5_I0_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I0_2(other_ops_6_I0_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I0_2(other_ops_7_I0_2),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .I1_2(other_ops_7_I1_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I0_2(other_ops_8_I0_2),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .I1_2(other_ops_8_I1_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I0_2(other_ops_9_I0_2),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .I1_2(other_ops_9_I1_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I0_2(other_ops_10_I0_2),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .I1_2(other_ops_10_I1_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I0_2(other_ops_11_I0_2),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .I1_2(other_ops_11_I1_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I0_2(other_ops_12_I0_2),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .I1_2(other_ops_12_I1_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I0_2(other_ops_13_I0_2),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .I1_2(other_ops_13_I1_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2)
  );
  SSeqTupleCreator_2 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I0_2(other_ops_14_I0_2),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .I1_2(other_ops_14_I1_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_2 = I0_3_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_2 = I0_4_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_2 = I0_5_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_2 = I0_6_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_2 = I0_7_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_2 = I0_8_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_2 = I1_8_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_2 = I0_9_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_2 = I1_9_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_2 = I0_10_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_2 = I1_10_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_2 = I0_11_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_2 = I1_11_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_2 = I0_12_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_2 = I1_12_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_2 = I0_13_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_2 = I1_13_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_2 = I0_14_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_2 = I1_14_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_2 = I0_15_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_2 = I1_15_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_2_2,
  input  [7:0] I0_3_0,
  input  [7:0] I0_3_1,
  input  [7:0] I0_3_2,
  input  [7:0] I0_4_0,
  input  [7:0] I0_4_1,
  input  [7:0] I0_4_2,
  input  [7:0] I0_5_0,
  input  [7:0] I0_5_1,
  input  [7:0] I0_5_2,
  input  [7:0] I0_6_0,
  input  [7:0] I0_6_1,
  input  [7:0] I0_6_2,
  input  [7:0] I0_7_0,
  input  [7:0] I0_7_1,
  input  [7:0] I0_7_2,
  input  [7:0] I0_8_0,
  input  [7:0] I0_8_1,
  input  [7:0] I0_8_2,
  input  [7:0] I0_9_0,
  input  [7:0] I0_9_1,
  input  [7:0] I0_9_2,
  input  [7:0] I0_10_0,
  input  [7:0] I0_10_1,
  input  [7:0] I0_10_2,
  input  [7:0] I0_11_0,
  input  [7:0] I0_11_1,
  input  [7:0] I0_11_2,
  input  [7:0] I0_12_0,
  input  [7:0] I0_12_1,
  input  [7:0] I0_12_2,
  input  [7:0] I0_13_0,
  input  [7:0] I0_13_1,
  input  [7:0] I0_13_2,
  input  [7:0] I0_14_0,
  input  [7:0] I0_14_1,
  input  [7:0] I0_14_2,
  input  [7:0] I0_15_0,
  input  [7:0] I0_15_1,
  input  [7:0] I0_15_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  input  [7:0] I1_2_0,
  input  [7:0] I1_2_1,
  input  [7:0] I1_2_2,
  input  [7:0] I1_3_0,
  input  [7:0] I1_3_1,
  input  [7:0] I1_3_2,
  input  [7:0] I1_4_0,
  input  [7:0] I1_4_1,
  input  [7:0] I1_4_2,
  input  [7:0] I1_5_0,
  input  [7:0] I1_5_1,
  input  [7:0] I1_5_2,
  input  [7:0] I1_6_0,
  input  [7:0] I1_6_1,
  input  [7:0] I1_6_2,
  input  [7:0] I1_7_0,
  input  [7:0] I1_7_1,
  input  [7:0] I1_7_2,
  input  [7:0] I1_8_0,
  input  [7:0] I1_8_1,
  input  [7:0] I1_8_2,
  input  [7:0] I1_9_0,
  input  [7:0] I1_9_1,
  input  [7:0] I1_9_2,
  input  [7:0] I1_10_0,
  input  [7:0] I1_10_1,
  input  [7:0] I1_10_2,
  input  [7:0] I1_11_0,
  input  [7:0] I1_11_1,
  input  [7:0] I1_11_2,
  input  [7:0] I1_12_0,
  input  [7:0] I1_12_1,
  input  [7:0] I1_12_2,
  input  [7:0] I1_13_0,
  input  [7:0] I1_13_1,
  input  [7:0] I1_13_2,
  input  [7:0] I1_14_0,
  input  [7:0] I1_14_1,
  input  [7:0] I1_14_2,
  input  [7:0] I1_15_0,
  input  [7:0] I1_15_1,
  input  [7:0] I1_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1_2; // @[Map2T.scala 8:20]
  Map2S_4 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_0_2(op_I0_0_2),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_1_2(op_I0_1_2),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_2_2(op_I0_2_2),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_3_2(op_I0_3_2),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_4_2(op_I0_4_2),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_5_2(op_I0_5_2),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_6_2(op_I0_6_2),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_7_2(op_I0_7_2),
    .I0_8_0(op_I0_8_0),
    .I0_8_1(op_I0_8_1),
    .I0_8_2(op_I0_8_2),
    .I0_9_0(op_I0_9_0),
    .I0_9_1(op_I0_9_1),
    .I0_9_2(op_I0_9_2),
    .I0_10_0(op_I0_10_0),
    .I0_10_1(op_I0_10_1),
    .I0_10_2(op_I0_10_2),
    .I0_11_0(op_I0_11_0),
    .I0_11_1(op_I0_11_1),
    .I0_11_2(op_I0_11_2),
    .I0_12_0(op_I0_12_0),
    .I0_12_1(op_I0_12_1),
    .I0_12_2(op_I0_12_2),
    .I0_13_0(op_I0_13_0),
    .I0_13_1(op_I0_13_1),
    .I0_13_2(op_I0_13_2),
    .I0_14_0(op_I0_14_0),
    .I0_14_1(op_I0_14_1),
    .I0_14_2(op_I0_14_2),
    .I0_15_0(op_I0_15_0),
    .I0_15_1(op_I0_15_1),
    .I0_15_2(op_I0_15_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .I1_8_0(op_I1_8_0),
    .I1_8_1(op_I1_8_1),
    .I1_8_2(op_I1_8_2),
    .I1_9_0(op_I1_9_0),
    .I1_9_1(op_I1_9_1),
    .I1_9_2(op_I1_9_2),
    .I1_10_0(op_I1_10_0),
    .I1_10_1(op_I1_10_1),
    .I1_10_2(op_I1_10_2),
    .I1_11_0(op_I1_11_0),
    .I1_11_1(op_I1_11_1),
    .I1_11_2(op_I1_11_2),
    .I1_12_0(op_I1_12_0),
    .I1_12_1(op_I1_12_1),
    .I1_12_2(op_I1_12_2),
    .I1_13_0(op_I1_13_0),
    .I1_13_1(op_I1_13_1),
    .I1_13_2(op_I1_13_2),
    .I1_14_0(op_I1_14_0),
    .I1_14_1(op_I1_14_1),
    .I1_14_2(op_I1_14_2),
    .I1_15_0(op_I1_15_0),
    .I1_15_1(op_I1_15_1),
    .I1_15_2(op_I1_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign O_8_0_0 = op_O_8_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_1 = op_O_8_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_2 = op_O_8_0_2; // @[Map2T.scala 17:7]
  assign O_8_1_0 = op_O_8_1_0; // @[Map2T.scala 17:7]
  assign O_8_1_1 = op_O_8_1_1; // @[Map2T.scala 17:7]
  assign O_8_1_2 = op_O_8_1_2; // @[Map2T.scala 17:7]
  assign O_9_0_0 = op_O_9_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_1 = op_O_9_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_2 = op_O_9_0_2; // @[Map2T.scala 17:7]
  assign O_9_1_0 = op_O_9_1_0; // @[Map2T.scala 17:7]
  assign O_9_1_1 = op_O_9_1_1; // @[Map2T.scala 17:7]
  assign O_9_1_2 = op_O_9_1_2; // @[Map2T.scala 17:7]
  assign O_10_0_0 = op_O_10_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_1 = op_O_10_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_2 = op_O_10_0_2; // @[Map2T.scala 17:7]
  assign O_10_1_0 = op_O_10_1_0; // @[Map2T.scala 17:7]
  assign O_10_1_1 = op_O_10_1_1; // @[Map2T.scala 17:7]
  assign O_10_1_2 = op_O_10_1_2; // @[Map2T.scala 17:7]
  assign O_11_0_0 = op_O_11_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_1 = op_O_11_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_2 = op_O_11_0_2; // @[Map2T.scala 17:7]
  assign O_11_1_0 = op_O_11_1_0; // @[Map2T.scala 17:7]
  assign O_11_1_1 = op_O_11_1_1; // @[Map2T.scala 17:7]
  assign O_11_1_2 = op_O_11_1_2; // @[Map2T.scala 17:7]
  assign O_12_0_0 = op_O_12_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_1 = op_O_12_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_2 = op_O_12_0_2; // @[Map2T.scala 17:7]
  assign O_12_1_0 = op_O_12_1_0; // @[Map2T.scala 17:7]
  assign O_12_1_1 = op_O_12_1_1; // @[Map2T.scala 17:7]
  assign O_12_1_2 = op_O_12_1_2; // @[Map2T.scala 17:7]
  assign O_13_0_0 = op_O_13_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_1 = op_O_13_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_2 = op_O_13_0_2; // @[Map2T.scala 17:7]
  assign O_13_1_0 = op_O_13_1_0; // @[Map2T.scala 17:7]
  assign O_13_1_1 = op_O_13_1_1; // @[Map2T.scala 17:7]
  assign O_13_1_2 = op_O_13_1_2; // @[Map2T.scala 17:7]
  assign O_14_0_0 = op_O_14_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_1 = op_O_14_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_2 = op_O_14_0_2; // @[Map2T.scala 17:7]
  assign O_14_1_0 = op_O_14_1_0; // @[Map2T.scala 17:7]
  assign O_14_1_1 = op_O_14_1_1; // @[Map2T.scala 17:7]
  assign O_14_1_2 = op_O_14_1_2; // @[Map2T.scala 17:7]
  assign O_15_0_0 = op_O_15_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_1 = op_O_15_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_2 = op_O_15_0_2; // @[Map2T.scala 17:7]
  assign O_15_1_0 = op_O_15_1_0; // @[Map2T.scala 17:7]
  assign O_15_1_1 = op_O_15_1_1; // @[Map2T.scala 17:7]
  assign O_15_1_2 = op_O_15_1_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_2 = I0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_2 = I0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_2_2 = I0_2_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_3_2 = I0_3_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_4_2 = I0_4_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_5_2 = I0_5_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_6_2 = I0_6_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_7_2 = I0_7_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0 = I0_8_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1 = I0_8_1; // @[Map2T.scala 15:11]
  assign op_I0_8_2 = I0_8_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0 = I0_9_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1 = I0_9_1; // @[Map2T.scala 15:11]
  assign op_I0_9_2 = I0_9_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0 = I0_10_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1 = I0_10_1; // @[Map2T.scala 15:11]
  assign op_I0_10_2 = I0_10_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0 = I0_11_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1 = I0_11_1; // @[Map2T.scala 15:11]
  assign op_I0_11_2 = I0_11_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0 = I0_12_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1 = I0_12_1; // @[Map2T.scala 15:11]
  assign op_I0_12_2 = I0_12_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0 = I0_13_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1 = I0_13_1; // @[Map2T.scala 15:11]
  assign op_I0_13_2 = I0_13_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0 = I0_14_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1 = I0_14_1; // @[Map2T.scala 15:11]
  assign op_I0_14_2 = I0_14_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0 = I0_15_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1 = I0_15_1; // @[Map2T.scala 15:11]
  assign op_I0_15_2 = I0_15_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
  assign op_I1_8_0 = I1_8_0; // @[Map2T.scala 16:11]
  assign op_I1_8_1 = I1_8_1; // @[Map2T.scala 16:11]
  assign op_I1_8_2 = I1_8_2; // @[Map2T.scala 16:11]
  assign op_I1_9_0 = I1_9_0; // @[Map2T.scala 16:11]
  assign op_I1_9_1 = I1_9_1; // @[Map2T.scala 16:11]
  assign op_I1_9_2 = I1_9_2; // @[Map2T.scala 16:11]
  assign op_I1_10_0 = I1_10_0; // @[Map2T.scala 16:11]
  assign op_I1_10_1 = I1_10_1; // @[Map2T.scala 16:11]
  assign op_I1_10_2 = I1_10_2; // @[Map2T.scala 16:11]
  assign op_I1_11_0 = I1_11_0; // @[Map2T.scala 16:11]
  assign op_I1_11_1 = I1_11_1; // @[Map2T.scala 16:11]
  assign op_I1_11_2 = I1_11_2; // @[Map2T.scala 16:11]
  assign op_I1_12_0 = I1_12_0; // @[Map2T.scala 16:11]
  assign op_I1_12_1 = I1_12_1; // @[Map2T.scala 16:11]
  assign op_I1_12_2 = I1_12_2; // @[Map2T.scala 16:11]
  assign op_I1_13_0 = I1_13_0; // @[Map2T.scala 16:11]
  assign op_I1_13_1 = I1_13_1; // @[Map2T.scala 16:11]
  assign op_I1_13_2 = I1_13_2; // @[Map2T.scala 16:11]
  assign op_I1_14_0 = I1_14_0; // @[Map2T.scala 16:11]
  assign op_I1_14_1 = I1_14_1; // @[Map2T.scala 16:11]
  assign op_I1_14_2 = I1_14_2; // @[Map2T.scala 16:11]
  assign op_I1_15_0 = I1_15_0; // @[Map2T.scala 16:11]
  assign op_I1_15_1 = I1_15_1; // @[Map2T.scala 16:11]
  assign op_I1_15_2 = I1_15_2; // @[Map2T.scala 16:11]
endmodule
module SSeqTupleAppender_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 28:14]
  assign O_0_0 = I0_0_0; // @[Tuple.scala 24:34]
  assign O_0_1 = I0_0_1; // @[Tuple.scala 24:34]
  assign O_0_2 = I0_0_2; // @[Tuple.scala 24:34]
  assign O_1_0 = I0_1_0; // @[Tuple.scala 24:34]
  assign O_1_1 = I0_1_1; // @[Tuple.scala 24:34]
  assign O_1_2 = I0_1_2; // @[Tuple.scala 24:34]
  assign O_2_0 = I1_0; // @[Tuple.scala 26:32]
  assign O_2_1 = I1_1; // @[Tuple.scala 26:32]
  assign O_2_2 = I1_2; // @[Tuple.scala 26:32]
endmodule
module Map2S_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_0_1_0,
  input  [7:0] I0_0_1_1,
  input  [7:0] I0_0_1_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_1_1_0,
  input  [7:0] I0_1_1_1,
  input  [7:0] I0_1_1_2,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_2_0_1,
  input  [7:0] I0_2_0_2,
  input  [7:0] I0_2_1_0,
  input  [7:0] I0_2_1_1,
  input  [7:0] I0_2_1_2,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_3_0_1,
  input  [7:0] I0_3_0_2,
  input  [7:0] I0_3_1_0,
  input  [7:0] I0_3_1_1,
  input  [7:0] I0_3_1_2,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_4_0_1,
  input  [7:0] I0_4_0_2,
  input  [7:0] I0_4_1_0,
  input  [7:0] I0_4_1_1,
  input  [7:0] I0_4_1_2,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_5_0_1,
  input  [7:0] I0_5_0_2,
  input  [7:0] I0_5_1_0,
  input  [7:0] I0_5_1_1,
  input  [7:0] I0_5_1_2,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_6_0_1,
  input  [7:0] I0_6_0_2,
  input  [7:0] I0_6_1_0,
  input  [7:0] I0_6_1_1,
  input  [7:0] I0_6_1_2,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_7_0_1,
  input  [7:0] I0_7_0_2,
  input  [7:0] I0_7_1_0,
  input  [7:0] I0_7_1_1,
  input  [7:0] I0_7_1_2,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_8_0_1,
  input  [7:0] I0_8_0_2,
  input  [7:0] I0_8_1_0,
  input  [7:0] I0_8_1_1,
  input  [7:0] I0_8_1_2,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_9_0_1,
  input  [7:0] I0_9_0_2,
  input  [7:0] I0_9_1_0,
  input  [7:0] I0_9_1_1,
  input  [7:0] I0_9_1_2,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_10_0_1,
  input  [7:0] I0_10_0_2,
  input  [7:0] I0_10_1_0,
  input  [7:0] I0_10_1_1,
  input  [7:0] I0_10_1_2,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_11_0_1,
  input  [7:0] I0_11_0_2,
  input  [7:0] I0_11_1_0,
  input  [7:0] I0_11_1_1,
  input  [7:0] I0_11_1_2,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_12_0_1,
  input  [7:0] I0_12_0_2,
  input  [7:0] I0_12_1_0,
  input  [7:0] I0_12_1_1,
  input  [7:0] I0_12_1_2,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_13_0_1,
  input  [7:0] I0_13_0_2,
  input  [7:0] I0_13_1_0,
  input  [7:0] I0_13_1_1,
  input  [7:0] I0_13_1_2,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_14_0_1,
  input  [7:0] I0_14_0_2,
  input  [7:0] I0_14_1_0,
  input  [7:0] I0_14_1_1,
  input  [7:0] I0_14_1_2,
  input  [7:0] I0_15_0_0,
  input  [7:0] I0_15_0_1,
  input  [7:0] I0_15_0_2,
  input  [7:0] I0_15_1_0,
  input  [7:0] I0_15_1_1,
  input  [7:0] I0_15_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  input  [7:0] I1_2_0,
  input  [7:0] I1_2_1,
  input  [7:0] I1_2_2,
  input  [7:0] I1_3_0,
  input  [7:0] I1_3_1,
  input  [7:0] I1_3_2,
  input  [7:0] I1_4_0,
  input  [7:0] I1_4_1,
  input  [7:0] I1_4_2,
  input  [7:0] I1_5_0,
  input  [7:0] I1_5_1,
  input  [7:0] I1_5_2,
  input  [7:0] I1_6_0,
  input  [7:0] I1_6_1,
  input  [7:0] I1_6_2,
  input  [7:0] I1_7_0,
  input  [7:0] I1_7_1,
  input  [7:0] I1_7_2,
  input  [7:0] I1_8_0,
  input  [7:0] I1_8_1,
  input  [7:0] I1_8_2,
  input  [7:0] I1_9_0,
  input  [7:0] I1_9_1,
  input  [7:0] I1_9_2,
  input  [7:0] I1_10_0,
  input  [7:0] I1_10_1,
  input  [7:0] I1_10_2,
  input  [7:0] I1_11_0,
  input  [7:0] I1_11_1,
  input  [7:0] I1_11_2,
  input  [7:0] I1_12_0,
  input  [7:0] I1_12_1,
  input  [7:0] I1_12_2,
  input  [7:0] I1_13_0,
  input  [7:0] I1_13_1,
  input  [7:0] I1_13_2,
  input  [7:0] I1_14_0,
  input  [7:0] I1_14_1,
  input  [7:0] I1_14_2,
  input  [7:0] I1_15_0,
  input  [7:0] I1_15_1,
  input  [7:0] I1_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_8_2_0,
  output [7:0] O_8_2_1,
  output [7:0] O_8_2_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_9_2_0,
  output [7:0] O_9_2_1,
  output [7:0] O_9_2_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_10_2_0,
  output [7:0] O_10_2_1,
  output [7:0] O_10_2_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_11_2_0,
  output [7:0] O_11_2_1,
  output [7:0] O_11_2_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_12_2_0,
  output [7:0] O_12_2_1,
  output [7:0] O_12_2_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_13_2_0,
  output [7:0] O_13_2_1,
  output [7:0] O_13_2_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_14_2_0,
  output [7:0] O_14_2_1,
  output [7:0] O_14_2_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2,
  output [7:0] O_15_2_0,
  output [7:0] O_15_2_1,
  output [7:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_2_2; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_2_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_2_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_2_2; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleAppender_3 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0_0(fst_op_I0_0_0),
    .I0_0_1(fst_op_I0_0_1),
    .I0_0_2(fst_op_I0_0_2),
    .I0_1_0(fst_op_I0_1_0),
    .I0_1_1(fst_op_I0_1_1),
    .I0_1_2(fst_op_I0_1_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0_0(other_ops_0_I0_0_0),
    .I0_0_1(other_ops_0_I0_0_1),
    .I0_0_2(other_ops_0_I0_0_2),
    .I0_1_0(other_ops_0_I0_1_0),
    .I0_1_1(other_ops_0_I0_1_1),
    .I0_1_2(other_ops_0_I0_1_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0_0(other_ops_1_I0_0_0),
    .I0_0_1(other_ops_1_I0_0_1),
    .I0_0_2(other_ops_1_I0_0_2),
    .I0_1_0(other_ops_1_I0_1_0),
    .I0_1_1(other_ops_1_I0_1_1),
    .I0_1_2(other_ops_1_I0_1_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0_0(other_ops_2_I0_0_0),
    .I0_0_1(other_ops_2_I0_0_1),
    .I0_0_2(other_ops_2_I0_0_2),
    .I0_1_0(other_ops_2_I0_1_0),
    .I0_1_1(other_ops_2_I0_1_1),
    .I0_1_2(other_ops_2_I0_1_2),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .I1_2(other_ops_2_I1_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0_0(other_ops_3_I0_0_0),
    .I0_0_1(other_ops_3_I0_0_1),
    .I0_0_2(other_ops_3_I0_0_2),
    .I0_1_0(other_ops_3_I0_1_0),
    .I0_1_1(other_ops_3_I0_1_1),
    .I0_1_2(other_ops_3_I0_1_2),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .I1_2(other_ops_3_I1_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0_0(other_ops_4_I0_0_0),
    .I0_0_1(other_ops_4_I0_0_1),
    .I0_0_2(other_ops_4_I0_0_2),
    .I0_1_0(other_ops_4_I0_1_0),
    .I0_1_1(other_ops_4_I0_1_1),
    .I0_1_2(other_ops_4_I0_1_2),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .I1_2(other_ops_4_I1_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0_0(other_ops_5_I0_0_0),
    .I0_0_1(other_ops_5_I0_0_1),
    .I0_0_2(other_ops_5_I0_0_2),
    .I0_1_0(other_ops_5_I0_1_0),
    .I0_1_1(other_ops_5_I0_1_1),
    .I0_1_2(other_ops_5_I0_1_2),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .I1_2(other_ops_5_I1_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0_0(other_ops_6_I0_0_0),
    .I0_0_1(other_ops_6_I0_0_1),
    .I0_0_2(other_ops_6_I0_0_2),
    .I0_1_0(other_ops_6_I0_1_0),
    .I0_1_1(other_ops_6_I0_1_1),
    .I0_1_2(other_ops_6_I0_1_2),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .I1_2(other_ops_6_I1_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0_0(other_ops_7_I0_0_0),
    .I0_0_1(other_ops_7_I0_0_1),
    .I0_0_2(other_ops_7_I0_0_2),
    .I0_1_0(other_ops_7_I0_1_0),
    .I0_1_1(other_ops_7_I0_1_1),
    .I0_1_2(other_ops_7_I0_1_2),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .I1_2(other_ops_7_I1_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0_0(other_ops_8_I0_0_0),
    .I0_0_1(other_ops_8_I0_0_1),
    .I0_0_2(other_ops_8_I0_0_2),
    .I0_1_0(other_ops_8_I0_1_0),
    .I0_1_1(other_ops_8_I0_1_1),
    .I0_1_2(other_ops_8_I0_1_2),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .I1_2(other_ops_8_I1_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0_0(other_ops_9_I0_0_0),
    .I0_0_1(other_ops_9_I0_0_1),
    .I0_0_2(other_ops_9_I0_0_2),
    .I0_1_0(other_ops_9_I0_1_0),
    .I0_1_1(other_ops_9_I0_1_1),
    .I0_1_2(other_ops_9_I0_1_2),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .I1_2(other_ops_9_I1_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0_0(other_ops_10_I0_0_0),
    .I0_0_1(other_ops_10_I0_0_1),
    .I0_0_2(other_ops_10_I0_0_2),
    .I0_1_0(other_ops_10_I0_1_0),
    .I0_1_1(other_ops_10_I0_1_1),
    .I0_1_2(other_ops_10_I0_1_2),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .I1_2(other_ops_10_I1_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0_0(other_ops_11_I0_0_0),
    .I0_0_1(other_ops_11_I0_0_1),
    .I0_0_2(other_ops_11_I0_0_2),
    .I0_1_0(other_ops_11_I0_1_0),
    .I0_1_1(other_ops_11_I0_1_1),
    .I0_1_2(other_ops_11_I0_1_2),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .I1_2(other_ops_11_I1_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0_0(other_ops_12_I0_0_0),
    .I0_0_1(other_ops_12_I0_0_1),
    .I0_0_2(other_ops_12_I0_0_2),
    .I0_1_0(other_ops_12_I0_1_0),
    .I0_1_1(other_ops_12_I0_1_1),
    .I0_1_2(other_ops_12_I0_1_2),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .I1_2(other_ops_12_I1_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0_0(other_ops_13_I0_0_0),
    .I0_0_1(other_ops_13_I0_0_1),
    .I0_0_2(other_ops_13_I0_0_2),
    .I0_1_0(other_ops_13_I0_1_0),
    .I0_1_1(other_ops_13_I0_1_1),
    .I0_1_2(other_ops_13_I0_1_2),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .I1_2(other_ops_13_I1_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  SSeqTupleAppender_3 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0_0(other_ops_14_I0_0_0),
    .I0_0_1(other_ops_14_I0_0_1),
    .I0_0_2(other_ops_14_I0_0_2),
    .I0_1_0(other_ops_14_I0_1_0),
    .I0_1_1(other_ops_14_I0_1_1),
    .I0_1_2(other_ops_14_I0_1_2),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .I1_2(other_ops_14_I1_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[Map2S.scala 19:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[Map2S.scala 19:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[Map2S.scala 19:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[Map2S.scala 24:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[Map2S.scala 24:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[Map2S.scala 24:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[Map2S.scala 24:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[Map2S.scala 24:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[Map2S.scala 24:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[Map2S.scala 24:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[Map2S.scala 24:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[Map2S.scala 24:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[Map2S.scala 24:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[Map2S.scala 24:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[Map2S.scala 24:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[Map2S.scala 24:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[Map2S.scala 24:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[Map2S.scala 24:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[Map2S.scala 24:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[Map2S.scala 24:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[Map2S.scala 24:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[Map2S.scala 24:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[Map2S.scala 24:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[Map2S.scala 24:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[Map2S.scala 24:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[Map2S.scala 24:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[Map2S.scala 24:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[Map2S.scala 24:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[Map2S.scala 24:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[Map2S.scala 24:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[Map2S.scala 24:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[Map2S.scala 24:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[Map2S.scala 24:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[Map2S.scala 24:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[Map2S.scala 24:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[Map2S.scala 24:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[Map2S.scala 24:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[Map2S.scala 24:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[Map2S.scala 24:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[Map2S.scala 24:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[Map2S.scala 24:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[Map2S.scala 24:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[Map2S.scala 24:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[Map2S.scala 24:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[Map2S.scala 24:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[Map2S.scala 24:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[Map2S.scala 24:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[Map2S.scala 24:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0_0 = I0_0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_1 = I0_0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_0_2 = I0_0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_0 = I0_0_1_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_1 = I0_0_1_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_1_2 = I0_0_1_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = I1_0_2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0_0 = I0_1_0_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_1 = I0_1_0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_0_2 = I0_1_0_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_0 = I0_1_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_1 = I0_1_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1_2 = I0_1_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = I1_1_2; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0_0 = I0_2_0_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_1 = I0_2_0_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_0_2 = I0_2_0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_0 = I0_2_1_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_1 = I0_2_1_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1_2 = I0_2_1_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = I1_2_2; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0_0 = I0_3_0_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_1 = I0_3_0_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_0_2 = I0_3_0_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_0 = I0_3_1_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_1 = I0_3_1_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1_2 = I0_3_1_2; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_2 = I1_3_2; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0_0 = I0_4_0_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_1 = I0_4_0_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_0_2 = I0_4_0_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_0 = I0_4_1_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_1 = I0_4_1_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1_2 = I0_4_1_2; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_2 = I1_4_2; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0_0 = I0_5_0_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_1 = I0_5_0_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_0_2 = I0_5_0_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_0 = I0_5_1_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_1 = I0_5_1_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1_2 = I0_5_1_2; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_2 = I1_5_2; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0_0 = I0_6_0_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_1 = I0_6_0_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_0_2 = I0_6_0_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_0 = I0_6_1_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_1 = I0_6_1_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1_2 = I0_6_1_2; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_2 = I1_6_2; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0_0 = I0_7_0_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_1 = I0_7_0_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_0_2 = I0_7_0_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_0 = I0_7_1_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_1 = I0_7_1_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1_2 = I0_7_1_2; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_2 = I1_7_2; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0_0 = I0_8_0_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_1 = I0_8_0_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_0_2 = I0_8_0_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_0 = I0_8_1_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_1 = I0_8_1_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1_2 = I0_8_1_2; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_2 = I1_8_2; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0_0 = I0_9_0_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_1 = I0_9_0_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_0_2 = I0_9_0_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_0 = I0_9_1_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_1 = I0_9_1_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1_2 = I0_9_1_2; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_2 = I1_9_2; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0_0 = I0_10_0_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_1 = I0_10_0_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_0_2 = I0_10_0_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_0 = I0_10_1_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_1 = I0_10_1_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1_2 = I0_10_1_2; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_2 = I1_10_2; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0_0 = I0_11_0_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_1 = I0_11_0_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_0_2 = I0_11_0_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_0 = I0_11_1_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_1 = I0_11_1_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1_2 = I0_11_1_2; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_2 = I1_11_2; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0_0 = I0_12_0_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_1 = I0_12_0_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_0_2 = I0_12_0_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_0 = I0_12_1_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_1 = I0_12_1_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1_2 = I0_12_1_2; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_2 = I1_12_2; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0_0 = I0_13_0_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_1 = I0_13_0_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_0_2 = I0_13_0_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_0 = I0_13_1_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_1 = I0_13_1_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1_2 = I0_13_1_2; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_2 = I1_13_2; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0_0 = I0_14_0_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_1 = I0_14_0_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_0_2 = I0_14_0_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_0 = I0_14_1_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_1 = I0_14_1_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1_2 = I0_14_1_2; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_2 = I1_14_2; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0_0 = I0_15_0_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_1 = I0_15_0_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_0_2 = I0_15_0_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_0 = I0_15_1_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_1 = I0_15_1_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1_2 = I0_15_1_2; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_2 = I1_15_2; // @[Map2S.scala 23:43]
endmodule
module Map2T_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0_0,
  input  [7:0] I0_0_0_1,
  input  [7:0] I0_0_0_2,
  input  [7:0] I0_0_1_0,
  input  [7:0] I0_0_1_1,
  input  [7:0] I0_0_1_2,
  input  [7:0] I0_1_0_0,
  input  [7:0] I0_1_0_1,
  input  [7:0] I0_1_0_2,
  input  [7:0] I0_1_1_0,
  input  [7:0] I0_1_1_1,
  input  [7:0] I0_1_1_2,
  input  [7:0] I0_2_0_0,
  input  [7:0] I0_2_0_1,
  input  [7:0] I0_2_0_2,
  input  [7:0] I0_2_1_0,
  input  [7:0] I0_2_1_1,
  input  [7:0] I0_2_1_2,
  input  [7:0] I0_3_0_0,
  input  [7:0] I0_3_0_1,
  input  [7:0] I0_3_0_2,
  input  [7:0] I0_3_1_0,
  input  [7:0] I0_3_1_1,
  input  [7:0] I0_3_1_2,
  input  [7:0] I0_4_0_0,
  input  [7:0] I0_4_0_1,
  input  [7:0] I0_4_0_2,
  input  [7:0] I0_4_1_0,
  input  [7:0] I0_4_1_1,
  input  [7:0] I0_4_1_2,
  input  [7:0] I0_5_0_0,
  input  [7:0] I0_5_0_1,
  input  [7:0] I0_5_0_2,
  input  [7:0] I0_5_1_0,
  input  [7:0] I0_5_1_1,
  input  [7:0] I0_5_1_2,
  input  [7:0] I0_6_0_0,
  input  [7:0] I0_6_0_1,
  input  [7:0] I0_6_0_2,
  input  [7:0] I0_6_1_0,
  input  [7:0] I0_6_1_1,
  input  [7:0] I0_6_1_2,
  input  [7:0] I0_7_0_0,
  input  [7:0] I0_7_0_1,
  input  [7:0] I0_7_0_2,
  input  [7:0] I0_7_1_0,
  input  [7:0] I0_7_1_1,
  input  [7:0] I0_7_1_2,
  input  [7:0] I0_8_0_0,
  input  [7:0] I0_8_0_1,
  input  [7:0] I0_8_0_2,
  input  [7:0] I0_8_1_0,
  input  [7:0] I0_8_1_1,
  input  [7:0] I0_8_1_2,
  input  [7:0] I0_9_0_0,
  input  [7:0] I0_9_0_1,
  input  [7:0] I0_9_0_2,
  input  [7:0] I0_9_1_0,
  input  [7:0] I0_9_1_1,
  input  [7:0] I0_9_1_2,
  input  [7:0] I0_10_0_0,
  input  [7:0] I0_10_0_1,
  input  [7:0] I0_10_0_2,
  input  [7:0] I0_10_1_0,
  input  [7:0] I0_10_1_1,
  input  [7:0] I0_10_1_2,
  input  [7:0] I0_11_0_0,
  input  [7:0] I0_11_0_1,
  input  [7:0] I0_11_0_2,
  input  [7:0] I0_11_1_0,
  input  [7:0] I0_11_1_1,
  input  [7:0] I0_11_1_2,
  input  [7:0] I0_12_0_0,
  input  [7:0] I0_12_0_1,
  input  [7:0] I0_12_0_2,
  input  [7:0] I0_12_1_0,
  input  [7:0] I0_12_1_1,
  input  [7:0] I0_12_1_2,
  input  [7:0] I0_13_0_0,
  input  [7:0] I0_13_0_1,
  input  [7:0] I0_13_0_2,
  input  [7:0] I0_13_1_0,
  input  [7:0] I0_13_1_1,
  input  [7:0] I0_13_1_2,
  input  [7:0] I0_14_0_0,
  input  [7:0] I0_14_0_1,
  input  [7:0] I0_14_0_2,
  input  [7:0] I0_14_1_0,
  input  [7:0] I0_14_1_1,
  input  [7:0] I0_14_1_2,
  input  [7:0] I0_15_0_0,
  input  [7:0] I0_15_0_1,
  input  [7:0] I0_15_0_2,
  input  [7:0] I0_15_1_0,
  input  [7:0] I0_15_1_1,
  input  [7:0] I0_15_1_2,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_0_2,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_1_2,
  input  [7:0] I1_2_0,
  input  [7:0] I1_2_1,
  input  [7:0] I1_2_2,
  input  [7:0] I1_3_0,
  input  [7:0] I1_3_1,
  input  [7:0] I1_3_2,
  input  [7:0] I1_4_0,
  input  [7:0] I1_4_1,
  input  [7:0] I1_4_2,
  input  [7:0] I1_5_0,
  input  [7:0] I1_5_1,
  input  [7:0] I1_5_2,
  input  [7:0] I1_6_0,
  input  [7:0] I1_6_1,
  input  [7:0] I1_6_2,
  input  [7:0] I1_7_0,
  input  [7:0] I1_7_1,
  input  [7:0] I1_7_2,
  input  [7:0] I1_8_0,
  input  [7:0] I1_8_1,
  input  [7:0] I1_8_2,
  input  [7:0] I1_9_0,
  input  [7:0] I1_9_1,
  input  [7:0] I1_9_2,
  input  [7:0] I1_10_0,
  input  [7:0] I1_10_1,
  input  [7:0] I1_10_2,
  input  [7:0] I1_11_0,
  input  [7:0] I1_11_1,
  input  [7:0] I1_11_2,
  input  [7:0] I1_12_0,
  input  [7:0] I1_12_1,
  input  [7:0] I1_12_2,
  input  [7:0] I1_13_0,
  input  [7:0] I1_13_1,
  input  [7:0] I1_13_2,
  input  [7:0] I1_14_0,
  input  [7:0] I1_14_1,
  input  [7:0] I1_14_2,
  input  [7:0] I1_15_0,
  input  [7:0] I1_15_1,
  input  [7:0] I1_15_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_8_2_0,
  output [7:0] O_8_2_1,
  output [7:0] O_8_2_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_9_2_0,
  output [7:0] O_9_2_1,
  output [7:0] O_9_2_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_10_2_0,
  output [7:0] O_10_2_1,
  output [7:0] O_10_2_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_11_2_0,
  output [7:0] O_11_2_1,
  output [7:0] O_11_2_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_12_2_0,
  output [7:0] O_12_2_1,
  output [7:0] O_12_2_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_13_2_0,
  output [7:0] O_13_2_1,
  output [7:0] O_13_2_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_14_2_0,
  output [7:0] O_14_2_1,
  output [7:0] O_14_2_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2,
  output [7:0] O_15_2_0,
  output [7:0] O_15_2_1,
  output [7:0] O_15_2_2
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_2; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_2_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1_2; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_2_2; // @[Map2T.scala 8:20]
  Map2S_7 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0_0(op_I0_0_0_0),
    .I0_0_0_1(op_I0_0_0_1),
    .I0_0_0_2(op_I0_0_0_2),
    .I0_0_1_0(op_I0_0_1_0),
    .I0_0_1_1(op_I0_0_1_1),
    .I0_0_1_2(op_I0_0_1_2),
    .I0_1_0_0(op_I0_1_0_0),
    .I0_1_0_1(op_I0_1_0_1),
    .I0_1_0_2(op_I0_1_0_2),
    .I0_1_1_0(op_I0_1_1_0),
    .I0_1_1_1(op_I0_1_1_1),
    .I0_1_1_2(op_I0_1_1_2),
    .I0_2_0_0(op_I0_2_0_0),
    .I0_2_0_1(op_I0_2_0_1),
    .I0_2_0_2(op_I0_2_0_2),
    .I0_2_1_0(op_I0_2_1_0),
    .I0_2_1_1(op_I0_2_1_1),
    .I0_2_1_2(op_I0_2_1_2),
    .I0_3_0_0(op_I0_3_0_0),
    .I0_3_0_1(op_I0_3_0_1),
    .I0_3_0_2(op_I0_3_0_2),
    .I0_3_1_0(op_I0_3_1_0),
    .I0_3_1_1(op_I0_3_1_1),
    .I0_3_1_2(op_I0_3_1_2),
    .I0_4_0_0(op_I0_4_0_0),
    .I0_4_0_1(op_I0_4_0_1),
    .I0_4_0_2(op_I0_4_0_2),
    .I0_4_1_0(op_I0_4_1_0),
    .I0_4_1_1(op_I0_4_1_1),
    .I0_4_1_2(op_I0_4_1_2),
    .I0_5_0_0(op_I0_5_0_0),
    .I0_5_0_1(op_I0_5_0_1),
    .I0_5_0_2(op_I0_5_0_2),
    .I0_5_1_0(op_I0_5_1_0),
    .I0_5_1_1(op_I0_5_1_1),
    .I0_5_1_2(op_I0_5_1_2),
    .I0_6_0_0(op_I0_6_0_0),
    .I0_6_0_1(op_I0_6_0_1),
    .I0_6_0_2(op_I0_6_0_2),
    .I0_6_1_0(op_I0_6_1_0),
    .I0_6_1_1(op_I0_6_1_1),
    .I0_6_1_2(op_I0_6_1_2),
    .I0_7_0_0(op_I0_7_0_0),
    .I0_7_0_1(op_I0_7_0_1),
    .I0_7_0_2(op_I0_7_0_2),
    .I0_7_1_0(op_I0_7_1_0),
    .I0_7_1_1(op_I0_7_1_1),
    .I0_7_1_2(op_I0_7_1_2),
    .I0_8_0_0(op_I0_8_0_0),
    .I0_8_0_1(op_I0_8_0_1),
    .I0_8_0_2(op_I0_8_0_2),
    .I0_8_1_0(op_I0_8_1_0),
    .I0_8_1_1(op_I0_8_1_1),
    .I0_8_1_2(op_I0_8_1_2),
    .I0_9_0_0(op_I0_9_0_0),
    .I0_9_0_1(op_I0_9_0_1),
    .I0_9_0_2(op_I0_9_0_2),
    .I0_9_1_0(op_I0_9_1_0),
    .I0_9_1_1(op_I0_9_1_1),
    .I0_9_1_2(op_I0_9_1_2),
    .I0_10_0_0(op_I0_10_0_0),
    .I0_10_0_1(op_I0_10_0_1),
    .I0_10_0_2(op_I0_10_0_2),
    .I0_10_1_0(op_I0_10_1_0),
    .I0_10_1_1(op_I0_10_1_1),
    .I0_10_1_2(op_I0_10_1_2),
    .I0_11_0_0(op_I0_11_0_0),
    .I0_11_0_1(op_I0_11_0_1),
    .I0_11_0_2(op_I0_11_0_2),
    .I0_11_1_0(op_I0_11_1_0),
    .I0_11_1_1(op_I0_11_1_1),
    .I0_11_1_2(op_I0_11_1_2),
    .I0_12_0_0(op_I0_12_0_0),
    .I0_12_0_1(op_I0_12_0_1),
    .I0_12_0_2(op_I0_12_0_2),
    .I0_12_1_0(op_I0_12_1_0),
    .I0_12_1_1(op_I0_12_1_1),
    .I0_12_1_2(op_I0_12_1_2),
    .I0_13_0_0(op_I0_13_0_0),
    .I0_13_0_1(op_I0_13_0_1),
    .I0_13_0_2(op_I0_13_0_2),
    .I0_13_1_0(op_I0_13_1_0),
    .I0_13_1_1(op_I0_13_1_1),
    .I0_13_1_2(op_I0_13_1_2),
    .I0_14_0_0(op_I0_14_0_0),
    .I0_14_0_1(op_I0_14_0_1),
    .I0_14_0_2(op_I0_14_0_2),
    .I0_14_1_0(op_I0_14_1_0),
    .I0_14_1_1(op_I0_14_1_1),
    .I0_14_1_2(op_I0_14_1_2),
    .I0_15_0_0(op_I0_15_0_0),
    .I0_15_0_1(op_I0_15_0_1),
    .I0_15_0_2(op_I0_15_0_2),
    .I0_15_1_0(op_I0_15_1_0),
    .I0_15_1_1(op_I0_15_1_1),
    .I0_15_1_2(op_I0_15_1_2),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_0_2(op_I1_0_2),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_1_2(op_I1_1_2),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_2_2(op_I1_2_2),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_3_2(op_I1_3_2),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_4_2(op_I1_4_2),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_5_2(op_I1_5_2),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_6_2(op_I1_6_2),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_7_2(op_I1_7_2),
    .I1_8_0(op_I1_8_0),
    .I1_8_1(op_I1_8_1),
    .I1_8_2(op_I1_8_2),
    .I1_9_0(op_I1_9_0),
    .I1_9_1(op_I1_9_1),
    .I1_9_2(op_I1_9_2),
    .I1_10_0(op_I1_10_0),
    .I1_10_1(op_I1_10_1),
    .I1_10_2(op_I1_10_2),
    .I1_11_0(op_I1_11_0),
    .I1_11_1(op_I1_11_1),
    .I1_11_2(op_I1_11_2),
    .I1_12_0(op_I1_12_0),
    .I1_12_1(op_I1_12_1),
    .I1_12_2(op_I1_12_2),
    .I1_13_0(op_I1_13_0),
    .I1_13_1(op_I1_13_1),
    .I1_13_2(op_I1_13_2),
    .I1_14_0(op_I1_14_0),
    .I1_14_1(op_I1_14_1),
    .I1_14_2(op_I1_14_2),
    .I1_15_0(op_I1_15_0),
    .I1_15_1(op_I1_15_1),
    .I1_15_2(op_I1_15_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_8_2_0(op_O_8_2_0),
    .O_8_2_1(op_O_8_2_1),
    .O_8_2_2(op_O_8_2_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_9_2_0(op_O_9_2_0),
    .O_9_2_1(op_O_9_2_1),
    .O_9_2_2(op_O_9_2_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_10_2_0(op_O_10_2_0),
    .O_10_2_1(op_O_10_2_1),
    .O_10_2_2(op_O_10_2_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_11_2_0(op_O_11_2_0),
    .O_11_2_1(op_O_11_2_1),
    .O_11_2_2(op_O_11_2_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_12_2_0(op_O_12_2_0),
    .O_12_2_1(op_O_12_2_1),
    .O_12_2_2(op_O_12_2_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_13_2_0(op_O_13_2_0),
    .O_13_2_1(op_O_13_2_1),
    .O_13_2_2(op_O_13_2_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_14_2_0(op_O_14_2_0),
    .O_14_2_1(op_O_14_2_1),
    .O_14_2_2(op_O_14_2_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2),
    .O_15_2_0(op_O_15_2_0),
    .O_15_2_1(op_O_15_2_1),
    .O_15_2_2(op_O_15_2_2)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_0_2 = op_O_0_0_2; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_0_1_2 = op_O_0_1_2; // @[Map2T.scala 17:7]
  assign O_0_2_0 = op_O_0_2_0; // @[Map2T.scala 17:7]
  assign O_0_2_1 = op_O_0_2_1; // @[Map2T.scala 17:7]
  assign O_0_2_2 = op_O_0_2_2; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_0_2 = op_O_1_0_2; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_1_1_2 = op_O_1_1_2; // @[Map2T.scala 17:7]
  assign O_1_2_0 = op_O_1_2_0; // @[Map2T.scala 17:7]
  assign O_1_2_1 = op_O_1_2_1; // @[Map2T.scala 17:7]
  assign O_1_2_2 = op_O_1_2_2; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_0_2 = op_O_2_0_2; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_2_1_2 = op_O_2_1_2; // @[Map2T.scala 17:7]
  assign O_2_2_0 = op_O_2_2_0; // @[Map2T.scala 17:7]
  assign O_2_2_1 = op_O_2_2_1; // @[Map2T.scala 17:7]
  assign O_2_2_2 = op_O_2_2_2; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_0_2 = op_O_3_0_2; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_3_1_2 = op_O_3_1_2; // @[Map2T.scala 17:7]
  assign O_3_2_0 = op_O_3_2_0; // @[Map2T.scala 17:7]
  assign O_3_2_1 = op_O_3_2_1; // @[Map2T.scala 17:7]
  assign O_3_2_2 = op_O_3_2_2; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_0_2 = op_O_4_0_2; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_4_1_2 = op_O_4_1_2; // @[Map2T.scala 17:7]
  assign O_4_2_0 = op_O_4_2_0; // @[Map2T.scala 17:7]
  assign O_4_2_1 = op_O_4_2_1; // @[Map2T.scala 17:7]
  assign O_4_2_2 = op_O_4_2_2; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_0_2 = op_O_5_0_2; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_5_1_2 = op_O_5_1_2; // @[Map2T.scala 17:7]
  assign O_5_2_0 = op_O_5_2_0; // @[Map2T.scala 17:7]
  assign O_5_2_1 = op_O_5_2_1; // @[Map2T.scala 17:7]
  assign O_5_2_2 = op_O_5_2_2; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_0_2 = op_O_6_0_2; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_6_1_2 = op_O_6_1_2; // @[Map2T.scala 17:7]
  assign O_6_2_0 = op_O_6_2_0; // @[Map2T.scala 17:7]
  assign O_6_2_1 = op_O_6_2_1; // @[Map2T.scala 17:7]
  assign O_6_2_2 = op_O_6_2_2; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_0_2 = op_O_7_0_2; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_7_1_2 = op_O_7_1_2; // @[Map2T.scala 17:7]
  assign O_7_2_0 = op_O_7_2_0; // @[Map2T.scala 17:7]
  assign O_7_2_1 = op_O_7_2_1; // @[Map2T.scala 17:7]
  assign O_7_2_2 = op_O_7_2_2; // @[Map2T.scala 17:7]
  assign O_8_0_0 = op_O_8_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_1 = op_O_8_0_1; // @[Map2T.scala 17:7]
  assign O_8_0_2 = op_O_8_0_2; // @[Map2T.scala 17:7]
  assign O_8_1_0 = op_O_8_1_0; // @[Map2T.scala 17:7]
  assign O_8_1_1 = op_O_8_1_1; // @[Map2T.scala 17:7]
  assign O_8_1_2 = op_O_8_1_2; // @[Map2T.scala 17:7]
  assign O_8_2_0 = op_O_8_2_0; // @[Map2T.scala 17:7]
  assign O_8_2_1 = op_O_8_2_1; // @[Map2T.scala 17:7]
  assign O_8_2_2 = op_O_8_2_2; // @[Map2T.scala 17:7]
  assign O_9_0_0 = op_O_9_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_1 = op_O_9_0_1; // @[Map2T.scala 17:7]
  assign O_9_0_2 = op_O_9_0_2; // @[Map2T.scala 17:7]
  assign O_9_1_0 = op_O_9_1_0; // @[Map2T.scala 17:7]
  assign O_9_1_1 = op_O_9_1_1; // @[Map2T.scala 17:7]
  assign O_9_1_2 = op_O_9_1_2; // @[Map2T.scala 17:7]
  assign O_9_2_0 = op_O_9_2_0; // @[Map2T.scala 17:7]
  assign O_9_2_1 = op_O_9_2_1; // @[Map2T.scala 17:7]
  assign O_9_2_2 = op_O_9_2_2; // @[Map2T.scala 17:7]
  assign O_10_0_0 = op_O_10_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_1 = op_O_10_0_1; // @[Map2T.scala 17:7]
  assign O_10_0_2 = op_O_10_0_2; // @[Map2T.scala 17:7]
  assign O_10_1_0 = op_O_10_1_0; // @[Map2T.scala 17:7]
  assign O_10_1_1 = op_O_10_1_1; // @[Map2T.scala 17:7]
  assign O_10_1_2 = op_O_10_1_2; // @[Map2T.scala 17:7]
  assign O_10_2_0 = op_O_10_2_0; // @[Map2T.scala 17:7]
  assign O_10_2_1 = op_O_10_2_1; // @[Map2T.scala 17:7]
  assign O_10_2_2 = op_O_10_2_2; // @[Map2T.scala 17:7]
  assign O_11_0_0 = op_O_11_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_1 = op_O_11_0_1; // @[Map2T.scala 17:7]
  assign O_11_0_2 = op_O_11_0_2; // @[Map2T.scala 17:7]
  assign O_11_1_0 = op_O_11_1_0; // @[Map2T.scala 17:7]
  assign O_11_1_1 = op_O_11_1_1; // @[Map2T.scala 17:7]
  assign O_11_1_2 = op_O_11_1_2; // @[Map2T.scala 17:7]
  assign O_11_2_0 = op_O_11_2_0; // @[Map2T.scala 17:7]
  assign O_11_2_1 = op_O_11_2_1; // @[Map2T.scala 17:7]
  assign O_11_2_2 = op_O_11_2_2; // @[Map2T.scala 17:7]
  assign O_12_0_0 = op_O_12_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_1 = op_O_12_0_1; // @[Map2T.scala 17:7]
  assign O_12_0_2 = op_O_12_0_2; // @[Map2T.scala 17:7]
  assign O_12_1_0 = op_O_12_1_0; // @[Map2T.scala 17:7]
  assign O_12_1_1 = op_O_12_1_1; // @[Map2T.scala 17:7]
  assign O_12_1_2 = op_O_12_1_2; // @[Map2T.scala 17:7]
  assign O_12_2_0 = op_O_12_2_0; // @[Map2T.scala 17:7]
  assign O_12_2_1 = op_O_12_2_1; // @[Map2T.scala 17:7]
  assign O_12_2_2 = op_O_12_2_2; // @[Map2T.scala 17:7]
  assign O_13_0_0 = op_O_13_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_1 = op_O_13_0_1; // @[Map2T.scala 17:7]
  assign O_13_0_2 = op_O_13_0_2; // @[Map2T.scala 17:7]
  assign O_13_1_0 = op_O_13_1_0; // @[Map2T.scala 17:7]
  assign O_13_1_1 = op_O_13_1_1; // @[Map2T.scala 17:7]
  assign O_13_1_2 = op_O_13_1_2; // @[Map2T.scala 17:7]
  assign O_13_2_0 = op_O_13_2_0; // @[Map2T.scala 17:7]
  assign O_13_2_1 = op_O_13_2_1; // @[Map2T.scala 17:7]
  assign O_13_2_2 = op_O_13_2_2; // @[Map2T.scala 17:7]
  assign O_14_0_0 = op_O_14_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_1 = op_O_14_0_1; // @[Map2T.scala 17:7]
  assign O_14_0_2 = op_O_14_0_2; // @[Map2T.scala 17:7]
  assign O_14_1_0 = op_O_14_1_0; // @[Map2T.scala 17:7]
  assign O_14_1_1 = op_O_14_1_1; // @[Map2T.scala 17:7]
  assign O_14_1_2 = op_O_14_1_2; // @[Map2T.scala 17:7]
  assign O_14_2_0 = op_O_14_2_0; // @[Map2T.scala 17:7]
  assign O_14_2_1 = op_O_14_2_1; // @[Map2T.scala 17:7]
  assign O_14_2_2 = op_O_14_2_2; // @[Map2T.scala 17:7]
  assign O_15_0_0 = op_O_15_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_1 = op_O_15_0_1; // @[Map2T.scala 17:7]
  assign O_15_0_2 = op_O_15_0_2; // @[Map2T.scala 17:7]
  assign O_15_1_0 = op_O_15_1_0; // @[Map2T.scala 17:7]
  assign O_15_1_1 = op_O_15_1_1; // @[Map2T.scala 17:7]
  assign O_15_1_2 = op_O_15_1_2; // @[Map2T.scala 17:7]
  assign O_15_2_0 = op_O_15_2_0; // @[Map2T.scala 17:7]
  assign O_15_2_1 = op_O_15_2_1; // @[Map2T.scala 17:7]
  assign O_15_2_2 = op_O_15_2_2; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0_0 = I0_0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_0_1 = I0_0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_0_0_2 = I0_0_0_2; // @[Map2T.scala 15:11]
  assign op_I0_0_1_0 = I0_0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1_1 = I0_0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_0_1_2 = I0_0_1_2; // @[Map2T.scala 15:11]
  assign op_I0_1_0_0 = I0_1_0_0; // @[Map2T.scala 15:11]
  assign op_I0_1_0_1 = I0_1_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0_2 = I0_1_0_2; // @[Map2T.scala 15:11]
  assign op_I0_1_1_0 = I0_1_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1_1 = I0_1_1_1; // @[Map2T.scala 15:11]
  assign op_I0_1_1_2 = I0_1_1_2; // @[Map2T.scala 15:11]
  assign op_I0_2_0_0 = I0_2_0_0; // @[Map2T.scala 15:11]
  assign op_I0_2_0_1 = I0_2_0_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0_2 = I0_2_0_2; // @[Map2T.scala 15:11]
  assign op_I0_2_1_0 = I0_2_1_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1_1 = I0_2_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_1_2 = I0_2_1_2; // @[Map2T.scala 15:11]
  assign op_I0_3_0_0 = I0_3_0_0; // @[Map2T.scala 15:11]
  assign op_I0_3_0_1 = I0_3_0_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0_2 = I0_3_0_2; // @[Map2T.scala 15:11]
  assign op_I0_3_1_0 = I0_3_1_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1_1 = I0_3_1_1; // @[Map2T.scala 15:11]
  assign op_I0_3_1_2 = I0_3_1_2; // @[Map2T.scala 15:11]
  assign op_I0_4_0_0 = I0_4_0_0; // @[Map2T.scala 15:11]
  assign op_I0_4_0_1 = I0_4_0_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0_2 = I0_4_0_2; // @[Map2T.scala 15:11]
  assign op_I0_4_1_0 = I0_4_1_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1_1 = I0_4_1_1; // @[Map2T.scala 15:11]
  assign op_I0_4_1_2 = I0_4_1_2; // @[Map2T.scala 15:11]
  assign op_I0_5_0_0 = I0_5_0_0; // @[Map2T.scala 15:11]
  assign op_I0_5_0_1 = I0_5_0_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0_2 = I0_5_0_2; // @[Map2T.scala 15:11]
  assign op_I0_5_1_0 = I0_5_1_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1_1 = I0_5_1_1; // @[Map2T.scala 15:11]
  assign op_I0_5_1_2 = I0_5_1_2; // @[Map2T.scala 15:11]
  assign op_I0_6_0_0 = I0_6_0_0; // @[Map2T.scala 15:11]
  assign op_I0_6_0_1 = I0_6_0_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0_2 = I0_6_0_2; // @[Map2T.scala 15:11]
  assign op_I0_6_1_0 = I0_6_1_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1_1 = I0_6_1_1; // @[Map2T.scala 15:11]
  assign op_I0_6_1_2 = I0_6_1_2; // @[Map2T.scala 15:11]
  assign op_I0_7_0_0 = I0_7_0_0; // @[Map2T.scala 15:11]
  assign op_I0_7_0_1 = I0_7_0_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0_2 = I0_7_0_2; // @[Map2T.scala 15:11]
  assign op_I0_7_1_0 = I0_7_1_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1_1 = I0_7_1_1; // @[Map2T.scala 15:11]
  assign op_I0_7_1_2 = I0_7_1_2; // @[Map2T.scala 15:11]
  assign op_I0_8_0_0 = I0_8_0_0; // @[Map2T.scala 15:11]
  assign op_I0_8_0_1 = I0_8_0_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0_2 = I0_8_0_2; // @[Map2T.scala 15:11]
  assign op_I0_8_1_0 = I0_8_1_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1_1 = I0_8_1_1; // @[Map2T.scala 15:11]
  assign op_I0_8_1_2 = I0_8_1_2; // @[Map2T.scala 15:11]
  assign op_I0_9_0_0 = I0_9_0_0; // @[Map2T.scala 15:11]
  assign op_I0_9_0_1 = I0_9_0_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0_2 = I0_9_0_2; // @[Map2T.scala 15:11]
  assign op_I0_9_1_0 = I0_9_1_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1_1 = I0_9_1_1; // @[Map2T.scala 15:11]
  assign op_I0_9_1_2 = I0_9_1_2; // @[Map2T.scala 15:11]
  assign op_I0_10_0_0 = I0_10_0_0; // @[Map2T.scala 15:11]
  assign op_I0_10_0_1 = I0_10_0_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0_2 = I0_10_0_2; // @[Map2T.scala 15:11]
  assign op_I0_10_1_0 = I0_10_1_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1_1 = I0_10_1_1; // @[Map2T.scala 15:11]
  assign op_I0_10_1_2 = I0_10_1_2; // @[Map2T.scala 15:11]
  assign op_I0_11_0_0 = I0_11_0_0; // @[Map2T.scala 15:11]
  assign op_I0_11_0_1 = I0_11_0_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0_2 = I0_11_0_2; // @[Map2T.scala 15:11]
  assign op_I0_11_1_0 = I0_11_1_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1_1 = I0_11_1_1; // @[Map2T.scala 15:11]
  assign op_I0_11_1_2 = I0_11_1_2; // @[Map2T.scala 15:11]
  assign op_I0_12_0_0 = I0_12_0_0; // @[Map2T.scala 15:11]
  assign op_I0_12_0_1 = I0_12_0_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0_2 = I0_12_0_2; // @[Map2T.scala 15:11]
  assign op_I0_12_1_0 = I0_12_1_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1_1 = I0_12_1_1; // @[Map2T.scala 15:11]
  assign op_I0_12_1_2 = I0_12_1_2; // @[Map2T.scala 15:11]
  assign op_I0_13_0_0 = I0_13_0_0; // @[Map2T.scala 15:11]
  assign op_I0_13_0_1 = I0_13_0_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0_2 = I0_13_0_2; // @[Map2T.scala 15:11]
  assign op_I0_13_1_0 = I0_13_1_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1_1 = I0_13_1_1; // @[Map2T.scala 15:11]
  assign op_I0_13_1_2 = I0_13_1_2; // @[Map2T.scala 15:11]
  assign op_I0_14_0_0 = I0_14_0_0; // @[Map2T.scala 15:11]
  assign op_I0_14_0_1 = I0_14_0_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0_2 = I0_14_0_2; // @[Map2T.scala 15:11]
  assign op_I0_14_1_0 = I0_14_1_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1_1 = I0_14_1_1; // @[Map2T.scala 15:11]
  assign op_I0_14_1_2 = I0_14_1_2; // @[Map2T.scala 15:11]
  assign op_I0_15_0_0 = I0_15_0_0; // @[Map2T.scala 15:11]
  assign op_I0_15_0_1 = I0_15_0_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0_2 = I0_15_0_2; // @[Map2T.scala 15:11]
  assign op_I0_15_1_0 = I0_15_1_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1_1 = I0_15_1_1; // @[Map2T.scala 15:11]
  assign op_I0_15_1_2 = I0_15_1_2; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_0_2 = I1_0_2; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_1_2 = I1_1_2; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_2_2 = I1_2_2; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_3_2 = I1_3_2; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_4_2 = I1_4_2; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_5_2 = I1_5_2; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_6_2 = I1_6_2; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_7_2 = I1_7_2; // @[Map2T.scala 16:11]
  assign op_I1_8_0 = I1_8_0; // @[Map2T.scala 16:11]
  assign op_I1_8_1 = I1_8_1; // @[Map2T.scala 16:11]
  assign op_I1_8_2 = I1_8_2; // @[Map2T.scala 16:11]
  assign op_I1_9_0 = I1_9_0; // @[Map2T.scala 16:11]
  assign op_I1_9_1 = I1_9_1; // @[Map2T.scala 16:11]
  assign op_I1_9_2 = I1_9_2; // @[Map2T.scala 16:11]
  assign op_I1_10_0 = I1_10_0; // @[Map2T.scala 16:11]
  assign op_I1_10_1 = I1_10_1; // @[Map2T.scala 16:11]
  assign op_I1_10_2 = I1_10_2; // @[Map2T.scala 16:11]
  assign op_I1_11_0 = I1_11_0; // @[Map2T.scala 16:11]
  assign op_I1_11_1 = I1_11_1; // @[Map2T.scala 16:11]
  assign op_I1_11_2 = I1_11_2; // @[Map2T.scala 16:11]
  assign op_I1_12_0 = I1_12_0; // @[Map2T.scala 16:11]
  assign op_I1_12_1 = I1_12_1; // @[Map2T.scala 16:11]
  assign op_I1_12_2 = I1_12_2; // @[Map2T.scala 16:11]
  assign op_I1_13_0 = I1_13_0; // @[Map2T.scala 16:11]
  assign op_I1_13_1 = I1_13_1; // @[Map2T.scala 16:11]
  assign op_I1_13_2 = I1_13_2; // @[Map2T.scala 16:11]
  assign op_I1_14_0 = I1_14_0; // @[Map2T.scala 16:11]
  assign op_I1_14_1 = I1_14_1; // @[Map2T.scala 16:11]
  assign op_I1_14_2 = I1_14_2; // @[Map2T.scala 16:11]
  assign op_I1_15_0 = I1_15_0; // @[Map2T.scala 16:11]
  assign op_I1_15_1 = I1_15_1; // @[Map2T.scala 16:11]
  assign op_I1_15_2 = I1_15_2; // @[Map2T.scala 16:11]
endmodule
module PartitionS_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_8_1_2,
  input  [7:0] I_8_2_0,
  input  [7:0] I_8_2_1,
  input  [7:0] I_8_2_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_9_1_2,
  input  [7:0] I_9_2_0,
  input  [7:0] I_9_2_1,
  input  [7:0] I_9_2_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_10_1_2,
  input  [7:0] I_10_2_0,
  input  [7:0] I_10_2_1,
  input  [7:0] I_10_2_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_11_1_2,
  input  [7:0] I_11_2_0,
  input  [7:0] I_11_2_1,
  input  [7:0] I_11_2_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_12_1_2,
  input  [7:0] I_12_2_0,
  input  [7:0] I_12_2_1,
  input  [7:0] I_12_2_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_13_1_2,
  input  [7:0] I_13_2_0,
  input  [7:0] I_13_2_1,
  input  [7:0] I_13_2_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_14_1_2,
  input  [7:0] I_14_2_0,
  input  [7:0] I_14_2_1,
  input  [7:0] I_14_2_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  input  [7:0] I_15_1_2,
  input  [7:0] I_15_2_0,
  input  [7:0] I_15_2_1,
  input  [7:0] I_15_2_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_2_0_2_0,
  output [7:0] O_2_0_2_1,
  output [7:0] O_2_0_2_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_3_0_2_0,
  output [7:0] O_3_0_2_1,
  output [7:0] O_3_0_2_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_4_0_2_0,
  output [7:0] O_4_0_2_1,
  output [7:0] O_4_0_2_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_5_0_2_0,
  output [7:0] O_5_0_2_1,
  output [7:0] O_5_0_2_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_6_0_2_0,
  output [7:0] O_6_0_2_1,
  output [7:0] O_6_0_2_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_7_0_2_0,
  output [7:0] O_7_0_2_1,
  output [7:0] O_7_0_2_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_8_0_1_2,
  output [7:0] O_8_0_2_0,
  output [7:0] O_8_0_2_1,
  output [7:0] O_8_0_2_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_9_0_1_2,
  output [7:0] O_9_0_2_0,
  output [7:0] O_9_0_2_1,
  output [7:0] O_9_0_2_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_10_0_1_2,
  output [7:0] O_10_0_2_0,
  output [7:0] O_10_0_2_1,
  output [7:0] O_10_0_2_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_11_0_1_2,
  output [7:0] O_11_0_2_0,
  output [7:0] O_11_0_2_1,
  output [7:0] O_11_0_2_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_12_0_1_2,
  output [7:0] O_12_0_2_0,
  output [7:0] O_12_0_2_1,
  output [7:0] O_12_0_2_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_13_0_1_2,
  output [7:0] O_13_0_2_0,
  output [7:0] O_13_0_2_1,
  output [7:0] O_13_0_2_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_14_0_1_2,
  output [7:0] O_14_0_2_0,
  output [7:0] O_14_0_2_1,
  output [7:0] O_14_0_2_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1,
  output [7:0] O_15_0_1_2,
  output [7:0] O_15_0_2_0,
  output [7:0] O_15_0_2_1,
  output [7:0] O_15_0_2_2
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_0_2 = I_0_0_2; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_0_0_1_2 = I_0_1_2; // @[Partition.scala 15:39]
  assign O_0_0_2_0 = I_0_2_0; // @[Partition.scala 15:39]
  assign O_0_0_2_1 = I_0_2_1; // @[Partition.scala 15:39]
  assign O_0_0_2_2 = I_0_2_2; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0_2 = I_1_0_2; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_1_0_1_2 = I_1_1_2; // @[Partition.scala 15:39]
  assign O_1_0_2_0 = I_1_2_0; // @[Partition.scala 15:39]
  assign O_1_0_2_1 = I_1_2_1; // @[Partition.scala 15:39]
  assign O_1_0_2_2 = I_1_2_2; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_0_2 = I_2_0_2; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_2_0_1_2 = I_2_1_2; // @[Partition.scala 15:39]
  assign O_2_0_2_0 = I_2_2_0; // @[Partition.scala 15:39]
  assign O_2_0_2_1 = I_2_2_1; // @[Partition.scala 15:39]
  assign O_2_0_2_2 = I_2_2_2; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_0_2 = I_3_0_2; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
  assign O_3_0_1_2 = I_3_1_2; // @[Partition.scala 15:39]
  assign O_3_0_2_0 = I_3_2_0; // @[Partition.scala 15:39]
  assign O_3_0_2_1 = I_3_2_1; // @[Partition.scala 15:39]
  assign O_3_0_2_2 = I_3_2_2; // @[Partition.scala 15:39]
  assign O_4_0_0_0 = I_4_0_0; // @[Partition.scala 15:39]
  assign O_4_0_0_1 = I_4_0_1; // @[Partition.scala 15:39]
  assign O_4_0_0_2 = I_4_0_2; // @[Partition.scala 15:39]
  assign O_4_0_1_0 = I_4_1_0; // @[Partition.scala 15:39]
  assign O_4_0_1_1 = I_4_1_1; // @[Partition.scala 15:39]
  assign O_4_0_1_2 = I_4_1_2; // @[Partition.scala 15:39]
  assign O_4_0_2_0 = I_4_2_0; // @[Partition.scala 15:39]
  assign O_4_0_2_1 = I_4_2_1; // @[Partition.scala 15:39]
  assign O_4_0_2_2 = I_4_2_2; // @[Partition.scala 15:39]
  assign O_5_0_0_0 = I_5_0_0; // @[Partition.scala 15:39]
  assign O_5_0_0_1 = I_5_0_1; // @[Partition.scala 15:39]
  assign O_5_0_0_2 = I_5_0_2; // @[Partition.scala 15:39]
  assign O_5_0_1_0 = I_5_1_0; // @[Partition.scala 15:39]
  assign O_5_0_1_1 = I_5_1_1; // @[Partition.scala 15:39]
  assign O_5_0_1_2 = I_5_1_2; // @[Partition.scala 15:39]
  assign O_5_0_2_0 = I_5_2_0; // @[Partition.scala 15:39]
  assign O_5_0_2_1 = I_5_2_1; // @[Partition.scala 15:39]
  assign O_5_0_2_2 = I_5_2_2; // @[Partition.scala 15:39]
  assign O_6_0_0_0 = I_6_0_0; // @[Partition.scala 15:39]
  assign O_6_0_0_1 = I_6_0_1; // @[Partition.scala 15:39]
  assign O_6_0_0_2 = I_6_0_2; // @[Partition.scala 15:39]
  assign O_6_0_1_0 = I_6_1_0; // @[Partition.scala 15:39]
  assign O_6_0_1_1 = I_6_1_1; // @[Partition.scala 15:39]
  assign O_6_0_1_2 = I_6_1_2; // @[Partition.scala 15:39]
  assign O_6_0_2_0 = I_6_2_0; // @[Partition.scala 15:39]
  assign O_6_0_2_1 = I_6_2_1; // @[Partition.scala 15:39]
  assign O_6_0_2_2 = I_6_2_2; // @[Partition.scala 15:39]
  assign O_7_0_0_0 = I_7_0_0; // @[Partition.scala 15:39]
  assign O_7_0_0_1 = I_7_0_1; // @[Partition.scala 15:39]
  assign O_7_0_0_2 = I_7_0_2; // @[Partition.scala 15:39]
  assign O_7_0_1_0 = I_7_1_0; // @[Partition.scala 15:39]
  assign O_7_0_1_1 = I_7_1_1; // @[Partition.scala 15:39]
  assign O_7_0_1_2 = I_7_1_2; // @[Partition.scala 15:39]
  assign O_7_0_2_0 = I_7_2_0; // @[Partition.scala 15:39]
  assign O_7_0_2_1 = I_7_2_1; // @[Partition.scala 15:39]
  assign O_7_0_2_2 = I_7_2_2; // @[Partition.scala 15:39]
  assign O_8_0_0_0 = I_8_0_0; // @[Partition.scala 15:39]
  assign O_8_0_0_1 = I_8_0_1; // @[Partition.scala 15:39]
  assign O_8_0_0_2 = I_8_0_2; // @[Partition.scala 15:39]
  assign O_8_0_1_0 = I_8_1_0; // @[Partition.scala 15:39]
  assign O_8_0_1_1 = I_8_1_1; // @[Partition.scala 15:39]
  assign O_8_0_1_2 = I_8_1_2; // @[Partition.scala 15:39]
  assign O_8_0_2_0 = I_8_2_0; // @[Partition.scala 15:39]
  assign O_8_0_2_1 = I_8_2_1; // @[Partition.scala 15:39]
  assign O_8_0_2_2 = I_8_2_2; // @[Partition.scala 15:39]
  assign O_9_0_0_0 = I_9_0_0; // @[Partition.scala 15:39]
  assign O_9_0_0_1 = I_9_0_1; // @[Partition.scala 15:39]
  assign O_9_0_0_2 = I_9_0_2; // @[Partition.scala 15:39]
  assign O_9_0_1_0 = I_9_1_0; // @[Partition.scala 15:39]
  assign O_9_0_1_1 = I_9_1_1; // @[Partition.scala 15:39]
  assign O_9_0_1_2 = I_9_1_2; // @[Partition.scala 15:39]
  assign O_9_0_2_0 = I_9_2_0; // @[Partition.scala 15:39]
  assign O_9_0_2_1 = I_9_2_1; // @[Partition.scala 15:39]
  assign O_9_0_2_2 = I_9_2_2; // @[Partition.scala 15:39]
  assign O_10_0_0_0 = I_10_0_0; // @[Partition.scala 15:39]
  assign O_10_0_0_1 = I_10_0_1; // @[Partition.scala 15:39]
  assign O_10_0_0_2 = I_10_0_2; // @[Partition.scala 15:39]
  assign O_10_0_1_0 = I_10_1_0; // @[Partition.scala 15:39]
  assign O_10_0_1_1 = I_10_1_1; // @[Partition.scala 15:39]
  assign O_10_0_1_2 = I_10_1_2; // @[Partition.scala 15:39]
  assign O_10_0_2_0 = I_10_2_0; // @[Partition.scala 15:39]
  assign O_10_0_2_1 = I_10_2_1; // @[Partition.scala 15:39]
  assign O_10_0_2_2 = I_10_2_2; // @[Partition.scala 15:39]
  assign O_11_0_0_0 = I_11_0_0; // @[Partition.scala 15:39]
  assign O_11_0_0_1 = I_11_0_1; // @[Partition.scala 15:39]
  assign O_11_0_0_2 = I_11_0_2; // @[Partition.scala 15:39]
  assign O_11_0_1_0 = I_11_1_0; // @[Partition.scala 15:39]
  assign O_11_0_1_1 = I_11_1_1; // @[Partition.scala 15:39]
  assign O_11_0_1_2 = I_11_1_2; // @[Partition.scala 15:39]
  assign O_11_0_2_0 = I_11_2_0; // @[Partition.scala 15:39]
  assign O_11_0_2_1 = I_11_2_1; // @[Partition.scala 15:39]
  assign O_11_0_2_2 = I_11_2_2; // @[Partition.scala 15:39]
  assign O_12_0_0_0 = I_12_0_0; // @[Partition.scala 15:39]
  assign O_12_0_0_1 = I_12_0_1; // @[Partition.scala 15:39]
  assign O_12_0_0_2 = I_12_0_2; // @[Partition.scala 15:39]
  assign O_12_0_1_0 = I_12_1_0; // @[Partition.scala 15:39]
  assign O_12_0_1_1 = I_12_1_1; // @[Partition.scala 15:39]
  assign O_12_0_1_2 = I_12_1_2; // @[Partition.scala 15:39]
  assign O_12_0_2_0 = I_12_2_0; // @[Partition.scala 15:39]
  assign O_12_0_2_1 = I_12_2_1; // @[Partition.scala 15:39]
  assign O_12_0_2_2 = I_12_2_2; // @[Partition.scala 15:39]
  assign O_13_0_0_0 = I_13_0_0; // @[Partition.scala 15:39]
  assign O_13_0_0_1 = I_13_0_1; // @[Partition.scala 15:39]
  assign O_13_0_0_2 = I_13_0_2; // @[Partition.scala 15:39]
  assign O_13_0_1_0 = I_13_1_0; // @[Partition.scala 15:39]
  assign O_13_0_1_1 = I_13_1_1; // @[Partition.scala 15:39]
  assign O_13_0_1_2 = I_13_1_2; // @[Partition.scala 15:39]
  assign O_13_0_2_0 = I_13_2_0; // @[Partition.scala 15:39]
  assign O_13_0_2_1 = I_13_2_1; // @[Partition.scala 15:39]
  assign O_13_0_2_2 = I_13_2_2; // @[Partition.scala 15:39]
  assign O_14_0_0_0 = I_14_0_0; // @[Partition.scala 15:39]
  assign O_14_0_0_1 = I_14_0_1; // @[Partition.scala 15:39]
  assign O_14_0_0_2 = I_14_0_2; // @[Partition.scala 15:39]
  assign O_14_0_1_0 = I_14_1_0; // @[Partition.scala 15:39]
  assign O_14_0_1_1 = I_14_1_1; // @[Partition.scala 15:39]
  assign O_14_0_1_2 = I_14_1_2; // @[Partition.scala 15:39]
  assign O_14_0_2_0 = I_14_2_0; // @[Partition.scala 15:39]
  assign O_14_0_2_1 = I_14_2_1; // @[Partition.scala 15:39]
  assign O_14_0_2_2 = I_14_2_2; // @[Partition.scala 15:39]
  assign O_15_0_0_0 = I_15_0_0; // @[Partition.scala 15:39]
  assign O_15_0_0_1 = I_15_0_1; // @[Partition.scala 15:39]
  assign O_15_0_0_2 = I_15_0_2; // @[Partition.scala 15:39]
  assign O_15_0_1_0 = I_15_1_0; // @[Partition.scala 15:39]
  assign O_15_0_1_1 = I_15_1_1; // @[Partition.scala 15:39]
  assign O_15_0_1_2 = I_15_1_2; // @[Partition.scala 15:39]
  assign O_15_0_2_0 = I_15_2_0; // @[Partition.scala 15:39]
  assign O_15_0_2_1 = I_15_2_1; // @[Partition.scala 15:39]
  assign O_15_0_2_2 = I_15_2_2; // @[Partition.scala 15:39]
endmodule
module MapT_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_8_1_2,
  input  [7:0] I_8_2_0,
  input  [7:0] I_8_2_1,
  input  [7:0] I_8_2_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_9_1_2,
  input  [7:0] I_9_2_0,
  input  [7:0] I_9_2_1,
  input  [7:0] I_9_2_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_10_1_2,
  input  [7:0] I_10_2_0,
  input  [7:0] I_10_2_1,
  input  [7:0] I_10_2_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_11_1_2,
  input  [7:0] I_11_2_0,
  input  [7:0] I_11_2_1,
  input  [7:0] I_11_2_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_12_1_2,
  input  [7:0] I_12_2_0,
  input  [7:0] I_12_2_1,
  input  [7:0] I_12_2_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_13_1_2,
  input  [7:0] I_13_2_0,
  input  [7:0] I_13_2_1,
  input  [7:0] I_13_2_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_14_1_2,
  input  [7:0] I_14_2_0,
  input  [7:0] I_14_2_1,
  input  [7:0] I_14_2_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  input  [7:0] I_15_1_2,
  input  [7:0] I_15_2_0,
  input  [7:0] I_15_2_1,
  input  [7:0] I_15_2_2,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_0_2,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_0_0_1_2,
  output [7:0] O_0_0_2_0,
  output [7:0] O_0_0_2_1,
  output [7:0] O_0_0_2_2,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_0_2,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_1_0_1_2,
  output [7:0] O_1_0_2_0,
  output [7:0] O_1_0_2_1,
  output [7:0] O_1_0_2_2,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_0_2,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_2_0_1_2,
  output [7:0] O_2_0_2_0,
  output [7:0] O_2_0_2_1,
  output [7:0] O_2_0_2_2,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_0_2,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_3_0_1_2,
  output [7:0] O_3_0_2_0,
  output [7:0] O_3_0_2_1,
  output [7:0] O_3_0_2_2,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_0_2,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_4_0_1_2,
  output [7:0] O_4_0_2_0,
  output [7:0] O_4_0_2_1,
  output [7:0] O_4_0_2_2,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_0_2,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_5_0_1_2,
  output [7:0] O_5_0_2_0,
  output [7:0] O_5_0_2_1,
  output [7:0] O_5_0_2_2,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_0_2,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_6_0_1_2,
  output [7:0] O_6_0_2_0,
  output [7:0] O_6_0_2_1,
  output [7:0] O_6_0_2_2,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_0_2,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_7_0_1_2,
  output [7:0] O_7_0_2_0,
  output [7:0] O_7_0_2_1,
  output [7:0] O_7_0_2_2,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_0_2,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_8_0_1_2,
  output [7:0] O_8_0_2_0,
  output [7:0] O_8_0_2_1,
  output [7:0] O_8_0_2_2,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_0_2,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_9_0_1_2,
  output [7:0] O_9_0_2_0,
  output [7:0] O_9_0_2_1,
  output [7:0] O_9_0_2_2,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_0_2,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_10_0_1_2,
  output [7:0] O_10_0_2_0,
  output [7:0] O_10_0_2_1,
  output [7:0] O_10_0_2_2,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_0_2,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_11_0_1_2,
  output [7:0] O_11_0_2_0,
  output [7:0] O_11_0_2_1,
  output [7:0] O_11_0_2_2,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_0_2,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_12_0_1_2,
  output [7:0] O_12_0_2_0,
  output [7:0] O_12_0_2_1,
  output [7:0] O_12_0_2_2,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_0_2,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_13_0_1_2,
  output [7:0] O_13_0_2_0,
  output [7:0] O_13_0_2_1,
  output [7:0] O_13_0_2_2,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_0_2,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_14_0_1_2,
  output [7:0] O_14_0_2_0,
  output [7:0] O_14_0_2_1,
  output [7:0] O_14_0_2_2,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_0_2,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1,
  output [7:0] O_15_0_1_2,
  output [7:0] O_15_0_2_0,
  output [7:0] O_15_0_2_1,
  output [7:0] O_15_0_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_2_2; // @[MapT.scala 8:20]
  PartitionS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_8_1_2(op_I_8_1_2),
    .I_8_2_0(op_I_8_2_0),
    .I_8_2_1(op_I_8_2_1),
    .I_8_2_2(op_I_8_2_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_9_1_2(op_I_9_1_2),
    .I_9_2_0(op_I_9_2_0),
    .I_9_2_1(op_I_9_2_1),
    .I_9_2_2(op_I_9_2_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_10_1_2(op_I_10_1_2),
    .I_10_2_0(op_I_10_2_0),
    .I_10_2_1(op_I_10_2_1),
    .I_10_2_2(op_I_10_2_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_11_1_2(op_I_11_1_2),
    .I_11_2_0(op_I_11_2_0),
    .I_11_2_1(op_I_11_2_1),
    .I_11_2_2(op_I_11_2_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_12_1_2(op_I_12_1_2),
    .I_12_2_0(op_I_12_2_0),
    .I_12_2_1(op_I_12_2_1),
    .I_12_2_2(op_I_12_2_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_13_1_2(op_I_13_1_2),
    .I_13_2_0(op_I_13_2_0),
    .I_13_2_1(op_I_13_2_1),
    .I_13_2_2(op_I_13_2_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_14_1_2(op_I_14_1_2),
    .I_14_2_0(op_I_14_2_0),
    .I_14_2_1(op_I_14_2_1),
    .I_14_2_2(op_I_14_2_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .I_15_1_2(op_I_15_1_2),
    .I_15_2_0(op_I_15_2_0),
    .I_15_2_1(op_I_15_2_1),
    .I_15_2_2(op_I_15_2_2),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_0_2(op_O_0_0_0_2),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_0_0_1_2(op_O_0_0_1_2),
    .O_0_0_2_0(op_O_0_0_2_0),
    .O_0_0_2_1(op_O_0_0_2_1),
    .O_0_0_2_2(op_O_0_0_2_2),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_0_2(op_O_1_0_0_2),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_1_0_1_2(op_O_1_0_1_2),
    .O_1_0_2_0(op_O_1_0_2_0),
    .O_1_0_2_1(op_O_1_0_2_1),
    .O_1_0_2_2(op_O_1_0_2_2),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_0_2(op_O_2_0_0_2),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_2_0_1_2(op_O_2_0_1_2),
    .O_2_0_2_0(op_O_2_0_2_0),
    .O_2_0_2_1(op_O_2_0_2_1),
    .O_2_0_2_2(op_O_2_0_2_2),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_0_2(op_O_3_0_0_2),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_3_0_1_2(op_O_3_0_1_2),
    .O_3_0_2_0(op_O_3_0_2_0),
    .O_3_0_2_1(op_O_3_0_2_1),
    .O_3_0_2_2(op_O_3_0_2_2),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_0_2(op_O_4_0_0_2),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_4_0_1_2(op_O_4_0_1_2),
    .O_4_0_2_0(op_O_4_0_2_0),
    .O_4_0_2_1(op_O_4_0_2_1),
    .O_4_0_2_2(op_O_4_0_2_2),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_0_2(op_O_5_0_0_2),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_5_0_1_2(op_O_5_0_1_2),
    .O_5_0_2_0(op_O_5_0_2_0),
    .O_5_0_2_1(op_O_5_0_2_1),
    .O_5_0_2_2(op_O_5_0_2_2),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_0_2(op_O_6_0_0_2),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_6_0_1_2(op_O_6_0_1_2),
    .O_6_0_2_0(op_O_6_0_2_0),
    .O_6_0_2_1(op_O_6_0_2_1),
    .O_6_0_2_2(op_O_6_0_2_2),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_0_2(op_O_7_0_0_2),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_7_0_1_2(op_O_7_0_1_2),
    .O_7_0_2_0(op_O_7_0_2_0),
    .O_7_0_2_1(op_O_7_0_2_1),
    .O_7_0_2_2(op_O_7_0_2_2),
    .O_8_0_0_0(op_O_8_0_0_0),
    .O_8_0_0_1(op_O_8_0_0_1),
    .O_8_0_0_2(op_O_8_0_0_2),
    .O_8_0_1_0(op_O_8_0_1_0),
    .O_8_0_1_1(op_O_8_0_1_1),
    .O_8_0_1_2(op_O_8_0_1_2),
    .O_8_0_2_0(op_O_8_0_2_0),
    .O_8_0_2_1(op_O_8_0_2_1),
    .O_8_0_2_2(op_O_8_0_2_2),
    .O_9_0_0_0(op_O_9_0_0_0),
    .O_9_0_0_1(op_O_9_0_0_1),
    .O_9_0_0_2(op_O_9_0_0_2),
    .O_9_0_1_0(op_O_9_0_1_0),
    .O_9_0_1_1(op_O_9_0_1_1),
    .O_9_0_1_2(op_O_9_0_1_2),
    .O_9_0_2_0(op_O_9_0_2_0),
    .O_9_0_2_1(op_O_9_0_2_1),
    .O_9_0_2_2(op_O_9_0_2_2),
    .O_10_0_0_0(op_O_10_0_0_0),
    .O_10_0_0_1(op_O_10_0_0_1),
    .O_10_0_0_2(op_O_10_0_0_2),
    .O_10_0_1_0(op_O_10_0_1_0),
    .O_10_0_1_1(op_O_10_0_1_1),
    .O_10_0_1_2(op_O_10_0_1_2),
    .O_10_0_2_0(op_O_10_0_2_0),
    .O_10_0_2_1(op_O_10_0_2_1),
    .O_10_0_2_2(op_O_10_0_2_2),
    .O_11_0_0_0(op_O_11_0_0_0),
    .O_11_0_0_1(op_O_11_0_0_1),
    .O_11_0_0_2(op_O_11_0_0_2),
    .O_11_0_1_0(op_O_11_0_1_0),
    .O_11_0_1_1(op_O_11_0_1_1),
    .O_11_0_1_2(op_O_11_0_1_2),
    .O_11_0_2_0(op_O_11_0_2_0),
    .O_11_0_2_1(op_O_11_0_2_1),
    .O_11_0_2_2(op_O_11_0_2_2),
    .O_12_0_0_0(op_O_12_0_0_0),
    .O_12_0_0_1(op_O_12_0_0_1),
    .O_12_0_0_2(op_O_12_0_0_2),
    .O_12_0_1_0(op_O_12_0_1_0),
    .O_12_0_1_1(op_O_12_0_1_1),
    .O_12_0_1_2(op_O_12_0_1_2),
    .O_12_0_2_0(op_O_12_0_2_0),
    .O_12_0_2_1(op_O_12_0_2_1),
    .O_12_0_2_2(op_O_12_0_2_2),
    .O_13_0_0_0(op_O_13_0_0_0),
    .O_13_0_0_1(op_O_13_0_0_1),
    .O_13_0_0_2(op_O_13_0_0_2),
    .O_13_0_1_0(op_O_13_0_1_0),
    .O_13_0_1_1(op_O_13_0_1_1),
    .O_13_0_1_2(op_O_13_0_1_2),
    .O_13_0_2_0(op_O_13_0_2_0),
    .O_13_0_2_1(op_O_13_0_2_1),
    .O_13_0_2_2(op_O_13_0_2_2),
    .O_14_0_0_0(op_O_14_0_0_0),
    .O_14_0_0_1(op_O_14_0_0_1),
    .O_14_0_0_2(op_O_14_0_0_2),
    .O_14_0_1_0(op_O_14_0_1_0),
    .O_14_0_1_1(op_O_14_0_1_1),
    .O_14_0_1_2(op_O_14_0_1_2),
    .O_14_0_2_0(op_O_14_0_2_0),
    .O_14_0_2_1(op_O_14_0_2_1),
    .O_14_0_2_2(op_O_14_0_2_2),
    .O_15_0_0_0(op_O_15_0_0_0),
    .O_15_0_0_1(op_O_15_0_0_1),
    .O_15_0_0_2(op_O_15_0_0_2),
    .O_15_0_1_0(op_O_15_0_1_0),
    .O_15_0_1_1(op_O_15_0_1_1),
    .O_15_0_1_2(op_O_15_0_1_2),
    .O_15_0_2_0(op_O_15_0_2_0),
    .O_15_0_2_1(op_O_15_0_2_1),
    .O_15_0_2_2(op_O_15_0_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_0_2 = op_O_0_0_0_2; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_0_0_1_2 = op_O_0_0_1_2; // @[MapT.scala 15:7]
  assign O_0_0_2_0 = op_O_0_0_2_0; // @[MapT.scala 15:7]
  assign O_0_0_2_1 = op_O_0_0_2_1; // @[MapT.scala 15:7]
  assign O_0_0_2_2 = op_O_0_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0_2 = op_O_1_0_0_2; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_1_2 = op_O_1_0_1_2; // @[MapT.scala 15:7]
  assign O_1_0_2_0 = op_O_1_0_2_0; // @[MapT.scala 15:7]
  assign O_1_0_2_1 = op_O_1_0_2_1; // @[MapT.scala 15:7]
  assign O_1_0_2_2 = op_O_1_0_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[MapT.scala 15:7]
  assign O_2_0_0_2 = op_O_2_0_0_2; // @[MapT.scala 15:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[MapT.scala 15:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[MapT.scala 15:7]
  assign O_2_0_1_2 = op_O_2_0_1_2; // @[MapT.scala 15:7]
  assign O_2_0_2_0 = op_O_2_0_2_0; // @[MapT.scala 15:7]
  assign O_2_0_2_1 = op_O_2_0_2_1; // @[MapT.scala 15:7]
  assign O_2_0_2_2 = op_O_2_0_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[MapT.scala 15:7]
  assign O_3_0_0_2 = op_O_3_0_0_2; // @[MapT.scala 15:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[MapT.scala 15:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[MapT.scala 15:7]
  assign O_3_0_1_2 = op_O_3_0_1_2; // @[MapT.scala 15:7]
  assign O_3_0_2_0 = op_O_3_0_2_0; // @[MapT.scala 15:7]
  assign O_3_0_2_1 = op_O_3_0_2_1; // @[MapT.scala 15:7]
  assign O_3_0_2_2 = op_O_3_0_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[MapT.scala 15:7]
  assign O_4_0_0_2 = op_O_4_0_0_2; // @[MapT.scala 15:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[MapT.scala 15:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[MapT.scala 15:7]
  assign O_4_0_1_2 = op_O_4_0_1_2; // @[MapT.scala 15:7]
  assign O_4_0_2_0 = op_O_4_0_2_0; // @[MapT.scala 15:7]
  assign O_4_0_2_1 = op_O_4_0_2_1; // @[MapT.scala 15:7]
  assign O_4_0_2_2 = op_O_4_0_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[MapT.scala 15:7]
  assign O_5_0_0_2 = op_O_5_0_0_2; // @[MapT.scala 15:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[MapT.scala 15:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[MapT.scala 15:7]
  assign O_5_0_1_2 = op_O_5_0_1_2; // @[MapT.scala 15:7]
  assign O_5_0_2_0 = op_O_5_0_2_0; // @[MapT.scala 15:7]
  assign O_5_0_2_1 = op_O_5_0_2_1; // @[MapT.scala 15:7]
  assign O_5_0_2_2 = op_O_5_0_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[MapT.scala 15:7]
  assign O_6_0_0_2 = op_O_6_0_0_2; // @[MapT.scala 15:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[MapT.scala 15:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[MapT.scala 15:7]
  assign O_6_0_1_2 = op_O_6_0_1_2; // @[MapT.scala 15:7]
  assign O_6_0_2_0 = op_O_6_0_2_0; // @[MapT.scala 15:7]
  assign O_6_0_2_1 = op_O_6_0_2_1; // @[MapT.scala 15:7]
  assign O_6_0_2_2 = op_O_6_0_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[MapT.scala 15:7]
  assign O_7_0_0_2 = op_O_7_0_0_2; // @[MapT.scala 15:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[MapT.scala 15:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[MapT.scala 15:7]
  assign O_7_0_1_2 = op_O_7_0_1_2; // @[MapT.scala 15:7]
  assign O_7_0_2_0 = op_O_7_0_2_0; // @[MapT.scala 15:7]
  assign O_7_0_2_1 = op_O_7_0_2_1; // @[MapT.scala 15:7]
  assign O_7_0_2_2 = op_O_7_0_2_2; // @[MapT.scala 15:7]
  assign O_8_0_0_0 = op_O_8_0_0_0; // @[MapT.scala 15:7]
  assign O_8_0_0_1 = op_O_8_0_0_1; // @[MapT.scala 15:7]
  assign O_8_0_0_2 = op_O_8_0_0_2; // @[MapT.scala 15:7]
  assign O_8_0_1_0 = op_O_8_0_1_0; // @[MapT.scala 15:7]
  assign O_8_0_1_1 = op_O_8_0_1_1; // @[MapT.scala 15:7]
  assign O_8_0_1_2 = op_O_8_0_1_2; // @[MapT.scala 15:7]
  assign O_8_0_2_0 = op_O_8_0_2_0; // @[MapT.scala 15:7]
  assign O_8_0_2_1 = op_O_8_0_2_1; // @[MapT.scala 15:7]
  assign O_8_0_2_2 = op_O_8_0_2_2; // @[MapT.scala 15:7]
  assign O_9_0_0_0 = op_O_9_0_0_0; // @[MapT.scala 15:7]
  assign O_9_0_0_1 = op_O_9_0_0_1; // @[MapT.scala 15:7]
  assign O_9_0_0_2 = op_O_9_0_0_2; // @[MapT.scala 15:7]
  assign O_9_0_1_0 = op_O_9_0_1_0; // @[MapT.scala 15:7]
  assign O_9_0_1_1 = op_O_9_0_1_1; // @[MapT.scala 15:7]
  assign O_9_0_1_2 = op_O_9_0_1_2; // @[MapT.scala 15:7]
  assign O_9_0_2_0 = op_O_9_0_2_0; // @[MapT.scala 15:7]
  assign O_9_0_2_1 = op_O_9_0_2_1; // @[MapT.scala 15:7]
  assign O_9_0_2_2 = op_O_9_0_2_2; // @[MapT.scala 15:7]
  assign O_10_0_0_0 = op_O_10_0_0_0; // @[MapT.scala 15:7]
  assign O_10_0_0_1 = op_O_10_0_0_1; // @[MapT.scala 15:7]
  assign O_10_0_0_2 = op_O_10_0_0_2; // @[MapT.scala 15:7]
  assign O_10_0_1_0 = op_O_10_0_1_0; // @[MapT.scala 15:7]
  assign O_10_0_1_1 = op_O_10_0_1_1; // @[MapT.scala 15:7]
  assign O_10_0_1_2 = op_O_10_0_1_2; // @[MapT.scala 15:7]
  assign O_10_0_2_0 = op_O_10_0_2_0; // @[MapT.scala 15:7]
  assign O_10_0_2_1 = op_O_10_0_2_1; // @[MapT.scala 15:7]
  assign O_10_0_2_2 = op_O_10_0_2_2; // @[MapT.scala 15:7]
  assign O_11_0_0_0 = op_O_11_0_0_0; // @[MapT.scala 15:7]
  assign O_11_0_0_1 = op_O_11_0_0_1; // @[MapT.scala 15:7]
  assign O_11_0_0_2 = op_O_11_0_0_2; // @[MapT.scala 15:7]
  assign O_11_0_1_0 = op_O_11_0_1_0; // @[MapT.scala 15:7]
  assign O_11_0_1_1 = op_O_11_0_1_1; // @[MapT.scala 15:7]
  assign O_11_0_1_2 = op_O_11_0_1_2; // @[MapT.scala 15:7]
  assign O_11_0_2_0 = op_O_11_0_2_0; // @[MapT.scala 15:7]
  assign O_11_0_2_1 = op_O_11_0_2_1; // @[MapT.scala 15:7]
  assign O_11_0_2_2 = op_O_11_0_2_2; // @[MapT.scala 15:7]
  assign O_12_0_0_0 = op_O_12_0_0_0; // @[MapT.scala 15:7]
  assign O_12_0_0_1 = op_O_12_0_0_1; // @[MapT.scala 15:7]
  assign O_12_0_0_2 = op_O_12_0_0_2; // @[MapT.scala 15:7]
  assign O_12_0_1_0 = op_O_12_0_1_0; // @[MapT.scala 15:7]
  assign O_12_0_1_1 = op_O_12_0_1_1; // @[MapT.scala 15:7]
  assign O_12_0_1_2 = op_O_12_0_1_2; // @[MapT.scala 15:7]
  assign O_12_0_2_0 = op_O_12_0_2_0; // @[MapT.scala 15:7]
  assign O_12_0_2_1 = op_O_12_0_2_1; // @[MapT.scala 15:7]
  assign O_12_0_2_2 = op_O_12_0_2_2; // @[MapT.scala 15:7]
  assign O_13_0_0_0 = op_O_13_0_0_0; // @[MapT.scala 15:7]
  assign O_13_0_0_1 = op_O_13_0_0_1; // @[MapT.scala 15:7]
  assign O_13_0_0_2 = op_O_13_0_0_2; // @[MapT.scala 15:7]
  assign O_13_0_1_0 = op_O_13_0_1_0; // @[MapT.scala 15:7]
  assign O_13_0_1_1 = op_O_13_0_1_1; // @[MapT.scala 15:7]
  assign O_13_0_1_2 = op_O_13_0_1_2; // @[MapT.scala 15:7]
  assign O_13_0_2_0 = op_O_13_0_2_0; // @[MapT.scala 15:7]
  assign O_13_0_2_1 = op_O_13_0_2_1; // @[MapT.scala 15:7]
  assign O_13_0_2_2 = op_O_13_0_2_2; // @[MapT.scala 15:7]
  assign O_14_0_0_0 = op_O_14_0_0_0; // @[MapT.scala 15:7]
  assign O_14_0_0_1 = op_O_14_0_0_1; // @[MapT.scala 15:7]
  assign O_14_0_0_2 = op_O_14_0_0_2; // @[MapT.scala 15:7]
  assign O_14_0_1_0 = op_O_14_0_1_0; // @[MapT.scala 15:7]
  assign O_14_0_1_1 = op_O_14_0_1_1; // @[MapT.scala 15:7]
  assign O_14_0_1_2 = op_O_14_0_1_2; // @[MapT.scala 15:7]
  assign O_14_0_2_0 = op_O_14_0_2_0; // @[MapT.scala 15:7]
  assign O_14_0_2_1 = op_O_14_0_2_1; // @[MapT.scala 15:7]
  assign O_14_0_2_2 = op_O_14_0_2_2; // @[MapT.scala 15:7]
  assign O_15_0_0_0 = op_O_15_0_0_0; // @[MapT.scala 15:7]
  assign O_15_0_0_1 = op_O_15_0_0_1; // @[MapT.scala 15:7]
  assign O_15_0_0_2 = op_O_15_0_0_2; // @[MapT.scala 15:7]
  assign O_15_0_1_0 = op_O_15_0_1_0; // @[MapT.scala 15:7]
  assign O_15_0_1_1 = op_O_15_0_1_1; // @[MapT.scala 15:7]
  assign O_15_0_1_2 = op_O_15_0_1_2; // @[MapT.scala 15:7]
  assign O_15_0_2_0 = op_O_15_0_2_0; // @[MapT.scala 15:7]
  assign O_15_0_2_1 = op_O_15_0_2_1; // @[MapT.scala 15:7]
  assign O_15_0_2_2 = op_O_15_0_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_8_1_2 = I_8_1_2; // @[MapT.scala 14:10]
  assign op_I_8_2_0 = I_8_2_0; // @[MapT.scala 14:10]
  assign op_I_8_2_1 = I_8_2_1; // @[MapT.scala 14:10]
  assign op_I_8_2_2 = I_8_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_9_1_2 = I_9_1_2; // @[MapT.scala 14:10]
  assign op_I_9_2_0 = I_9_2_0; // @[MapT.scala 14:10]
  assign op_I_9_2_1 = I_9_2_1; // @[MapT.scala 14:10]
  assign op_I_9_2_2 = I_9_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_10_1_2 = I_10_1_2; // @[MapT.scala 14:10]
  assign op_I_10_2_0 = I_10_2_0; // @[MapT.scala 14:10]
  assign op_I_10_2_1 = I_10_2_1; // @[MapT.scala 14:10]
  assign op_I_10_2_2 = I_10_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_11_1_2 = I_11_1_2; // @[MapT.scala 14:10]
  assign op_I_11_2_0 = I_11_2_0; // @[MapT.scala 14:10]
  assign op_I_11_2_1 = I_11_2_1; // @[MapT.scala 14:10]
  assign op_I_11_2_2 = I_11_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_12_1_2 = I_12_1_2; // @[MapT.scala 14:10]
  assign op_I_12_2_0 = I_12_2_0; // @[MapT.scala 14:10]
  assign op_I_12_2_1 = I_12_2_1; // @[MapT.scala 14:10]
  assign op_I_12_2_2 = I_12_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_13_1_2 = I_13_1_2; // @[MapT.scala 14:10]
  assign op_I_13_2_0 = I_13_2_0; // @[MapT.scala 14:10]
  assign op_I_13_2_1 = I_13_2_1; // @[MapT.scala 14:10]
  assign op_I_13_2_2 = I_13_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_14_1_2 = I_14_1_2; // @[MapT.scala 14:10]
  assign op_I_14_2_0 = I_14_2_0; // @[MapT.scala 14:10]
  assign op_I_14_2_1 = I_14_2_1; // @[MapT.scala 14:10]
  assign op_I_14_2_2 = I_14_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
  assign op_I_15_1_2 = I_15_1_2; // @[MapT.scala 14:10]
  assign op_I_15_2_0 = I_15_2_0; // @[MapT.scala 14:10]
  assign op_I_15_2_1 = I_15_2_1; // @[MapT.scala 14:10]
  assign op_I_15_2_2 = I_15_2_2; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_0_2 = I_0_2; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
  assign O_1_2 = I_1_2; // @[Tuple.scala 41:5]
  assign O_2_0 = I_2_0; // @[Tuple.scala 41:5]
  assign O_2_1 = I_2_1; // @[Tuple.scala 41:5]
  assign O_2_2 = I_2_2; // @[Tuple.scala 41:5]
endmodule
module Remove1S_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_2_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_2; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_2_2; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_3 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_0_2(op_inst_I_0_2),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .I_1_2(op_inst_I_1_2),
    .I_2_0(op_inst_I_2_0),
    .I_2_1(op_inst_I_2_1),
    .I_2_2(op_inst_I_2_2),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_0_2(op_inst_O_0_2),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1),
    .O_1_2(op_inst_O_1_2),
    .O_2_0(op_inst_O_2_0),
    .O_2_1(op_inst_O_2_1),
    .O_2_2(op_inst_O_2_2)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_0_2 = op_inst_O_0_2; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign O_1_2 = op_inst_O_1_2; // @[Remove1S.scala 14:5]
  assign O_2_0 = op_inst_O_2_0; // @[Remove1S.scala 14:5]
  assign O_2_1 = op_inst_O_2_1; // @[Remove1S.scala 14:5]
  assign O_2_2 = op_inst_O_2_2; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_2 = I_0_0_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_2 = I_0_1_2; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_0 = I_0_2_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_1 = I_0_2_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_2_2 = I_0_2_2; // @[Remove1S.scala 13:13]
endmodule
module MapS_3(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_2_0_1_2,
  input  [7:0] I_2_0_2_0,
  input  [7:0] I_2_0_2_1,
  input  [7:0] I_2_0_2_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_3_0_1_2,
  input  [7:0] I_3_0_2_0,
  input  [7:0] I_3_0_2_1,
  input  [7:0] I_3_0_2_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_4_0_1_2,
  input  [7:0] I_4_0_2_0,
  input  [7:0] I_4_0_2_1,
  input  [7:0] I_4_0_2_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_5_0_1_2,
  input  [7:0] I_5_0_2_0,
  input  [7:0] I_5_0_2_1,
  input  [7:0] I_5_0_2_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_6_0_1_2,
  input  [7:0] I_6_0_2_0,
  input  [7:0] I_6_0_2_1,
  input  [7:0] I_6_0_2_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_7_0_1_2,
  input  [7:0] I_7_0_2_0,
  input  [7:0] I_7_0_2_1,
  input  [7:0] I_7_0_2_2,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_0_2,
  input  [7:0] I_8_0_1_0,
  input  [7:0] I_8_0_1_1,
  input  [7:0] I_8_0_1_2,
  input  [7:0] I_8_0_2_0,
  input  [7:0] I_8_0_2_1,
  input  [7:0] I_8_0_2_2,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_0_2,
  input  [7:0] I_9_0_1_0,
  input  [7:0] I_9_0_1_1,
  input  [7:0] I_9_0_1_2,
  input  [7:0] I_9_0_2_0,
  input  [7:0] I_9_0_2_1,
  input  [7:0] I_9_0_2_2,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_0_2,
  input  [7:0] I_10_0_1_0,
  input  [7:0] I_10_0_1_1,
  input  [7:0] I_10_0_1_2,
  input  [7:0] I_10_0_2_0,
  input  [7:0] I_10_0_2_1,
  input  [7:0] I_10_0_2_2,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_0_2,
  input  [7:0] I_11_0_1_0,
  input  [7:0] I_11_0_1_1,
  input  [7:0] I_11_0_1_2,
  input  [7:0] I_11_0_2_0,
  input  [7:0] I_11_0_2_1,
  input  [7:0] I_11_0_2_2,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_0_2,
  input  [7:0] I_12_0_1_0,
  input  [7:0] I_12_0_1_1,
  input  [7:0] I_12_0_1_2,
  input  [7:0] I_12_0_2_0,
  input  [7:0] I_12_0_2_1,
  input  [7:0] I_12_0_2_2,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_0_2,
  input  [7:0] I_13_0_1_0,
  input  [7:0] I_13_0_1_1,
  input  [7:0] I_13_0_1_2,
  input  [7:0] I_13_0_2_0,
  input  [7:0] I_13_0_2_1,
  input  [7:0] I_13_0_2_2,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_0_2,
  input  [7:0] I_14_0_1_0,
  input  [7:0] I_14_0_1_1,
  input  [7:0] I_14_0_1_2,
  input  [7:0] I_14_0_2_0,
  input  [7:0] I_14_0_2_1,
  input  [7:0] I_14_0_2_2,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_0_2,
  input  [7:0] I_15_0_1_0,
  input  [7:0] I_15_0_1_1,
  input  [7:0] I_15_0_1_2,
  input  [7:0] I_15_0_2_0,
  input  [7:0] I_15_0_2_1,
  input  [7:0] I_15_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_8_2_0,
  output [7:0] O_8_2_1,
  output [7:0] O_8_2_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_9_2_0,
  output [7:0] O_9_2_1,
  output [7:0] O_9_2_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_10_2_0,
  output [7:0] O_10_2_1,
  output [7:0] O_10_2_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_11_2_0,
  output [7:0] O_11_2_1,
  output [7:0] O_11_2_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_12_2_0,
  output [7:0] O_12_2_1,
  output [7:0] O_12_2_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_13_2_0,
  output [7:0] O_13_2_1,
  output [7:0] O_13_2_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_14_2_0,
  output [7:0] O_14_2_1,
  output [7:0] O_14_2_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2,
  output [7:0] O_15_2_0,
  output [7:0] O_15_2_1,
  output [7:0] O_15_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_2_2; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_2_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S_3 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_0_2(fst_op_I_0_0_2),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .I_0_1_2(fst_op_I_0_1_2),
    .I_0_2_0(fst_op_I_0_2_0),
    .I_0_2_1(fst_op_I_0_2_1),
    .I_0_2_2(fst_op_I_0_2_2),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_0_2(fst_op_O_0_2),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1),
    .O_1_2(fst_op_O_1_2),
    .O_2_0(fst_op_O_2_0),
    .O_2_1(fst_op_O_2_1),
    .O_2_2(fst_op_O_2_2)
  );
  Remove1S_3 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_0_2(other_ops_0_I_0_0_2),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .I_0_1_2(other_ops_0_I_0_1_2),
    .I_0_2_0(other_ops_0_I_0_2_0),
    .I_0_2_1(other_ops_0_I_0_2_1),
    .I_0_2_2(other_ops_0_I_0_2_2),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_0_2(other_ops_0_O_0_2),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1),
    .O_1_2(other_ops_0_O_1_2),
    .O_2_0(other_ops_0_O_2_0),
    .O_2_1(other_ops_0_O_2_1),
    .O_2_2(other_ops_0_O_2_2)
  );
  Remove1S_3 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_0_2(other_ops_1_I_0_0_2),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .I_0_1_2(other_ops_1_I_0_1_2),
    .I_0_2_0(other_ops_1_I_0_2_0),
    .I_0_2_1(other_ops_1_I_0_2_1),
    .I_0_2_2(other_ops_1_I_0_2_2),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_0_2(other_ops_1_O_0_2),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1),
    .O_1_2(other_ops_1_O_1_2),
    .O_2_0(other_ops_1_O_2_0),
    .O_2_1(other_ops_1_O_2_1),
    .O_2_2(other_ops_1_O_2_2)
  );
  Remove1S_3 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_0_2(other_ops_2_I_0_0_2),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .I_0_1_2(other_ops_2_I_0_1_2),
    .I_0_2_0(other_ops_2_I_0_2_0),
    .I_0_2_1(other_ops_2_I_0_2_1),
    .I_0_2_2(other_ops_2_I_0_2_2),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_0_2(other_ops_2_O_0_2),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1),
    .O_1_2(other_ops_2_O_1_2),
    .O_2_0(other_ops_2_O_2_0),
    .O_2_1(other_ops_2_O_2_1),
    .O_2_2(other_ops_2_O_2_2)
  );
  Remove1S_3 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_0_2(other_ops_3_I_0_0_2),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .I_0_1_2(other_ops_3_I_0_1_2),
    .I_0_2_0(other_ops_3_I_0_2_0),
    .I_0_2_1(other_ops_3_I_0_2_1),
    .I_0_2_2(other_ops_3_I_0_2_2),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_0_2(other_ops_3_O_0_2),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1),
    .O_1_2(other_ops_3_O_1_2),
    .O_2_0(other_ops_3_O_2_0),
    .O_2_1(other_ops_3_O_2_1),
    .O_2_2(other_ops_3_O_2_2)
  );
  Remove1S_3 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_0_2(other_ops_4_I_0_0_2),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .I_0_1_2(other_ops_4_I_0_1_2),
    .I_0_2_0(other_ops_4_I_0_2_0),
    .I_0_2_1(other_ops_4_I_0_2_1),
    .I_0_2_2(other_ops_4_I_0_2_2),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_0_2(other_ops_4_O_0_2),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1),
    .O_1_2(other_ops_4_O_1_2),
    .O_2_0(other_ops_4_O_2_0),
    .O_2_1(other_ops_4_O_2_1),
    .O_2_2(other_ops_4_O_2_2)
  );
  Remove1S_3 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_0_2(other_ops_5_I_0_0_2),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .I_0_1_2(other_ops_5_I_0_1_2),
    .I_0_2_0(other_ops_5_I_0_2_0),
    .I_0_2_1(other_ops_5_I_0_2_1),
    .I_0_2_2(other_ops_5_I_0_2_2),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_0_2(other_ops_5_O_0_2),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1),
    .O_1_2(other_ops_5_O_1_2),
    .O_2_0(other_ops_5_O_2_0),
    .O_2_1(other_ops_5_O_2_1),
    .O_2_2(other_ops_5_O_2_2)
  );
  Remove1S_3 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_0_2(other_ops_6_I_0_0_2),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .I_0_1_2(other_ops_6_I_0_1_2),
    .I_0_2_0(other_ops_6_I_0_2_0),
    .I_0_2_1(other_ops_6_I_0_2_1),
    .I_0_2_2(other_ops_6_I_0_2_2),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_0_2(other_ops_6_O_0_2),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1),
    .O_1_2(other_ops_6_O_1_2),
    .O_2_0(other_ops_6_O_2_0),
    .O_2_1(other_ops_6_O_2_1),
    .O_2_2(other_ops_6_O_2_2)
  );
  Remove1S_3 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0_0(other_ops_7_I_0_0_0),
    .I_0_0_1(other_ops_7_I_0_0_1),
    .I_0_0_2(other_ops_7_I_0_0_2),
    .I_0_1_0(other_ops_7_I_0_1_0),
    .I_0_1_1(other_ops_7_I_0_1_1),
    .I_0_1_2(other_ops_7_I_0_1_2),
    .I_0_2_0(other_ops_7_I_0_2_0),
    .I_0_2_1(other_ops_7_I_0_2_1),
    .I_0_2_2(other_ops_7_I_0_2_2),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_0_2(other_ops_7_O_0_2),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1),
    .O_1_2(other_ops_7_O_1_2),
    .O_2_0(other_ops_7_O_2_0),
    .O_2_1(other_ops_7_O_2_1),
    .O_2_2(other_ops_7_O_2_2)
  );
  Remove1S_3 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0_0(other_ops_8_I_0_0_0),
    .I_0_0_1(other_ops_8_I_0_0_1),
    .I_0_0_2(other_ops_8_I_0_0_2),
    .I_0_1_0(other_ops_8_I_0_1_0),
    .I_0_1_1(other_ops_8_I_0_1_1),
    .I_0_1_2(other_ops_8_I_0_1_2),
    .I_0_2_0(other_ops_8_I_0_2_0),
    .I_0_2_1(other_ops_8_I_0_2_1),
    .I_0_2_2(other_ops_8_I_0_2_2),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_0_2(other_ops_8_O_0_2),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1),
    .O_1_2(other_ops_8_O_1_2),
    .O_2_0(other_ops_8_O_2_0),
    .O_2_1(other_ops_8_O_2_1),
    .O_2_2(other_ops_8_O_2_2)
  );
  Remove1S_3 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0_0(other_ops_9_I_0_0_0),
    .I_0_0_1(other_ops_9_I_0_0_1),
    .I_0_0_2(other_ops_9_I_0_0_2),
    .I_0_1_0(other_ops_9_I_0_1_0),
    .I_0_1_1(other_ops_9_I_0_1_1),
    .I_0_1_2(other_ops_9_I_0_1_2),
    .I_0_2_0(other_ops_9_I_0_2_0),
    .I_0_2_1(other_ops_9_I_0_2_1),
    .I_0_2_2(other_ops_9_I_0_2_2),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_0_2(other_ops_9_O_0_2),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1),
    .O_1_2(other_ops_9_O_1_2),
    .O_2_0(other_ops_9_O_2_0),
    .O_2_1(other_ops_9_O_2_1),
    .O_2_2(other_ops_9_O_2_2)
  );
  Remove1S_3 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0_0(other_ops_10_I_0_0_0),
    .I_0_0_1(other_ops_10_I_0_0_1),
    .I_0_0_2(other_ops_10_I_0_0_2),
    .I_0_1_0(other_ops_10_I_0_1_0),
    .I_0_1_1(other_ops_10_I_0_1_1),
    .I_0_1_2(other_ops_10_I_0_1_2),
    .I_0_2_0(other_ops_10_I_0_2_0),
    .I_0_2_1(other_ops_10_I_0_2_1),
    .I_0_2_2(other_ops_10_I_0_2_2),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_0_2(other_ops_10_O_0_2),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1),
    .O_1_2(other_ops_10_O_1_2),
    .O_2_0(other_ops_10_O_2_0),
    .O_2_1(other_ops_10_O_2_1),
    .O_2_2(other_ops_10_O_2_2)
  );
  Remove1S_3 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0_0(other_ops_11_I_0_0_0),
    .I_0_0_1(other_ops_11_I_0_0_1),
    .I_0_0_2(other_ops_11_I_0_0_2),
    .I_0_1_0(other_ops_11_I_0_1_0),
    .I_0_1_1(other_ops_11_I_0_1_1),
    .I_0_1_2(other_ops_11_I_0_1_2),
    .I_0_2_0(other_ops_11_I_0_2_0),
    .I_0_2_1(other_ops_11_I_0_2_1),
    .I_0_2_2(other_ops_11_I_0_2_2),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_0_2(other_ops_11_O_0_2),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1),
    .O_1_2(other_ops_11_O_1_2),
    .O_2_0(other_ops_11_O_2_0),
    .O_2_1(other_ops_11_O_2_1),
    .O_2_2(other_ops_11_O_2_2)
  );
  Remove1S_3 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0_0(other_ops_12_I_0_0_0),
    .I_0_0_1(other_ops_12_I_0_0_1),
    .I_0_0_2(other_ops_12_I_0_0_2),
    .I_0_1_0(other_ops_12_I_0_1_0),
    .I_0_1_1(other_ops_12_I_0_1_1),
    .I_0_1_2(other_ops_12_I_0_1_2),
    .I_0_2_0(other_ops_12_I_0_2_0),
    .I_0_2_1(other_ops_12_I_0_2_1),
    .I_0_2_2(other_ops_12_I_0_2_2),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_0_2(other_ops_12_O_0_2),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1),
    .O_1_2(other_ops_12_O_1_2),
    .O_2_0(other_ops_12_O_2_0),
    .O_2_1(other_ops_12_O_2_1),
    .O_2_2(other_ops_12_O_2_2)
  );
  Remove1S_3 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0_0(other_ops_13_I_0_0_0),
    .I_0_0_1(other_ops_13_I_0_0_1),
    .I_0_0_2(other_ops_13_I_0_0_2),
    .I_0_1_0(other_ops_13_I_0_1_0),
    .I_0_1_1(other_ops_13_I_0_1_1),
    .I_0_1_2(other_ops_13_I_0_1_2),
    .I_0_2_0(other_ops_13_I_0_2_0),
    .I_0_2_1(other_ops_13_I_0_2_1),
    .I_0_2_2(other_ops_13_I_0_2_2),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_0_2(other_ops_13_O_0_2),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1),
    .O_1_2(other_ops_13_O_1_2),
    .O_2_0(other_ops_13_O_2_0),
    .O_2_1(other_ops_13_O_2_1),
    .O_2_2(other_ops_13_O_2_2)
  );
  Remove1S_3 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0_0(other_ops_14_I_0_0_0),
    .I_0_0_1(other_ops_14_I_0_0_1),
    .I_0_0_2(other_ops_14_I_0_0_2),
    .I_0_1_0(other_ops_14_I_0_1_0),
    .I_0_1_1(other_ops_14_I_0_1_1),
    .I_0_1_2(other_ops_14_I_0_1_2),
    .I_0_2_0(other_ops_14_I_0_2_0),
    .I_0_2_1(other_ops_14_I_0_2_1),
    .I_0_2_2(other_ops_14_I_0_2_2),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_0_2(other_ops_14_O_0_2),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1),
    .O_1_2(other_ops_14_O_1_2),
    .O_2_0(other_ops_14_O_2_0),
    .O_2_1(other_ops_14_O_2_1),
    .O_2_2(other_ops_14_O_2_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_0_2 = fst_op_O_0_2; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_0_1_2 = fst_op_O_1_2; // @[MapS.scala 17:8]
  assign O_0_2_0 = fst_op_O_2_0; // @[MapS.scala 17:8]
  assign O_0_2_1 = fst_op_O_2_1; // @[MapS.scala 17:8]
  assign O_0_2_2 = fst_op_O_2_2; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_0_2 = other_ops_0_O_0_2; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_1_1_2 = other_ops_0_O_1_2; // @[MapS.scala 21:12]
  assign O_1_2_0 = other_ops_0_O_2_0; // @[MapS.scala 21:12]
  assign O_1_2_1 = other_ops_0_O_2_1; // @[MapS.scala 21:12]
  assign O_1_2_2 = other_ops_0_O_2_2; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_0_2 = other_ops_1_O_0_2; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_2_1_2 = other_ops_1_O_1_2; // @[MapS.scala 21:12]
  assign O_2_2_0 = other_ops_1_O_2_0; // @[MapS.scala 21:12]
  assign O_2_2_1 = other_ops_1_O_2_1; // @[MapS.scala 21:12]
  assign O_2_2_2 = other_ops_1_O_2_2; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_0_2 = other_ops_2_O_0_2; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_3_1_2 = other_ops_2_O_1_2; // @[MapS.scala 21:12]
  assign O_3_2_0 = other_ops_2_O_2_0; // @[MapS.scala 21:12]
  assign O_3_2_1 = other_ops_2_O_2_1; // @[MapS.scala 21:12]
  assign O_3_2_2 = other_ops_2_O_2_2; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_0_2 = other_ops_3_O_0_2; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_4_1_2 = other_ops_3_O_1_2; // @[MapS.scala 21:12]
  assign O_4_2_0 = other_ops_3_O_2_0; // @[MapS.scala 21:12]
  assign O_4_2_1 = other_ops_3_O_2_1; // @[MapS.scala 21:12]
  assign O_4_2_2 = other_ops_3_O_2_2; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_0_2 = other_ops_4_O_0_2; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_5_1_2 = other_ops_4_O_1_2; // @[MapS.scala 21:12]
  assign O_5_2_0 = other_ops_4_O_2_0; // @[MapS.scala 21:12]
  assign O_5_2_1 = other_ops_4_O_2_1; // @[MapS.scala 21:12]
  assign O_5_2_2 = other_ops_4_O_2_2; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_0_2 = other_ops_5_O_0_2; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_6_1_2 = other_ops_5_O_1_2; // @[MapS.scala 21:12]
  assign O_6_2_0 = other_ops_5_O_2_0; // @[MapS.scala 21:12]
  assign O_6_2_1 = other_ops_5_O_2_1; // @[MapS.scala 21:12]
  assign O_6_2_2 = other_ops_5_O_2_2; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_0_2 = other_ops_6_O_0_2; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_7_1_2 = other_ops_6_O_1_2; // @[MapS.scala 21:12]
  assign O_7_2_0 = other_ops_6_O_2_0; // @[MapS.scala 21:12]
  assign O_7_2_1 = other_ops_6_O_2_1; // @[MapS.scala 21:12]
  assign O_7_2_2 = other_ops_6_O_2_2; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[MapS.scala 21:12]
  assign O_8_0_2 = other_ops_7_O_0_2; // @[MapS.scala 21:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[MapS.scala 21:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[MapS.scala 21:12]
  assign O_8_1_2 = other_ops_7_O_1_2; // @[MapS.scala 21:12]
  assign O_8_2_0 = other_ops_7_O_2_0; // @[MapS.scala 21:12]
  assign O_8_2_1 = other_ops_7_O_2_1; // @[MapS.scala 21:12]
  assign O_8_2_2 = other_ops_7_O_2_2; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[MapS.scala 21:12]
  assign O_9_0_2 = other_ops_8_O_0_2; // @[MapS.scala 21:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[MapS.scala 21:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[MapS.scala 21:12]
  assign O_9_1_2 = other_ops_8_O_1_2; // @[MapS.scala 21:12]
  assign O_9_2_0 = other_ops_8_O_2_0; // @[MapS.scala 21:12]
  assign O_9_2_1 = other_ops_8_O_2_1; // @[MapS.scala 21:12]
  assign O_9_2_2 = other_ops_8_O_2_2; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[MapS.scala 21:12]
  assign O_10_0_2 = other_ops_9_O_0_2; // @[MapS.scala 21:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[MapS.scala 21:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[MapS.scala 21:12]
  assign O_10_1_2 = other_ops_9_O_1_2; // @[MapS.scala 21:12]
  assign O_10_2_0 = other_ops_9_O_2_0; // @[MapS.scala 21:12]
  assign O_10_2_1 = other_ops_9_O_2_1; // @[MapS.scala 21:12]
  assign O_10_2_2 = other_ops_9_O_2_2; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[MapS.scala 21:12]
  assign O_11_0_2 = other_ops_10_O_0_2; // @[MapS.scala 21:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[MapS.scala 21:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[MapS.scala 21:12]
  assign O_11_1_2 = other_ops_10_O_1_2; // @[MapS.scala 21:12]
  assign O_11_2_0 = other_ops_10_O_2_0; // @[MapS.scala 21:12]
  assign O_11_2_1 = other_ops_10_O_2_1; // @[MapS.scala 21:12]
  assign O_11_2_2 = other_ops_10_O_2_2; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[MapS.scala 21:12]
  assign O_12_0_2 = other_ops_11_O_0_2; // @[MapS.scala 21:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[MapS.scala 21:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[MapS.scala 21:12]
  assign O_12_1_2 = other_ops_11_O_1_2; // @[MapS.scala 21:12]
  assign O_12_2_0 = other_ops_11_O_2_0; // @[MapS.scala 21:12]
  assign O_12_2_1 = other_ops_11_O_2_1; // @[MapS.scala 21:12]
  assign O_12_2_2 = other_ops_11_O_2_2; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[MapS.scala 21:12]
  assign O_13_0_2 = other_ops_12_O_0_2; // @[MapS.scala 21:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[MapS.scala 21:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[MapS.scala 21:12]
  assign O_13_1_2 = other_ops_12_O_1_2; // @[MapS.scala 21:12]
  assign O_13_2_0 = other_ops_12_O_2_0; // @[MapS.scala 21:12]
  assign O_13_2_1 = other_ops_12_O_2_1; // @[MapS.scala 21:12]
  assign O_13_2_2 = other_ops_12_O_2_2; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[MapS.scala 21:12]
  assign O_14_0_2 = other_ops_13_O_0_2; // @[MapS.scala 21:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[MapS.scala 21:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[MapS.scala 21:12]
  assign O_14_1_2 = other_ops_13_O_1_2; // @[MapS.scala 21:12]
  assign O_14_2_0 = other_ops_13_O_2_0; // @[MapS.scala 21:12]
  assign O_14_2_1 = other_ops_13_O_2_1; // @[MapS.scala 21:12]
  assign O_14_2_2 = other_ops_13_O_2_2; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[MapS.scala 21:12]
  assign O_15_0_2 = other_ops_14_O_0_2; // @[MapS.scala 21:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[MapS.scala 21:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[MapS.scala 21:12]
  assign O_15_1_2 = other_ops_14_O_1_2; // @[MapS.scala 21:12]
  assign O_15_2_0 = other_ops_14_O_2_0; // @[MapS.scala 21:12]
  assign O_15_2_1 = other_ops_14_O_2_1; // @[MapS.scala 21:12]
  assign O_15_2_2 = other_ops_14_O_2_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_2 = I_0_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_2 = I_0_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_0 = I_0_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_1 = I_0_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2_2 = I_0_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_2 = I_1_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_2 = I_1_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_0 = I_1_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_1 = I_1_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2_2 = I_1_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_2 = I_2_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_2 = I_2_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_0 = I_2_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_1 = I_2_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2_2 = I_2_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_2 = I_3_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_2 = I_3_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_0 = I_3_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_1 = I_3_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2_2 = I_3_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_2 = I_4_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_2 = I_4_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_0 = I_4_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_1 = I_4_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2_2 = I_4_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_2 = I_5_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_2 = I_5_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_0 = I_5_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_1 = I_5_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2_2 = I_5_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_2 = I_6_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_2 = I_6_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_0 = I_6_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_1 = I_6_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2_2 = I_6_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_2 = I_7_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_2 = I_7_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_0 = I_7_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_1 = I_7_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2_2 = I_7_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0_0 = I_8_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_1 = I_8_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_2 = I_8_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_0 = I_8_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_1 = I_8_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_2 = I_8_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_0 = I_8_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_1 = I_8_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2_2 = I_8_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0_0 = I_9_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_1 = I_9_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_2 = I_9_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_0 = I_9_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_1 = I_9_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_2 = I_9_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_0 = I_9_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_1 = I_9_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2_2 = I_9_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0_0 = I_10_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_1 = I_10_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_2 = I_10_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_0 = I_10_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_1 = I_10_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_2 = I_10_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_0 = I_10_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_1 = I_10_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2_2 = I_10_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0_0 = I_11_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_1 = I_11_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_2 = I_11_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_0 = I_11_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_1 = I_11_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_2 = I_11_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_0 = I_11_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_1 = I_11_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2_2 = I_11_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0_0 = I_12_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_1 = I_12_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_2 = I_12_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_0 = I_12_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_1 = I_12_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_2 = I_12_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_0 = I_12_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_1 = I_12_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2_2 = I_12_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0_0 = I_13_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_1 = I_13_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_2 = I_13_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_0 = I_13_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_1 = I_13_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_2 = I_13_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_0 = I_13_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_1 = I_13_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2_2 = I_13_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0_0 = I_14_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_1 = I_14_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_2 = I_14_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_0 = I_14_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_1 = I_14_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_2 = I_14_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_0 = I_14_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_1 = I_14_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2_2 = I_14_0_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0_0 = I_15_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_1 = I_15_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_2 = I_15_0_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_0 = I_15_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_1 = I_15_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_2 = I_15_0_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_0 = I_15_0_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_1 = I_15_0_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2_2 = I_15_0_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_0_2,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_0_0_1_2,
  input  [7:0] I_0_0_2_0,
  input  [7:0] I_0_0_2_1,
  input  [7:0] I_0_0_2_2,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_0_2,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_1_0_1_2,
  input  [7:0] I_1_0_2_0,
  input  [7:0] I_1_0_2_1,
  input  [7:0] I_1_0_2_2,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_0_2,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_2_0_1_2,
  input  [7:0] I_2_0_2_0,
  input  [7:0] I_2_0_2_1,
  input  [7:0] I_2_0_2_2,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_0_2,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_3_0_1_2,
  input  [7:0] I_3_0_2_0,
  input  [7:0] I_3_0_2_1,
  input  [7:0] I_3_0_2_2,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_0_2,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_4_0_1_2,
  input  [7:0] I_4_0_2_0,
  input  [7:0] I_4_0_2_1,
  input  [7:0] I_4_0_2_2,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_0_2,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_5_0_1_2,
  input  [7:0] I_5_0_2_0,
  input  [7:0] I_5_0_2_1,
  input  [7:0] I_5_0_2_2,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_0_2,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_6_0_1_2,
  input  [7:0] I_6_0_2_0,
  input  [7:0] I_6_0_2_1,
  input  [7:0] I_6_0_2_2,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_0_2,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_7_0_1_2,
  input  [7:0] I_7_0_2_0,
  input  [7:0] I_7_0_2_1,
  input  [7:0] I_7_0_2_2,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_0_2,
  input  [7:0] I_8_0_1_0,
  input  [7:0] I_8_0_1_1,
  input  [7:0] I_8_0_1_2,
  input  [7:0] I_8_0_2_0,
  input  [7:0] I_8_0_2_1,
  input  [7:0] I_8_0_2_2,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_0_2,
  input  [7:0] I_9_0_1_0,
  input  [7:0] I_9_0_1_1,
  input  [7:0] I_9_0_1_2,
  input  [7:0] I_9_0_2_0,
  input  [7:0] I_9_0_2_1,
  input  [7:0] I_9_0_2_2,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_0_2,
  input  [7:0] I_10_0_1_0,
  input  [7:0] I_10_0_1_1,
  input  [7:0] I_10_0_1_2,
  input  [7:0] I_10_0_2_0,
  input  [7:0] I_10_0_2_1,
  input  [7:0] I_10_0_2_2,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_0_2,
  input  [7:0] I_11_0_1_0,
  input  [7:0] I_11_0_1_1,
  input  [7:0] I_11_0_1_2,
  input  [7:0] I_11_0_2_0,
  input  [7:0] I_11_0_2_1,
  input  [7:0] I_11_0_2_2,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_0_2,
  input  [7:0] I_12_0_1_0,
  input  [7:0] I_12_0_1_1,
  input  [7:0] I_12_0_1_2,
  input  [7:0] I_12_0_2_0,
  input  [7:0] I_12_0_2_1,
  input  [7:0] I_12_0_2_2,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_0_2,
  input  [7:0] I_13_0_1_0,
  input  [7:0] I_13_0_1_1,
  input  [7:0] I_13_0_1_2,
  input  [7:0] I_13_0_2_0,
  input  [7:0] I_13_0_2_1,
  input  [7:0] I_13_0_2_2,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_0_2,
  input  [7:0] I_14_0_1_0,
  input  [7:0] I_14_0_1_1,
  input  [7:0] I_14_0_1_2,
  input  [7:0] I_14_0_2_0,
  input  [7:0] I_14_0_2_1,
  input  [7:0] I_14_0_2_2,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_0_2,
  input  [7:0] I_15_0_1_0,
  input  [7:0] I_15_0_1_1,
  input  [7:0] I_15_0_1_2,
  input  [7:0] I_15_0_2_0,
  input  [7:0] I_15_0_2_1,
  input  [7:0] I_15_0_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_0_2,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_0_1_2,
  output [7:0] O_0_2_0,
  output [7:0] O_0_2_1,
  output [7:0] O_0_2_2,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_0_2,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_1_1_2,
  output [7:0] O_1_2_0,
  output [7:0] O_1_2_1,
  output [7:0] O_1_2_2,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_0_2,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_2_1_2,
  output [7:0] O_2_2_0,
  output [7:0] O_2_2_1,
  output [7:0] O_2_2_2,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_0_2,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_3_1_2,
  output [7:0] O_3_2_0,
  output [7:0] O_3_2_1,
  output [7:0] O_3_2_2,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_0_2,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_4_1_2,
  output [7:0] O_4_2_0,
  output [7:0] O_4_2_1,
  output [7:0] O_4_2_2,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_0_2,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_5_1_2,
  output [7:0] O_5_2_0,
  output [7:0] O_5_2_1,
  output [7:0] O_5_2_2,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_0_2,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_6_1_2,
  output [7:0] O_6_2_0,
  output [7:0] O_6_2_1,
  output [7:0] O_6_2_2,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_0_2,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_7_1_2,
  output [7:0] O_7_2_0,
  output [7:0] O_7_2_1,
  output [7:0] O_7_2_2,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_0_2,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_8_1_2,
  output [7:0] O_8_2_0,
  output [7:0] O_8_2_1,
  output [7:0] O_8_2_2,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_0_2,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_9_1_2,
  output [7:0] O_9_2_0,
  output [7:0] O_9_2_1,
  output [7:0] O_9_2_2,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_0_2,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_10_1_2,
  output [7:0] O_10_2_0,
  output [7:0] O_10_2_1,
  output [7:0] O_10_2_2,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_0_2,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_11_1_2,
  output [7:0] O_11_2_0,
  output [7:0] O_11_2_1,
  output [7:0] O_11_2_2,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_0_2,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_12_1_2,
  output [7:0] O_12_2_0,
  output [7:0] O_12_2_1,
  output [7:0] O_12_2_2,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_0_2,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_13_1_2,
  output [7:0] O_13_2_0,
  output [7:0] O_13_2_1,
  output [7:0] O_13_2_2,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_0_2,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_14_1_2,
  output [7:0] O_14_2_0,
  output [7:0] O_14_2_1,
  output [7:0] O_14_2_2,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_0_2,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1,
  output [7:0] O_15_1_2,
  output [7:0] O_15_2_0,
  output [7:0] O_15_2_1,
  output [7:0] O_15_2_2
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_2_2; // @[MapT.scala 8:20]
  MapS_3 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_0_2(op_I_0_0_0_2),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_0_0_1_2(op_I_0_0_1_2),
    .I_0_0_2_0(op_I_0_0_2_0),
    .I_0_0_2_1(op_I_0_0_2_1),
    .I_0_0_2_2(op_I_0_0_2_2),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_0_2(op_I_1_0_0_2),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_1_0_1_2(op_I_1_0_1_2),
    .I_1_0_2_0(op_I_1_0_2_0),
    .I_1_0_2_1(op_I_1_0_2_1),
    .I_1_0_2_2(op_I_1_0_2_2),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_0_2(op_I_2_0_0_2),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_2_0_1_2(op_I_2_0_1_2),
    .I_2_0_2_0(op_I_2_0_2_0),
    .I_2_0_2_1(op_I_2_0_2_1),
    .I_2_0_2_2(op_I_2_0_2_2),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_0_2(op_I_3_0_0_2),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_3_0_1_2(op_I_3_0_1_2),
    .I_3_0_2_0(op_I_3_0_2_0),
    .I_3_0_2_1(op_I_3_0_2_1),
    .I_3_0_2_2(op_I_3_0_2_2),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_0_2(op_I_4_0_0_2),
    .I_4_0_1_0(op_I_4_0_1_0),
    .I_4_0_1_1(op_I_4_0_1_1),
    .I_4_0_1_2(op_I_4_0_1_2),
    .I_4_0_2_0(op_I_4_0_2_0),
    .I_4_0_2_1(op_I_4_0_2_1),
    .I_4_0_2_2(op_I_4_0_2_2),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_0_2(op_I_5_0_0_2),
    .I_5_0_1_0(op_I_5_0_1_0),
    .I_5_0_1_1(op_I_5_0_1_1),
    .I_5_0_1_2(op_I_5_0_1_2),
    .I_5_0_2_0(op_I_5_0_2_0),
    .I_5_0_2_1(op_I_5_0_2_1),
    .I_5_0_2_2(op_I_5_0_2_2),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_0_2(op_I_6_0_0_2),
    .I_6_0_1_0(op_I_6_0_1_0),
    .I_6_0_1_1(op_I_6_0_1_1),
    .I_6_0_1_2(op_I_6_0_1_2),
    .I_6_0_2_0(op_I_6_0_2_0),
    .I_6_0_2_1(op_I_6_0_2_1),
    .I_6_0_2_2(op_I_6_0_2_2),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_0_2(op_I_7_0_0_2),
    .I_7_0_1_0(op_I_7_0_1_0),
    .I_7_0_1_1(op_I_7_0_1_1),
    .I_7_0_1_2(op_I_7_0_1_2),
    .I_7_0_2_0(op_I_7_0_2_0),
    .I_7_0_2_1(op_I_7_0_2_1),
    .I_7_0_2_2(op_I_7_0_2_2),
    .I_8_0_0_0(op_I_8_0_0_0),
    .I_8_0_0_1(op_I_8_0_0_1),
    .I_8_0_0_2(op_I_8_0_0_2),
    .I_8_0_1_0(op_I_8_0_1_0),
    .I_8_0_1_1(op_I_8_0_1_1),
    .I_8_0_1_2(op_I_8_0_1_2),
    .I_8_0_2_0(op_I_8_0_2_0),
    .I_8_0_2_1(op_I_8_0_2_1),
    .I_8_0_2_2(op_I_8_0_2_2),
    .I_9_0_0_0(op_I_9_0_0_0),
    .I_9_0_0_1(op_I_9_0_0_1),
    .I_9_0_0_2(op_I_9_0_0_2),
    .I_9_0_1_0(op_I_9_0_1_0),
    .I_9_0_1_1(op_I_9_0_1_1),
    .I_9_0_1_2(op_I_9_0_1_2),
    .I_9_0_2_0(op_I_9_0_2_0),
    .I_9_0_2_1(op_I_9_0_2_1),
    .I_9_0_2_2(op_I_9_0_2_2),
    .I_10_0_0_0(op_I_10_0_0_0),
    .I_10_0_0_1(op_I_10_0_0_1),
    .I_10_0_0_2(op_I_10_0_0_2),
    .I_10_0_1_0(op_I_10_0_1_0),
    .I_10_0_1_1(op_I_10_0_1_1),
    .I_10_0_1_2(op_I_10_0_1_2),
    .I_10_0_2_0(op_I_10_0_2_0),
    .I_10_0_2_1(op_I_10_0_2_1),
    .I_10_0_2_2(op_I_10_0_2_2),
    .I_11_0_0_0(op_I_11_0_0_0),
    .I_11_0_0_1(op_I_11_0_0_1),
    .I_11_0_0_2(op_I_11_0_0_2),
    .I_11_0_1_0(op_I_11_0_1_0),
    .I_11_0_1_1(op_I_11_0_1_1),
    .I_11_0_1_2(op_I_11_0_1_2),
    .I_11_0_2_0(op_I_11_0_2_0),
    .I_11_0_2_1(op_I_11_0_2_1),
    .I_11_0_2_2(op_I_11_0_2_2),
    .I_12_0_0_0(op_I_12_0_0_0),
    .I_12_0_0_1(op_I_12_0_0_1),
    .I_12_0_0_2(op_I_12_0_0_2),
    .I_12_0_1_0(op_I_12_0_1_0),
    .I_12_0_1_1(op_I_12_0_1_1),
    .I_12_0_1_2(op_I_12_0_1_2),
    .I_12_0_2_0(op_I_12_0_2_0),
    .I_12_0_2_1(op_I_12_0_2_1),
    .I_12_0_2_2(op_I_12_0_2_2),
    .I_13_0_0_0(op_I_13_0_0_0),
    .I_13_0_0_1(op_I_13_0_0_1),
    .I_13_0_0_2(op_I_13_0_0_2),
    .I_13_0_1_0(op_I_13_0_1_0),
    .I_13_0_1_1(op_I_13_0_1_1),
    .I_13_0_1_2(op_I_13_0_1_2),
    .I_13_0_2_0(op_I_13_0_2_0),
    .I_13_0_2_1(op_I_13_0_2_1),
    .I_13_0_2_2(op_I_13_0_2_2),
    .I_14_0_0_0(op_I_14_0_0_0),
    .I_14_0_0_1(op_I_14_0_0_1),
    .I_14_0_0_2(op_I_14_0_0_2),
    .I_14_0_1_0(op_I_14_0_1_0),
    .I_14_0_1_1(op_I_14_0_1_1),
    .I_14_0_1_2(op_I_14_0_1_2),
    .I_14_0_2_0(op_I_14_0_2_0),
    .I_14_0_2_1(op_I_14_0_2_1),
    .I_14_0_2_2(op_I_14_0_2_2),
    .I_15_0_0_0(op_I_15_0_0_0),
    .I_15_0_0_1(op_I_15_0_0_1),
    .I_15_0_0_2(op_I_15_0_0_2),
    .I_15_0_1_0(op_I_15_0_1_0),
    .I_15_0_1_1(op_I_15_0_1_1),
    .I_15_0_1_2(op_I_15_0_1_2),
    .I_15_0_2_0(op_I_15_0_2_0),
    .I_15_0_2_1(op_I_15_0_2_1),
    .I_15_0_2_2(op_I_15_0_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_0_2(op_O_0_0_2),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_0_1_2(op_O_0_1_2),
    .O_0_2_0(op_O_0_2_0),
    .O_0_2_1(op_O_0_2_1),
    .O_0_2_2(op_O_0_2_2),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_0_2(op_O_1_0_2),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_1_1_2(op_O_1_1_2),
    .O_1_2_0(op_O_1_2_0),
    .O_1_2_1(op_O_1_2_1),
    .O_1_2_2(op_O_1_2_2),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_0_2(op_O_2_0_2),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_2_1_2(op_O_2_1_2),
    .O_2_2_0(op_O_2_2_0),
    .O_2_2_1(op_O_2_2_1),
    .O_2_2_2(op_O_2_2_2),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_0_2(op_O_3_0_2),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_3_1_2(op_O_3_1_2),
    .O_3_2_0(op_O_3_2_0),
    .O_3_2_1(op_O_3_2_1),
    .O_3_2_2(op_O_3_2_2),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_0_2(op_O_4_0_2),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_4_1_2(op_O_4_1_2),
    .O_4_2_0(op_O_4_2_0),
    .O_4_2_1(op_O_4_2_1),
    .O_4_2_2(op_O_4_2_2),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_0_2(op_O_5_0_2),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_5_1_2(op_O_5_1_2),
    .O_5_2_0(op_O_5_2_0),
    .O_5_2_1(op_O_5_2_1),
    .O_5_2_2(op_O_5_2_2),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_0_2(op_O_6_0_2),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_6_1_2(op_O_6_1_2),
    .O_6_2_0(op_O_6_2_0),
    .O_6_2_1(op_O_6_2_1),
    .O_6_2_2(op_O_6_2_2),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_0_2(op_O_7_0_2),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_7_1_2(op_O_7_1_2),
    .O_7_2_0(op_O_7_2_0),
    .O_7_2_1(op_O_7_2_1),
    .O_7_2_2(op_O_7_2_2),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_0_2(op_O_8_0_2),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_8_1_2(op_O_8_1_2),
    .O_8_2_0(op_O_8_2_0),
    .O_8_2_1(op_O_8_2_1),
    .O_8_2_2(op_O_8_2_2),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_0_2(op_O_9_0_2),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_9_1_2(op_O_9_1_2),
    .O_9_2_0(op_O_9_2_0),
    .O_9_2_1(op_O_9_2_1),
    .O_9_2_2(op_O_9_2_2),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_0_2(op_O_10_0_2),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_10_1_2(op_O_10_1_2),
    .O_10_2_0(op_O_10_2_0),
    .O_10_2_1(op_O_10_2_1),
    .O_10_2_2(op_O_10_2_2),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_0_2(op_O_11_0_2),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_11_1_2(op_O_11_1_2),
    .O_11_2_0(op_O_11_2_0),
    .O_11_2_1(op_O_11_2_1),
    .O_11_2_2(op_O_11_2_2),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_0_2(op_O_12_0_2),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_12_1_2(op_O_12_1_2),
    .O_12_2_0(op_O_12_2_0),
    .O_12_2_1(op_O_12_2_1),
    .O_12_2_2(op_O_12_2_2),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_0_2(op_O_13_0_2),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_13_1_2(op_O_13_1_2),
    .O_13_2_0(op_O_13_2_0),
    .O_13_2_1(op_O_13_2_1),
    .O_13_2_2(op_O_13_2_2),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_0_2(op_O_14_0_2),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_14_1_2(op_O_14_1_2),
    .O_14_2_0(op_O_14_2_0),
    .O_14_2_1(op_O_14_2_1),
    .O_14_2_2(op_O_14_2_2),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_0_2(op_O_15_0_2),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1),
    .O_15_1_2(op_O_15_1_2),
    .O_15_2_0(op_O_15_2_0),
    .O_15_2_1(op_O_15_2_1),
    .O_15_2_2(op_O_15_2_2)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_2 = op_O_0_0_2; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_0_1_2 = op_O_0_1_2; // @[MapT.scala 15:7]
  assign O_0_2_0 = op_O_0_2_0; // @[MapT.scala 15:7]
  assign O_0_2_1 = op_O_0_2_1; // @[MapT.scala 15:7]
  assign O_0_2_2 = op_O_0_2_2; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_0_2 = op_O_1_0_2; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_1_1_2 = op_O_1_1_2; // @[MapT.scala 15:7]
  assign O_1_2_0 = op_O_1_2_0; // @[MapT.scala 15:7]
  assign O_1_2_1 = op_O_1_2_1; // @[MapT.scala 15:7]
  assign O_1_2_2 = op_O_1_2_2; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_0_2 = op_O_2_0_2; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_2_1_2 = op_O_2_1_2; // @[MapT.scala 15:7]
  assign O_2_2_0 = op_O_2_2_0; // @[MapT.scala 15:7]
  assign O_2_2_1 = op_O_2_2_1; // @[MapT.scala 15:7]
  assign O_2_2_2 = op_O_2_2_2; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_0_2 = op_O_3_0_2; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_3_1_2 = op_O_3_1_2; // @[MapT.scala 15:7]
  assign O_3_2_0 = op_O_3_2_0; // @[MapT.scala 15:7]
  assign O_3_2_1 = op_O_3_2_1; // @[MapT.scala 15:7]
  assign O_3_2_2 = op_O_3_2_2; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_0_2 = op_O_4_0_2; // @[MapT.scala 15:7]
  assign O_4_1_0 = op_O_4_1_0; // @[MapT.scala 15:7]
  assign O_4_1_1 = op_O_4_1_1; // @[MapT.scala 15:7]
  assign O_4_1_2 = op_O_4_1_2; // @[MapT.scala 15:7]
  assign O_4_2_0 = op_O_4_2_0; // @[MapT.scala 15:7]
  assign O_4_2_1 = op_O_4_2_1; // @[MapT.scala 15:7]
  assign O_4_2_2 = op_O_4_2_2; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_0_2 = op_O_5_0_2; // @[MapT.scala 15:7]
  assign O_5_1_0 = op_O_5_1_0; // @[MapT.scala 15:7]
  assign O_5_1_1 = op_O_5_1_1; // @[MapT.scala 15:7]
  assign O_5_1_2 = op_O_5_1_2; // @[MapT.scala 15:7]
  assign O_5_2_0 = op_O_5_2_0; // @[MapT.scala 15:7]
  assign O_5_2_1 = op_O_5_2_1; // @[MapT.scala 15:7]
  assign O_5_2_2 = op_O_5_2_2; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_0_2 = op_O_6_0_2; // @[MapT.scala 15:7]
  assign O_6_1_0 = op_O_6_1_0; // @[MapT.scala 15:7]
  assign O_6_1_1 = op_O_6_1_1; // @[MapT.scala 15:7]
  assign O_6_1_2 = op_O_6_1_2; // @[MapT.scala 15:7]
  assign O_6_2_0 = op_O_6_2_0; // @[MapT.scala 15:7]
  assign O_6_2_1 = op_O_6_2_1; // @[MapT.scala 15:7]
  assign O_6_2_2 = op_O_6_2_2; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_0_2 = op_O_7_0_2; // @[MapT.scala 15:7]
  assign O_7_1_0 = op_O_7_1_0; // @[MapT.scala 15:7]
  assign O_7_1_1 = op_O_7_1_1; // @[MapT.scala 15:7]
  assign O_7_1_2 = op_O_7_1_2; // @[MapT.scala 15:7]
  assign O_7_2_0 = op_O_7_2_0; // @[MapT.scala 15:7]
  assign O_7_2_1 = op_O_7_2_1; // @[MapT.scala 15:7]
  assign O_7_2_2 = op_O_7_2_2; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_0_2 = op_O_8_0_2; // @[MapT.scala 15:7]
  assign O_8_1_0 = op_O_8_1_0; // @[MapT.scala 15:7]
  assign O_8_1_1 = op_O_8_1_1; // @[MapT.scala 15:7]
  assign O_8_1_2 = op_O_8_1_2; // @[MapT.scala 15:7]
  assign O_8_2_0 = op_O_8_2_0; // @[MapT.scala 15:7]
  assign O_8_2_1 = op_O_8_2_1; // @[MapT.scala 15:7]
  assign O_8_2_2 = op_O_8_2_2; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_0_2 = op_O_9_0_2; // @[MapT.scala 15:7]
  assign O_9_1_0 = op_O_9_1_0; // @[MapT.scala 15:7]
  assign O_9_1_1 = op_O_9_1_1; // @[MapT.scala 15:7]
  assign O_9_1_2 = op_O_9_1_2; // @[MapT.scala 15:7]
  assign O_9_2_0 = op_O_9_2_0; // @[MapT.scala 15:7]
  assign O_9_2_1 = op_O_9_2_1; // @[MapT.scala 15:7]
  assign O_9_2_2 = op_O_9_2_2; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_0_2 = op_O_10_0_2; // @[MapT.scala 15:7]
  assign O_10_1_0 = op_O_10_1_0; // @[MapT.scala 15:7]
  assign O_10_1_1 = op_O_10_1_1; // @[MapT.scala 15:7]
  assign O_10_1_2 = op_O_10_1_2; // @[MapT.scala 15:7]
  assign O_10_2_0 = op_O_10_2_0; // @[MapT.scala 15:7]
  assign O_10_2_1 = op_O_10_2_1; // @[MapT.scala 15:7]
  assign O_10_2_2 = op_O_10_2_2; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_0_2 = op_O_11_0_2; // @[MapT.scala 15:7]
  assign O_11_1_0 = op_O_11_1_0; // @[MapT.scala 15:7]
  assign O_11_1_1 = op_O_11_1_1; // @[MapT.scala 15:7]
  assign O_11_1_2 = op_O_11_1_2; // @[MapT.scala 15:7]
  assign O_11_2_0 = op_O_11_2_0; // @[MapT.scala 15:7]
  assign O_11_2_1 = op_O_11_2_1; // @[MapT.scala 15:7]
  assign O_11_2_2 = op_O_11_2_2; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_0_2 = op_O_12_0_2; // @[MapT.scala 15:7]
  assign O_12_1_0 = op_O_12_1_0; // @[MapT.scala 15:7]
  assign O_12_1_1 = op_O_12_1_1; // @[MapT.scala 15:7]
  assign O_12_1_2 = op_O_12_1_2; // @[MapT.scala 15:7]
  assign O_12_2_0 = op_O_12_2_0; // @[MapT.scala 15:7]
  assign O_12_2_1 = op_O_12_2_1; // @[MapT.scala 15:7]
  assign O_12_2_2 = op_O_12_2_2; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_0_2 = op_O_13_0_2; // @[MapT.scala 15:7]
  assign O_13_1_0 = op_O_13_1_0; // @[MapT.scala 15:7]
  assign O_13_1_1 = op_O_13_1_1; // @[MapT.scala 15:7]
  assign O_13_1_2 = op_O_13_1_2; // @[MapT.scala 15:7]
  assign O_13_2_0 = op_O_13_2_0; // @[MapT.scala 15:7]
  assign O_13_2_1 = op_O_13_2_1; // @[MapT.scala 15:7]
  assign O_13_2_2 = op_O_13_2_2; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_0_2 = op_O_14_0_2; // @[MapT.scala 15:7]
  assign O_14_1_0 = op_O_14_1_0; // @[MapT.scala 15:7]
  assign O_14_1_1 = op_O_14_1_1; // @[MapT.scala 15:7]
  assign O_14_1_2 = op_O_14_1_2; // @[MapT.scala 15:7]
  assign O_14_2_0 = op_O_14_2_0; // @[MapT.scala 15:7]
  assign O_14_2_1 = op_O_14_2_1; // @[MapT.scala 15:7]
  assign O_14_2_2 = op_O_14_2_2; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_0_2 = op_O_15_0_2; // @[MapT.scala 15:7]
  assign O_15_1_0 = op_O_15_1_0; // @[MapT.scala 15:7]
  assign O_15_1_1 = op_O_15_1_1; // @[MapT.scala 15:7]
  assign O_15_1_2 = op_O_15_1_2; // @[MapT.scala 15:7]
  assign O_15_2_0 = op_O_15_2_0; // @[MapT.scala 15:7]
  assign O_15_2_1 = op_O_15_2_1; // @[MapT.scala 15:7]
  assign O_15_2_2 = op_O_15_2_2; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_0_2 = I_0_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_2 = I_0_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_0_2_0 = I_0_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_0_2_1 = I_0_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2_2 = I_0_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_2 = I_1_0_0_2; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_2 = I_1_0_1_2; // @[MapT.scala 14:10]
  assign op_I_1_0_2_0 = I_1_0_2_0; // @[MapT.scala 14:10]
  assign op_I_1_0_2_1 = I_1_0_2_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2_2 = I_1_0_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_2 = I_2_0_0_2; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_2 = I_2_0_1_2; // @[MapT.scala 14:10]
  assign op_I_2_0_2_0 = I_2_0_2_0; // @[MapT.scala 14:10]
  assign op_I_2_0_2_1 = I_2_0_2_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2_2 = I_2_0_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_2 = I_3_0_0_2; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_2 = I_3_0_1_2; // @[MapT.scala 14:10]
  assign op_I_3_0_2_0 = I_3_0_2_0; // @[MapT.scala 14:10]
  assign op_I_3_0_2_1 = I_3_0_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2_2 = I_3_0_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_2 = I_4_0_0_2; // @[MapT.scala 14:10]
  assign op_I_4_0_1_0 = I_4_0_1_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1_1 = I_4_0_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_1_2 = I_4_0_1_2; // @[MapT.scala 14:10]
  assign op_I_4_0_2_0 = I_4_0_2_0; // @[MapT.scala 14:10]
  assign op_I_4_0_2_1 = I_4_0_2_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2_2 = I_4_0_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_2 = I_5_0_0_2; // @[MapT.scala 14:10]
  assign op_I_5_0_1_0 = I_5_0_1_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1_1 = I_5_0_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_1_2 = I_5_0_1_2; // @[MapT.scala 14:10]
  assign op_I_5_0_2_0 = I_5_0_2_0; // @[MapT.scala 14:10]
  assign op_I_5_0_2_1 = I_5_0_2_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2_2 = I_5_0_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_2 = I_6_0_0_2; // @[MapT.scala 14:10]
  assign op_I_6_0_1_0 = I_6_0_1_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1_1 = I_6_0_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_1_2 = I_6_0_1_2; // @[MapT.scala 14:10]
  assign op_I_6_0_2_0 = I_6_0_2_0; // @[MapT.scala 14:10]
  assign op_I_6_0_2_1 = I_6_0_2_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2_2 = I_6_0_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_2 = I_7_0_0_2; // @[MapT.scala 14:10]
  assign op_I_7_0_1_0 = I_7_0_1_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1_1 = I_7_0_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_1_2 = I_7_0_1_2; // @[MapT.scala 14:10]
  assign op_I_7_0_2_0 = I_7_0_2_0; // @[MapT.scala 14:10]
  assign op_I_7_0_2_1 = I_7_0_2_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2_2 = I_7_0_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0_0 = I_8_0_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_0_1 = I_8_0_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0_2 = I_8_0_0_2; // @[MapT.scala 14:10]
  assign op_I_8_0_1_0 = I_8_0_1_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1_1 = I_8_0_1_1; // @[MapT.scala 14:10]
  assign op_I_8_0_1_2 = I_8_0_1_2; // @[MapT.scala 14:10]
  assign op_I_8_0_2_0 = I_8_0_2_0; // @[MapT.scala 14:10]
  assign op_I_8_0_2_1 = I_8_0_2_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2_2 = I_8_0_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0_0 = I_9_0_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_0_1 = I_9_0_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0_2 = I_9_0_0_2; // @[MapT.scala 14:10]
  assign op_I_9_0_1_0 = I_9_0_1_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1_1 = I_9_0_1_1; // @[MapT.scala 14:10]
  assign op_I_9_0_1_2 = I_9_0_1_2; // @[MapT.scala 14:10]
  assign op_I_9_0_2_0 = I_9_0_2_0; // @[MapT.scala 14:10]
  assign op_I_9_0_2_1 = I_9_0_2_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2_2 = I_9_0_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0_0 = I_10_0_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_0_1 = I_10_0_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0_2 = I_10_0_0_2; // @[MapT.scala 14:10]
  assign op_I_10_0_1_0 = I_10_0_1_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1_1 = I_10_0_1_1; // @[MapT.scala 14:10]
  assign op_I_10_0_1_2 = I_10_0_1_2; // @[MapT.scala 14:10]
  assign op_I_10_0_2_0 = I_10_0_2_0; // @[MapT.scala 14:10]
  assign op_I_10_0_2_1 = I_10_0_2_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2_2 = I_10_0_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0_0 = I_11_0_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_0_1 = I_11_0_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0_2 = I_11_0_0_2; // @[MapT.scala 14:10]
  assign op_I_11_0_1_0 = I_11_0_1_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1_1 = I_11_0_1_1; // @[MapT.scala 14:10]
  assign op_I_11_0_1_2 = I_11_0_1_2; // @[MapT.scala 14:10]
  assign op_I_11_0_2_0 = I_11_0_2_0; // @[MapT.scala 14:10]
  assign op_I_11_0_2_1 = I_11_0_2_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2_2 = I_11_0_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0_0 = I_12_0_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_0_1 = I_12_0_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0_2 = I_12_0_0_2; // @[MapT.scala 14:10]
  assign op_I_12_0_1_0 = I_12_0_1_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1_1 = I_12_0_1_1; // @[MapT.scala 14:10]
  assign op_I_12_0_1_2 = I_12_0_1_2; // @[MapT.scala 14:10]
  assign op_I_12_0_2_0 = I_12_0_2_0; // @[MapT.scala 14:10]
  assign op_I_12_0_2_1 = I_12_0_2_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2_2 = I_12_0_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0_0 = I_13_0_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_0_1 = I_13_0_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0_2 = I_13_0_0_2; // @[MapT.scala 14:10]
  assign op_I_13_0_1_0 = I_13_0_1_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1_1 = I_13_0_1_1; // @[MapT.scala 14:10]
  assign op_I_13_0_1_2 = I_13_0_1_2; // @[MapT.scala 14:10]
  assign op_I_13_0_2_0 = I_13_0_2_0; // @[MapT.scala 14:10]
  assign op_I_13_0_2_1 = I_13_0_2_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2_2 = I_13_0_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0_0 = I_14_0_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_0_1 = I_14_0_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0_2 = I_14_0_0_2; // @[MapT.scala 14:10]
  assign op_I_14_0_1_0 = I_14_0_1_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1_1 = I_14_0_1_1; // @[MapT.scala 14:10]
  assign op_I_14_0_1_2 = I_14_0_1_2; // @[MapT.scala 14:10]
  assign op_I_14_0_2_0 = I_14_0_2_0; // @[MapT.scala 14:10]
  assign op_I_14_0_2_1 = I_14_0_2_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2_2 = I_14_0_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0_0 = I_15_0_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_0_1 = I_15_0_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0_2 = I_15_0_0_2; // @[MapT.scala 14:10]
  assign op_I_15_0_1_0 = I_15_0_1_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1_1 = I_15_0_1_1; // @[MapT.scala 14:10]
  assign op_I_15_0_1_2 = I_15_0_1_2; // @[MapT.scala 14:10]
  assign op_I_15_0_2_0 = I_15_0_2_0; // @[MapT.scala 14:10]
  assign op_I_15_0_2_1 = I_15_0_2_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2_2 = I_15_0_2_2; // @[MapT.scala 14:10]
endmodule
module InitialDelayCounter(
  input   clock,
  input   reset,
  output  valid_down
);
  reg  value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire  _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 1'h1; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 1'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 1'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module AtomTuple(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0,
  input  [7:0] I1,
  output [7:0] O_t0b,
  output [7:0] O_t1b
);
  assign valid_down = valid_up; // @[Tuple.scala 51:14]
  assign O_t0b = I0; // @[Tuple.scala 49:9]
  assign O_t1b = I1; // @[Tuple.scala 50:9]
endmodule
module Map2S_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I0_2,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  input  [7:0] I1_2,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b,
  output [7:0] O_2_t0b,
  output [7:0] O_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  AtomTuple other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0(other_ops_1_I0),
    .I1(other_ops_1_I1),
    .O_t0b(other_ops_1_O_t0b),
    .O_t1b(other_ops_1_O_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign O_2_t0b = other_ops_1_O_t0b; // @[Map2S.scala 24:12]
  assign O_2_t1b = other_ops_1_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0 = I0_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1 = I1_2; // @[Map2S.scala 23:43]
endmodule
module Map2S_9(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_0_2,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_1_2,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_2_2,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b,
  output [7:0] O_0_1_t0b,
  output [7:0] O_0_1_t1b,
  output [7:0] O_0_2_t0b,
  output [7:0] O_0_2_t1b,
  output [7:0] O_1_0_t0b,
  output [7:0] O_1_0_t1b,
  output [7:0] O_1_1_t0b,
  output [7:0] O_1_1_t1b,
  output [7:0] O_1_2_t0b,
  output [7:0] O_1_2_t1b,
  output [7:0] O_2_0_t0b,
  output [7:0] O_2_0_t1b,
  output [7:0] O_2_1_t0b,
  output [7:0] O_2_1_t1b,
  output [7:0] O_2_2_t0b,
  output [7:0] O_2_2_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_2; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_2_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_2_t1b; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_2; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_2_t1b; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  Map2S_8 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I0_2(fst_op_I0_2),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .I1_2(fst_op_I1_2),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b),
    .O_2_t0b(fst_op_O_2_t0b),
    .O_2_t1b(fst_op_O_2_t1b)
  );
  Map2S_8 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I0_2(other_ops_0_I0_2),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .I1_2(other_ops_0_I1_2),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b),
    .O_2_t0b(other_ops_0_O_2_t0b),
    .O_2_t1b(other_ops_0_O_2_t1b)
  );
  Map2S_8 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I0_2(other_ops_1_I0_2),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .I1_2(other_ops_1_I1_2),
    .O_0_t0b(other_ops_1_O_0_t0b),
    .O_0_t1b(other_ops_1_O_0_t1b),
    .O_1_t0b(other_ops_1_O_1_t0b),
    .O_1_t1b(other_ops_1_O_1_t1b),
    .O_2_t0b(other_ops_1_O_2_t0b),
    .O_2_t1b(other_ops_1_O_2_t1b)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_0_2_t0b = fst_op_O_2_t0b; // @[Map2S.scala 19:8]
  assign O_0_2_t1b = fst_op_O_2_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_1_2_t0b = other_ops_0_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_1_2_t1b = other_ops_0_O_2_t1b; // @[Map2S.scala 24:12]
  assign O_2_0_t0b = other_ops_1_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_2_0_t1b = other_ops_1_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_2_1_t0b = other_ops_1_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_2_1_t1b = other_ops_1_O_1_t1b; // @[Map2S.scala 24:12]
  assign O_2_2_t0b = other_ops_1_O_2_t0b; // @[Map2S.scala 24:12]
  assign O_2_2_t1b = other_ops_1_O_2_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I0_2 = I0_0_2; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 8'h0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 8'h1; // @[Map2S.scala 18:13]
  assign fst_op_I1_2 = 8'h0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_2 = I0_1_2; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 8'h2; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_2 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_2 = I0_2_2; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = 8'h0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_2 = 8'h0; // @[Map2S.scala 23:43]
endmodule
module LShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  wire [262:0] _GEN_0; // @[Arithmetic.scala 301:25]
  wire [262:0] _T; // @[Arithmetic.scala 301:25]
  assign _GEN_0 = {{255'd0}, I_t0b}; // @[Arithmetic.scala 301:25]
  assign _T = _GEN_0 << I_t1b; // @[Arithmetic.scala 301:25]
  assign valid_down = valid_up; // @[Arithmetic.scala 303:14]
  assign O = _T[7:0]; // @[Arithmetic.scala 301:7]
endmodule
module MapS_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  input  [7:0] I_2_t0b,
  input  [7:0] I_2_t1b,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  LShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  LShift other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  LShift other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_t0b(other_ops_1_I_t0b),
    .I_t1b(other_ops_1_I_t1b),
    .O(other_ops_1_O)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign O_2 = other_ops_1_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_t0b = I_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_t1b = I_2_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_5(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  input  [7:0] I_0_1_t0b,
  input  [7:0] I_0_1_t1b,
  input  [7:0] I_0_2_t0b,
  input  [7:0] I_0_2_t1b,
  input  [7:0] I_1_0_t0b,
  input  [7:0] I_1_0_t1b,
  input  [7:0] I_1_1_t0b,
  input  [7:0] I_1_1_t1b,
  input  [7:0] I_1_2_t0b,
  input  [7:0] I_1_2_t1b,
  input  [7:0] I_2_0_t0b,
  input  [7:0] I_2_0_t1b,
  input  [7:0] I_2_1_t0b,
  input  [7:0] I_2_1_t1b,
  input  [7:0] I_2_2_t0b,
  input  [7:0] I_2_2_t1b,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_0_2,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_1_2,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_2_2
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_2; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_2; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_2; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  MapS_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .I_2_t0b(fst_op_I_2_t0b),
    .I_2_t1b(fst_op_I_2_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1),
    .O_2(fst_op_O_2)
  );
  MapS_4 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .I_2_t0b(other_ops_0_I_2_t0b),
    .I_2_t1b(other_ops_0_I_2_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1),
    .O_2(other_ops_0_O_2)
  );
  MapS_4 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_t0b(other_ops_1_I_0_t0b),
    .I_0_t1b(other_ops_1_I_0_t1b),
    .I_1_t0b(other_ops_1_I_1_t0b),
    .I_1_t1b(other_ops_1_I_1_t1b),
    .I_2_t0b(other_ops_1_I_2_t0b),
    .I_2_t1b(other_ops_1_I_2_t1b),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1),
    .O_2(other_ops_1_O_2)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_0_2 = fst_op_O_2; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_1_2 = other_ops_0_O_2; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_2_2 = other_ops_1_O_2; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t0b = I_0_2_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_2_t1b = I_0_2_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t0b = I_1_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_t1b = I_1_2_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_t0b = I_2_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_t1b = I_2_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t0b = I_2_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_t1b = I_2_1_t1b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t0b = I_2_2_t0b; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_t1b = I_2_2_t1b; // @[MapS.scala 20:41]
endmodule
module AddNoValid(
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign O = I_t0b + I_t1b; // @[Arithmetic.scala 122:7]
endmodule
module ReduceS(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  output [7:0] O_0
);
  wire [7:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_1_O; // @[ReduceS.scala 20:43]
  reg [7:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  AddNoValid AddNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_1_I_t0b),
    .I_t1b(AddNoValid_1_I_t1b),
    .O(AddNoValid_1_O)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = I_2; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = AddNoValid_1_O; // @[ReduceS.scala 36:18]
  assign AddNoValid_1_I_t0b = I_0; // @[ReduceS.scala 43:18]
  assign AddNoValid_1_I_t1b = I_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module MapS_6(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0,
  output [7:0] O_1_0,
  output [7:0] O_2_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  ReduceS fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .I_2(fst_op_I_2),
    .O_0(fst_op_O_0)
  );
  ReduceS other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .I_2(other_ops_0_I_2),
    .O_0(other_ops_0_O_0)
  );
  ReduceS other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0(other_ops_1_I_0),
    .I_1(other_ops_1_I_1),
    .I_2(other_ops_1_I_2),
    .O_0(other_ops_1_O_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T & other_ops_1_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_2 = I_0_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2 = I_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0 = I_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1 = I_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2 = I_2_2; // @[MapS.scala 20:41]
endmodule
module MapSNoValid(
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 28:22]
  wire [7:0] fst_op_O; // @[MapS.scala 28:22]
  AddNoValid fst_op ( // @[MapS.scala 28:22]
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign O_0 = fst_op_O; // @[MapS.scala 35:8]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 34:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 34:12]
endmodule
module ReduceS_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  input  [7:0] I_2_0,
  output [7:0] O_0_0
);
  wire [7:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_1_O_0; // @[ReduceS.scala 20:43]
  reg [7:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  MapSNoValid MapSNoValid_1 ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_1_I_0_t0b),
    .I_0_t1b(MapSNoValid_1_I_0_t1b),
    .O_0(MapSNoValid_1_O_0)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = I_2_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = MapSNoValid_1_O_0; // @[ReduceS.scala 36:18]
  assign MapSNoValid_1_I_0_t0b = I_0_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_1_I_0_t1b = I_1_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module InitialDelayCounter_1(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [1:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [1:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 2'h3; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 2'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 2'h3; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 2'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Map2S_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I1_0,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
endmodule
module Map2S_11(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I1_0_0,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  Map2S_10 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I1_0(fst_op_I1_0),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b)
  );
  assign valid_down = fst_op_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
endmodule
module RShift(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_t0b,
  input  [7:0] I_t1b,
  output [7:0] O
);
  assign valid_down = valid_up; // @[Arithmetic.scala 272:14]
  assign O = I_t0b >> I_t1b; // @[Arithmetic.scala 270:7]
endmodule
module MapS_7(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  output [7:0] O_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  RShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
endmodule
module MapS_8(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  output [7:0] O_0_0
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  MapS_7 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .O_0(fst_op_O_0)
  );
  assign valid_down = fst_op_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
endmodule
module Module_0(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_0_2,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_1_2,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_2_2,
  output [7:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n110_valid_up; // @[Top.scala 17:22]
  wire  n110_valid_down; // @[Top.scala 17:22]
  wire [7:0] n110_I0_0_0; // @[Top.scala 17:22]
  wire [7:0] n110_I0_0_1; // @[Top.scala 17:22]
  wire [7:0] n110_I0_0_2; // @[Top.scala 17:22]
  wire [7:0] n110_I0_1_0; // @[Top.scala 17:22]
  wire [7:0] n110_I0_1_1; // @[Top.scala 17:22]
  wire [7:0] n110_I0_1_2; // @[Top.scala 17:22]
  wire [7:0] n110_I0_2_0; // @[Top.scala 17:22]
  wire [7:0] n110_I0_2_1; // @[Top.scala 17:22]
  wire [7:0] n110_I0_2_2; // @[Top.scala 17:22]
  wire [7:0] n110_O_0_0_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_0_0_t1b; // @[Top.scala 17:22]
  wire [7:0] n110_O_0_1_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_0_1_t1b; // @[Top.scala 17:22]
  wire [7:0] n110_O_0_2_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_0_2_t1b; // @[Top.scala 17:22]
  wire [7:0] n110_O_1_0_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_1_0_t1b; // @[Top.scala 17:22]
  wire [7:0] n110_O_1_1_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_1_1_t1b; // @[Top.scala 17:22]
  wire [7:0] n110_O_1_2_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_1_2_t1b; // @[Top.scala 17:22]
  wire [7:0] n110_O_2_0_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_2_0_t1b; // @[Top.scala 17:22]
  wire [7:0] n110_O_2_1_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_2_1_t1b; // @[Top.scala 17:22]
  wire [7:0] n110_O_2_2_t0b; // @[Top.scala 17:22]
  wire [7:0] n110_O_2_2_t1b; // @[Top.scala 17:22]
  wire  n121_valid_up; // @[Top.scala 21:22]
  wire  n121_valid_down; // @[Top.scala 21:22]
  wire [7:0] n121_I_0_0_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_0_0_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_I_0_1_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_0_1_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_I_0_2_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_0_2_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_I_1_0_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_1_0_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_I_1_1_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_1_1_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_I_1_2_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_1_2_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_I_2_0_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_2_0_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_I_2_1_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_2_1_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_I_2_2_t0b; // @[Top.scala 21:22]
  wire [7:0] n121_I_2_2_t1b; // @[Top.scala 21:22]
  wire [7:0] n121_O_0_0; // @[Top.scala 21:22]
  wire [7:0] n121_O_0_1; // @[Top.scala 21:22]
  wire [7:0] n121_O_0_2; // @[Top.scala 21:22]
  wire [7:0] n121_O_1_0; // @[Top.scala 21:22]
  wire [7:0] n121_O_1_1; // @[Top.scala 21:22]
  wire [7:0] n121_O_1_2; // @[Top.scala 21:22]
  wire [7:0] n121_O_2_0; // @[Top.scala 21:22]
  wire [7:0] n121_O_2_1; // @[Top.scala 21:22]
  wire [7:0] n121_O_2_2; // @[Top.scala 21:22]
  wire  n126_clock; // @[Top.scala 24:22]
  wire  n126_reset; // @[Top.scala 24:22]
  wire  n126_valid_up; // @[Top.scala 24:22]
  wire  n126_valid_down; // @[Top.scala 24:22]
  wire [7:0] n126_I_0_0; // @[Top.scala 24:22]
  wire [7:0] n126_I_0_1; // @[Top.scala 24:22]
  wire [7:0] n126_I_0_2; // @[Top.scala 24:22]
  wire [7:0] n126_I_1_0; // @[Top.scala 24:22]
  wire [7:0] n126_I_1_1; // @[Top.scala 24:22]
  wire [7:0] n126_I_1_2; // @[Top.scala 24:22]
  wire [7:0] n126_I_2_0; // @[Top.scala 24:22]
  wire [7:0] n126_I_2_1; // @[Top.scala 24:22]
  wire [7:0] n126_I_2_2; // @[Top.scala 24:22]
  wire [7:0] n126_O_0_0; // @[Top.scala 24:22]
  wire [7:0] n126_O_1_0; // @[Top.scala 24:22]
  wire [7:0] n126_O_2_0; // @[Top.scala 24:22]
  wire  n131_clock; // @[Top.scala 27:22]
  wire  n131_reset; // @[Top.scala 27:22]
  wire  n131_valid_up; // @[Top.scala 27:22]
  wire  n131_valid_down; // @[Top.scala 27:22]
  wire [7:0] n131_I_0_0; // @[Top.scala 27:22]
  wire [7:0] n131_I_1_0; // @[Top.scala 27:22]
  wire [7:0] n131_I_2_0; // @[Top.scala 27:22]
  wire [7:0] n131_O_0_0; // @[Top.scala 27:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n134_valid_up; // @[Top.scala 31:22]
  wire  n134_valid_down; // @[Top.scala 31:22]
  wire [7:0] n134_I0_0_0; // @[Top.scala 31:22]
  wire [7:0] n134_I1_0_0; // @[Top.scala 31:22]
  wire [7:0] n134_O_0_0_t0b; // @[Top.scala 31:22]
  wire [7:0] n134_O_0_0_t1b; // @[Top.scala 31:22]
  wire  n145_valid_up; // @[Top.scala 35:22]
  wire  n145_valid_down; // @[Top.scala 35:22]
  wire [7:0] n145_I_0_0_t0b; // @[Top.scala 35:22]
  wire [7:0] n145_I_0_0_t1b; // @[Top.scala 35:22]
  wire [7:0] n145_O_0_0; // @[Top.scala 35:22]
  InitialDelayCounter InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_9 n110 ( // @[Top.scala 17:22]
    .valid_up(n110_valid_up),
    .valid_down(n110_valid_down),
    .I0_0_0(n110_I0_0_0),
    .I0_0_1(n110_I0_0_1),
    .I0_0_2(n110_I0_0_2),
    .I0_1_0(n110_I0_1_0),
    .I0_1_1(n110_I0_1_1),
    .I0_1_2(n110_I0_1_2),
    .I0_2_0(n110_I0_2_0),
    .I0_2_1(n110_I0_2_1),
    .I0_2_2(n110_I0_2_2),
    .O_0_0_t0b(n110_O_0_0_t0b),
    .O_0_0_t1b(n110_O_0_0_t1b),
    .O_0_1_t0b(n110_O_0_1_t0b),
    .O_0_1_t1b(n110_O_0_1_t1b),
    .O_0_2_t0b(n110_O_0_2_t0b),
    .O_0_2_t1b(n110_O_0_2_t1b),
    .O_1_0_t0b(n110_O_1_0_t0b),
    .O_1_0_t1b(n110_O_1_0_t1b),
    .O_1_1_t0b(n110_O_1_1_t0b),
    .O_1_1_t1b(n110_O_1_1_t1b),
    .O_1_2_t0b(n110_O_1_2_t0b),
    .O_1_2_t1b(n110_O_1_2_t1b),
    .O_2_0_t0b(n110_O_2_0_t0b),
    .O_2_0_t1b(n110_O_2_0_t1b),
    .O_2_1_t0b(n110_O_2_1_t0b),
    .O_2_1_t1b(n110_O_2_1_t1b),
    .O_2_2_t0b(n110_O_2_2_t0b),
    .O_2_2_t1b(n110_O_2_2_t1b)
  );
  MapS_5 n121 ( // @[Top.scala 21:22]
    .valid_up(n121_valid_up),
    .valid_down(n121_valid_down),
    .I_0_0_t0b(n121_I_0_0_t0b),
    .I_0_0_t1b(n121_I_0_0_t1b),
    .I_0_1_t0b(n121_I_0_1_t0b),
    .I_0_1_t1b(n121_I_0_1_t1b),
    .I_0_2_t0b(n121_I_0_2_t0b),
    .I_0_2_t1b(n121_I_0_2_t1b),
    .I_1_0_t0b(n121_I_1_0_t0b),
    .I_1_0_t1b(n121_I_1_0_t1b),
    .I_1_1_t0b(n121_I_1_1_t0b),
    .I_1_1_t1b(n121_I_1_1_t1b),
    .I_1_2_t0b(n121_I_1_2_t0b),
    .I_1_2_t1b(n121_I_1_2_t1b),
    .I_2_0_t0b(n121_I_2_0_t0b),
    .I_2_0_t1b(n121_I_2_0_t1b),
    .I_2_1_t0b(n121_I_2_1_t0b),
    .I_2_1_t1b(n121_I_2_1_t1b),
    .I_2_2_t0b(n121_I_2_2_t0b),
    .I_2_2_t1b(n121_I_2_2_t1b),
    .O_0_0(n121_O_0_0),
    .O_0_1(n121_O_0_1),
    .O_0_2(n121_O_0_2),
    .O_1_0(n121_O_1_0),
    .O_1_1(n121_O_1_1),
    .O_1_2(n121_O_1_2),
    .O_2_0(n121_O_2_0),
    .O_2_1(n121_O_2_1),
    .O_2_2(n121_O_2_2)
  );
  MapS_6 n126 ( // @[Top.scala 24:22]
    .clock(n126_clock),
    .reset(n126_reset),
    .valid_up(n126_valid_up),
    .valid_down(n126_valid_down),
    .I_0_0(n126_I_0_0),
    .I_0_1(n126_I_0_1),
    .I_0_2(n126_I_0_2),
    .I_1_0(n126_I_1_0),
    .I_1_1(n126_I_1_1),
    .I_1_2(n126_I_1_2),
    .I_2_0(n126_I_2_0),
    .I_2_1(n126_I_2_1),
    .I_2_2(n126_I_2_2),
    .O_0_0(n126_O_0_0),
    .O_1_0(n126_O_1_0),
    .O_2_0(n126_O_2_0)
  );
  ReduceS_1 n131 ( // @[Top.scala 27:22]
    .clock(n131_clock),
    .reset(n131_reset),
    .valid_up(n131_valid_up),
    .valid_down(n131_valid_down),
    .I_0_0(n131_I_0_0),
    .I_1_0(n131_I_1_0),
    .I_2_0(n131_I_2_0),
    .O_0_0(n131_O_0_0)
  );
  InitialDelayCounter_1 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_11 n134 ( // @[Top.scala 31:22]
    .valid_up(n134_valid_up),
    .valid_down(n134_valid_down),
    .I0_0_0(n134_I0_0_0),
    .I1_0_0(n134_I1_0_0),
    .O_0_0_t0b(n134_O_0_0_t0b),
    .O_0_0_t1b(n134_O_0_0_t1b)
  );
  MapS_8 n145 ( // @[Top.scala 35:22]
    .valid_up(n145_valid_up),
    .valid_down(n145_valid_down),
    .I_0_0_t0b(n145_I_0_0_t0b),
    .I_0_0_t1b(n145_I_0_0_t1b),
    .O_0_0(n145_O_0_0)
  );
  assign valid_down = n145_valid_down; // @[Top.scala 39:16]
  assign O_0_0 = n145_O_0_0; // @[Top.scala 38:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n110_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 20:19]
  assign n110_I0_0_0 = I_0_0; // @[Top.scala 18:13]
  assign n110_I0_0_1 = I_0_1; // @[Top.scala 18:13]
  assign n110_I0_0_2 = I_0_2; // @[Top.scala 18:13]
  assign n110_I0_1_0 = I_1_0; // @[Top.scala 18:13]
  assign n110_I0_1_1 = I_1_1; // @[Top.scala 18:13]
  assign n110_I0_1_2 = I_1_2; // @[Top.scala 18:13]
  assign n110_I0_2_0 = I_2_0; // @[Top.scala 18:13]
  assign n110_I0_2_1 = I_2_1; // @[Top.scala 18:13]
  assign n110_I0_2_2 = I_2_2; // @[Top.scala 18:13]
  assign n121_valid_up = n110_valid_down; // @[Top.scala 23:19]
  assign n121_I_0_0_t0b = n110_O_0_0_t0b; // @[Top.scala 22:12]
  assign n121_I_0_0_t1b = n110_O_0_0_t1b; // @[Top.scala 22:12]
  assign n121_I_0_1_t0b = n110_O_0_1_t0b; // @[Top.scala 22:12]
  assign n121_I_0_1_t1b = n110_O_0_1_t1b; // @[Top.scala 22:12]
  assign n121_I_0_2_t0b = n110_O_0_2_t0b; // @[Top.scala 22:12]
  assign n121_I_0_2_t1b = n110_O_0_2_t1b; // @[Top.scala 22:12]
  assign n121_I_1_0_t0b = n110_O_1_0_t0b; // @[Top.scala 22:12]
  assign n121_I_1_0_t1b = n110_O_1_0_t1b; // @[Top.scala 22:12]
  assign n121_I_1_1_t0b = n110_O_1_1_t0b; // @[Top.scala 22:12]
  assign n121_I_1_1_t1b = n110_O_1_1_t1b; // @[Top.scala 22:12]
  assign n121_I_1_2_t0b = n110_O_1_2_t0b; // @[Top.scala 22:12]
  assign n121_I_1_2_t1b = n110_O_1_2_t1b; // @[Top.scala 22:12]
  assign n121_I_2_0_t0b = n110_O_2_0_t0b; // @[Top.scala 22:12]
  assign n121_I_2_0_t1b = n110_O_2_0_t1b; // @[Top.scala 22:12]
  assign n121_I_2_1_t0b = n110_O_2_1_t0b; // @[Top.scala 22:12]
  assign n121_I_2_1_t1b = n110_O_2_1_t1b; // @[Top.scala 22:12]
  assign n121_I_2_2_t0b = n110_O_2_2_t0b; // @[Top.scala 22:12]
  assign n121_I_2_2_t1b = n110_O_2_2_t1b; // @[Top.scala 22:12]
  assign n126_clock = clock;
  assign n126_reset = reset;
  assign n126_valid_up = n121_valid_down; // @[Top.scala 26:19]
  assign n126_I_0_0 = n121_O_0_0; // @[Top.scala 25:12]
  assign n126_I_0_1 = n121_O_0_1; // @[Top.scala 25:12]
  assign n126_I_0_2 = n121_O_0_2; // @[Top.scala 25:12]
  assign n126_I_1_0 = n121_O_1_0; // @[Top.scala 25:12]
  assign n126_I_1_1 = n121_O_1_1; // @[Top.scala 25:12]
  assign n126_I_1_2 = n121_O_1_2; // @[Top.scala 25:12]
  assign n126_I_2_0 = n121_O_2_0; // @[Top.scala 25:12]
  assign n126_I_2_1 = n121_O_2_1; // @[Top.scala 25:12]
  assign n126_I_2_2 = n121_O_2_2; // @[Top.scala 25:12]
  assign n131_clock = clock;
  assign n131_reset = reset;
  assign n131_valid_up = n126_valid_down; // @[Top.scala 29:19]
  assign n131_I_0_0 = n126_O_0_0; // @[Top.scala 28:12]
  assign n131_I_1_0 = n126_O_1_0; // @[Top.scala 28:12]
  assign n131_I_2_0 = n126_O_2_0; // @[Top.scala 28:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n134_valid_up = n131_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 34:19]
  assign n134_I0_0_0 = n131_O_0_0; // @[Top.scala 32:13]
  assign n134_I1_0_0 = 8'h4; // @[Top.scala 33:13]
  assign n145_valid_up = n134_valid_down; // @[Top.scala 37:19]
  assign n145_I_0_0_t0b = n134_O_0_0_t0b; // @[Top.scala 36:12]
  assign n145_I_0_0_t1b = n134_O_0_0_t1b; // @[Top.scala 36:12]
endmodule
module MapS_9(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_8_1_2,
  input  [7:0] I_8_2_0,
  input  [7:0] I_8_2_1,
  input  [7:0] I_8_2_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_9_1_2,
  input  [7:0] I_9_2_0,
  input  [7:0] I_9_2_1,
  input  [7:0] I_9_2_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_10_1_2,
  input  [7:0] I_10_2_0,
  input  [7:0] I_10_2_1,
  input  [7:0] I_10_2_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_11_1_2,
  input  [7:0] I_11_2_0,
  input  [7:0] I_11_2_1,
  input  [7:0] I_11_2_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_12_1_2,
  input  [7:0] I_12_2_0,
  input  [7:0] I_12_2_1,
  input  [7:0] I_12_2_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_13_1_2,
  input  [7:0] I_13_2_0,
  input  [7:0] I_13_2_1,
  input  [7:0] I_13_2_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_14_1_2,
  input  [7:0] I_14_2_0,
  input  [7:0] I_14_2_1,
  input  [7:0] I_14_2_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  input  [7:0] I_15_1_2,
  input  [7:0] I_15_2_0,
  input  [7:0] I_15_2_1,
  input  [7:0] I_15_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_2_2; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_7_clock; // @[MapS.scala 10:86]
  wire  other_ops_7_reset; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_8_clock; // @[MapS.scala 10:86]
  wire  other_ops_8_reset; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_9_clock; // @[MapS.scala 10:86]
  wire  other_ops_9_reset; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_10_clock; // @[MapS.scala 10:86]
  wire  other_ops_10_reset; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_11_clock; // @[MapS.scala 10:86]
  wire  other_ops_11_reset; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_12_clock; // @[MapS.scala 10:86]
  wire  other_ops_12_reset; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_13_clock; // @[MapS.scala 10:86]
  wire  other_ops_13_reset; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_14_clock; // @[MapS.scala 10:86]
  wire  other_ops_14_reset; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_2_2; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Module_0 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_0_2(fst_op_I_0_2),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .I_1_2(fst_op_I_1_2),
    .I_2_0(fst_op_I_2_0),
    .I_2_1(fst_op_I_2_1),
    .I_2_2(fst_op_I_2_2),
    .O_0_0(fst_op_O_0_0)
  );
  Module_0 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_0_2(other_ops_0_I_0_2),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .I_1_2(other_ops_0_I_1_2),
    .I_2_0(other_ops_0_I_2_0),
    .I_2_1(other_ops_0_I_2_1),
    .I_2_2(other_ops_0_I_2_2),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_0 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_0_2(other_ops_1_I_0_2),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .I_1_2(other_ops_1_I_1_2),
    .I_2_0(other_ops_1_I_2_0),
    .I_2_1(other_ops_1_I_2_1),
    .I_2_2(other_ops_1_I_2_2),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_0 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_0_2(other_ops_2_I_0_2),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .I_1_2(other_ops_2_I_1_2),
    .I_2_0(other_ops_2_I_2_0),
    .I_2_1(other_ops_2_I_2_1),
    .I_2_2(other_ops_2_I_2_2),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_0 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_0_2(other_ops_3_I_0_2),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .I_1_2(other_ops_3_I_1_2),
    .I_2_0(other_ops_3_I_2_0),
    .I_2_1(other_ops_3_I_2_1),
    .I_2_2(other_ops_3_I_2_2),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_0 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_0_2(other_ops_4_I_0_2),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .I_1_2(other_ops_4_I_1_2),
    .I_2_0(other_ops_4_I_2_0),
    .I_2_1(other_ops_4_I_2_1),
    .I_2_2(other_ops_4_I_2_2),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_0 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_0_2(other_ops_5_I_0_2),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .I_1_2(other_ops_5_I_1_2),
    .I_2_0(other_ops_5_I_2_0),
    .I_2_1(other_ops_5_I_2_1),
    .I_2_2(other_ops_5_I_2_2),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_0 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_0_2(other_ops_6_I_0_2),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .I_1_2(other_ops_6_I_1_2),
    .I_2_0(other_ops_6_I_2_0),
    .I_2_1(other_ops_6_I_2_1),
    .I_2_2(other_ops_6_I_2_2),
    .O_0_0(other_ops_6_O_0_0)
  );
  Module_0 other_ops_7 ( // @[MapS.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_0_2(other_ops_7_I_0_2),
    .I_1_0(other_ops_7_I_1_0),
    .I_1_1(other_ops_7_I_1_1),
    .I_1_2(other_ops_7_I_1_2),
    .I_2_0(other_ops_7_I_2_0),
    .I_2_1(other_ops_7_I_2_1),
    .I_2_2(other_ops_7_I_2_2),
    .O_0_0(other_ops_7_O_0_0)
  );
  Module_0 other_ops_8 ( // @[MapS.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_0_2(other_ops_8_I_0_2),
    .I_1_0(other_ops_8_I_1_0),
    .I_1_1(other_ops_8_I_1_1),
    .I_1_2(other_ops_8_I_1_2),
    .I_2_0(other_ops_8_I_2_0),
    .I_2_1(other_ops_8_I_2_1),
    .I_2_2(other_ops_8_I_2_2),
    .O_0_0(other_ops_8_O_0_0)
  );
  Module_0 other_ops_9 ( // @[MapS.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_0_2(other_ops_9_I_0_2),
    .I_1_0(other_ops_9_I_1_0),
    .I_1_1(other_ops_9_I_1_1),
    .I_1_2(other_ops_9_I_1_2),
    .I_2_0(other_ops_9_I_2_0),
    .I_2_1(other_ops_9_I_2_1),
    .I_2_2(other_ops_9_I_2_2),
    .O_0_0(other_ops_9_O_0_0)
  );
  Module_0 other_ops_10 ( // @[MapS.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_0_2(other_ops_10_I_0_2),
    .I_1_0(other_ops_10_I_1_0),
    .I_1_1(other_ops_10_I_1_1),
    .I_1_2(other_ops_10_I_1_2),
    .I_2_0(other_ops_10_I_2_0),
    .I_2_1(other_ops_10_I_2_1),
    .I_2_2(other_ops_10_I_2_2),
    .O_0_0(other_ops_10_O_0_0)
  );
  Module_0 other_ops_11 ( // @[MapS.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_0_2(other_ops_11_I_0_2),
    .I_1_0(other_ops_11_I_1_0),
    .I_1_1(other_ops_11_I_1_1),
    .I_1_2(other_ops_11_I_1_2),
    .I_2_0(other_ops_11_I_2_0),
    .I_2_1(other_ops_11_I_2_1),
    .I_2_2(other_ops_11_I_2_2),
    .O_0_0(other_ops_11_O_0_0)
  );
  Module_0 other_ops_12 ( // @[MapS.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_0_2(other_ops_12_I_0_2),
    .I_1_0(other_ops_12_I_1_0),
    .I_1_1(other_ops_12_I_1_1),
    .I_1_2(other_ops_12_I_1_2),
    .I_2_0(other_ops_12_I_2_0),
    .I_2_1(other_ops_12_I_2_1),
    .I_2_2(other_ops_12_I_2_2),
    .O_0_0(other_ops_12_O_0_0)
  );
  Module_0 other_ops_13 ( // @[MapS.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_0_2(other_ops_13_I_0_2),
    .I_1_0(other_ops_13_I_1_0),
    .I_1_1(other_ops_13_I_1_1),
    .I_1_2(other_ops_13_I_1_2),
    .I_2_0(other_ops_13_I_2_0),
    .I_2_1(other_ops_13_I_2_1),
    .I_2_2(other_ops_13_I_2_2),
    .O_0_0(other_ops_13_O_0_0)
  );
  Module_0 other_ops_14 ( // @[MapS.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_0_2(other_ops_14_I_0_2),
    .I_1_0(other_ops_14_I_1_0),
    .I_1_1(other_ops_14_I_1_1),
    .I_1_2(other_ops_14_I_1_2),
    .I_2_0(other_ops_14_I_2_0),
    .I_2_1(other_ops_14_I_2_1),
    .I_2_2(other_ops_14_I_2_2),
    .O_0_0(other_ops_14_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_2 = I_0_0_2; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_2 = I_0_1_2; // @[MapS.scala 16:12]
  assign fst_op_I_2_0 = I_0_2_0; // @[MapS.scala 16:12]
  assign fst_op_I_2_1 = I_0_2_1; // @[MapS.scala 16:12]
  assign fst_op_I_2_2 = I_0_2_2; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_2 = I_1_0_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_2 = I_1_1_2; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_0 = I_1_2_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_1 = I_1_2_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_2_2 = I_1_2_2; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_2 = I_2_0_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_2 = I_2_1_2; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_0 = I_2_2_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_1 = I_2_2_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_2_2 = I_2_2_2; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_2 = I_3_0_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_2 = I_3_1_2; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_0 = I_3_2_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_1 = I_3_2_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_2_2 = I_3_2_2; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_2 = I_4_0_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_2 = I_4_1_2; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_0 = I_4_2_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_1 = I_4_2_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_2_2 = I_4_2_2; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_2 = I_5_0_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_2 = I_5_1_2; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_0 = I_5_2_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_1 = I_5_2_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_2_2 = I_5_2_2; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_2 = I_6_0_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_2 = I_6_1_2; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_0 = I_6_2_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_1 = I_6_2_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_2_2 = I_6_2_2; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_2 = I_7_0_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_2 = I_7_1_2; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_0 = I_7_2_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_1 = I_7_2_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_2_2 = I_7_2_2; // @[MapS.scala 20:41]
  assign other_ops_7_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_7_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_2 = I_8_0_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_0 = I_8_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_1 = I_8_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_2 = I_8_1_2; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_0 = I_8_2_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_1 = I_8_2_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_2_2 = I_8_2_2; // @[MapS.scala 20:41]
  assign other_ops_8_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_8_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_2 = I_9_0_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_0 = I_9_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_1 = I_9_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_2 = I_9_1_2; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_0 = I_9_2_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_1 = I_9_2_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_2_2 = I_9_2_2; // @[MapS.scala 20:41]
  assign other_ops_9_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_9_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_2 = I_10_0_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_0 = I_10_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_1 = I_10_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_2 = I_10_1_2; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_0 = I_10_2_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_1 = I_10_2_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_2_2 = I_10_2_2; // @[MapS.scala 20:41]
  assign other_ops_10_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_10_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_2 = I_11_0_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_0 = I_11_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_1 = I_11_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_2 = I_11_1_2; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_0 = I_11_2_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_1 = I_11_2_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_2_2 = I_11_2_2; // @[MapS.scala 20:41]
  assign other_ops_11_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_11_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_2 = I_12_0_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_0 = I_12_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_1 = I_12_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_2 = I_12_1_2; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_0 = I_12_2_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_1 = I_12_2_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_2_2 = I_12_2_2; // @[MapS.scala 20:41]
  assign other_ops_12_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_12_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_2 = I_13_0_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_0 = I_13_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_1 = I_13_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_2 = I_13_1_2; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_0 = I_13_2_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_1 = I_13_2_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_2_2 = I_13_2_2; // @[MapS.scala 20:41]
  assign other_ops_13_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_13_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_2 = I_14_0_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_0 = I_14_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_1 = I_14_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_2 = I_14_1_2; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_0 = I_14_2_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_1 = I_14_2_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_2_2 = I_14_2_2; // @[MapS.scala 20:41]
  assign other_ops_14_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_14_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_2 = I_15_0_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_0 = I_15_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_1 = I_15_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_2 = I_15_1_2; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_0 = I_15_2_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_1 = I_15_2_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_2_2 = I_15_2_2; // @[MapS.scala 20:41]
endmodule
module MapT_8(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_0_2,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_0_1_2,
  input  [7:0] I_0_2_0,
  input  [7:0] I_0_2_1,
  input  [7:0] I_0_2_2,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_0_2,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_1_1_2,
  input  [7:0] I_1_2_0,
  input  [7:0] I_1_2_1,
  input  [7:0] I_1_2_2,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_0_2,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_2_1_2,
  input  [7:0] I_2_2_0,
  input  [7:0] I_2_2_1,
  input  [7:0] I_2_2_2,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_0_2,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_3_1_2,
  input  [7:0] I_3_2_0,
  input  [7:0] I_3_2_1,
  input  [7:0] I_3_2_2,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_0_2,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_4_1_2,
  input  [7:0] I_4_2_0,
  input  [7:0] I_4_2_1,
  input  [7:0] I_4_2_2,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_0_2,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_5_1_2,
  input  [7:0] I_5_2_0,
  input  [7:0] I_5_2_1,
  input  [7:0] I_5_2_2,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_0_2,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_6_1_2,
  input  [7:0] I_6_2_0,
  input  [7:0] I_6_2_1,
  input  [7:0] I_6_2_2,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_0_2,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_7_1_2,
  input  [7:0] I_7_2_0,
  input  [7:0] I_7_2_1,
  input  [7:0] I_7_2_2,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_0_2,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_8_1_2,
  input  [7:0] I_8_2_0,
  input  [7:0] I_8_2_1,
  input  [7:0] I_8_2_2,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_0_2,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_9_1_2,
  input  [7:0] I_9_2_0,
  input  [7:0] I_9_2_1,
  input  [7:0] I_9_2_2,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_0_2,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_10_1_2,
  input  [7:0] I_10_2_0,
  input  [7:0] I_10_2_1,
  input  [7:0] I_10_2_2,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_0_2,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_11_1_2,
  input  [7:0] I_11_2_0,
  input  [7:0] I_11_2_1,
  input  [7:0] I_11_2_2,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_0_2,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_12_1_2,
  input  [7:0] I_12_2_0,
  input  [7:0] I_12_2_1,
  input  [7:0] I_12_2_2,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_0_2,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_13_1_2,
  input  [7:0] I_13_2_0,
  input  [7:0] I_13_2_1,
  input  [7:0] I_13_2_2,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_0_2,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_14_1_2,
  input  [7:0] I_14_2_0,
  input  [7:0] I_14_2_1,
  input  [7:0] I_14_2_2,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_0_2,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  input  [7:0] I_15_1_2,
  input  [7:0] I_15_2_0,
  input  [7:0] I_15_2_1,
  input  [7:0] I_15_2_2,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_2; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_2_2; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  MapS_9 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_0_2(op_I_0_0_2),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_0_1_2(op_I_0_1_2),
    .I_0_2_0(op_I_0_2_0),
    .I_0_2_1(op_I_0_2_1),
    .I_0_2_2(op_I_0_2_2),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_0_2(op_I_1_0_2),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_1_1_2(op_I_1_1_2),
    .I_1_2_0(op_I_1_2_0),
    .I_1_2_1(op_I_1_2_1),
    .I_1_2_2(op_I_1_2_2),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_0_2(op_I_2_0_2),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_2_1_2(op_I_2_1_2),
    .I_2_2_0(op_I_2_2_0),
    .I_2_2_1(op_I_2_2_1),
    .I_2_2_2(op_I_2_2_2),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_0_2(op_I_3_0_2),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_3_1_2(op_I_3_1_2),
    .I_3_2_0(op_I_3_2_0),
    .I_3_2_1(op_I_3_2_1),
    .I_3_2_2(op_I_3_2_2),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_0_2(op_I_4_0_2),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_4_1_2(op_I_4_1_2),
    .I_4_2_0(op_I_4_2_0),
    .I_4_2_1(op_I_4_2_1),
    .I_4_2_2(op_I_4_2_2),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_0_2(op_I_5_0_2),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_5_1_2(op_I_5_1_2),
    .I_5_2_0(op_I_5_2_0),
    .I_5_2_1(op_I_5_2_1),
    .I_5_2_2(op_I_5_2_2),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_0_2(op_I_6_0_2),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_6_1_2(op_I_6_1_2),
    .I_6_2_0(op_I_6_2_0),
    .I_6_2_1(op_I_6_2_1),
    .I_6_2_2(op_I_6_2_2),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_0_2(op_I_7_0_2),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_7_1_2(op_I_7_1_2),
    .I_7_2_0(op_I_7_2_0),
    .I_7_2_1(op_I_7_2_1),
    .I_7_2_2(op_I_7_2_2),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_0_2(op_I_8_0_2),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_8_1_2(op_I_8_1_2),
    .I_8_2_0(op_I_8_2_0),
    .I_8_2_1(op_I_8_2_1),
    .I_8_2_2(op_I_8_2_2),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_0_2(op_I_9_0_2),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_9_1_2(op_I_9_1_2),
    .I_9_2_0(op_I_9_2_0),
    .I_9_2_1(op_I_9_2_1),
    .I_9_2_2(op_I_9_2_2),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_0_2(op_I_10_0_2),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_10_1_2(op_I_10_1_2),
    .I_10_2_0(op_I_10_2_0),
    .I_10_2_1(op_I_10_2_1),
    .I_10_2_2(op_I_10_2_2),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_0_2(op_I_11_0_2),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_11_1_2(op_I_11_1_2),
    .I_11_2_0(op_I_11_2_0),
    .I_11_2_1(op_I_11_2_1),
    .I_11_2_2(op_I_11_2_2),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_0_2(op_I_12_0_2),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_12_1_2(op_I_12_1_2),
    .I_12_2_0(op_I_12_2_0),
    .I_12_2_1(op_I_12_2_1),
    .I_12_2_2(op_I_12_2_2),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_0_2(op_I_13_0_2),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_13_1_2(op_I_13_1_2),
    .I_13_2_0(op_I_13_2_0),
    .I_13_2_1(op_I_13_2_1),
    .I_13_2_2(op_I_13_2_2),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_0_2(op_I_14_0_2),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_14_1_2(op_I_14_1_2),
    .I_14_2_0(op_I_14_2_0),
    .I_14_2_1(op_I_14_2_1),
    .I_14_2_2(op_I_14_2_2),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_0_2(op_I_15_0_2),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .I_15_1_2(op_I_15_1_2),
    .I_15_2_0(op_I_15_2_0),
    .I_15_2_1(op_I_15_2_1),
    .I_15_2_2(op_I_15_2_2),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0),
    .O_8_0_0(op_O_8_0_0),
    .O_9_0_0(op_O_9_0_0),
    .O_10_0_0(op_O_10_0_0),
    .O_11_0_0(op_O_11_0_0),
    .O_12_0_0(op_O_12_0_0),
    .O_13_0_0(op_O_13_0_0),
    .O_14_0_0(op_O_14_0_0),
    .O_15_0_0(op_O_15_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_2 = I_0_0_2; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_0_1_2 = I_0_1_2; // @[MapT.scala 14:10]
  assign op_I_0_2_0 = I_0_2_0; // @[MapT.scala 14:10]
  assign op_I_0_2_1 = I_0_2_1; // @[MapT.scala 14:10]
  assign op_I_0_2_2 = I_0_2_2; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_2 = I_1_0_2; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_1_1_2 = I_1_1_2; // @[MapT.scala 14:10]
  assign op_I_1_2_0 = I_1_2_0; // @[MapT.scala 14:10]
  assign op_I_1_2_1 = I_1_2_1; // @[MapT.scala 14:10]
  assign op_I_1_2_2 = I_1_2_2; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_2 = I_2_0_2; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_2_1_2 = I_2_1_2; // @[MapT.scala 14:10]
  assign op_I_2_2_0 = I_2_2_0; // @[MapT.scala 14:10]
  assign op_I_2_2_1 = I_2_2_1; // @[MapT.scala 14:10]
  assign op_I_2_2_2 = I_2_2_2; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_2 = I_3_0_2; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_3_1_2 = I_3_1_2; // @[MapT.scala 14:10]
  assign op_I_3_2_0 = I_3_2_0; // @[MapT.scala 14:10]
  assign op_I_3_2_1 = I_3_2_1; // @[MapT.scala 14:10]
  assign op_I_3_2_2 = I_3_2_2; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_2 = I_4_0_2; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_4_1_2 = I_4_1_2; // @[MapT.scala 14:10]
  assign op_I_4_2_0 = I_4_2_0; // @[MapT.scala 14:10]
  assign op_I_4_2_1 = I_4_2_1; // @[MapT.scala 14:10]
  assign op_I_4_2_2 = I_4_2_2; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_2 = I_5_0_2; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_5_1_2 = I_5_1_2; // @[MapT.scala 14:10]
  assign op_I_5_2_0 = I_5_2_0; // @[MapT.scala 14:10]
  assign op_I_5_2_1 = I_5_2_1; // @[MapT.scala 14:10]
  assign op_I_5_2_2 = I_5_2_2; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_2 = I_6_0_2; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_6_1_2 = I_6_1_2; // @[MapT.scala 14:10]
  assign op_I_6_2_0 = I_6_2_0; // @[MapT.scala 14:10]
  assign op_I_6_2_1 = I_6_2_1; // @[MapT.scala 14:10]
  assign op_I_6_2_2 = I_6_2_2; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_2 = I_7_0_2; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_7_1_2 = I_7_1_2; // @[MapT.scala 14:10]
  assign op_I_7_2_0 = I_7_2_0; // @[MapT.scala 14:10]
  assign op_I_7_2_1 = I_7_2_1; // @[MapT.scala 14:10]
  assign op_I_7_2_2 = I_7_2_2; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_2 = I_8_0_2; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_8_1_2 = I_8_1_2; // @[MapT.scala 14:10]
  assign op_I_8_2_0 = I_8_2_0; // @[MapT.scala 14:10]
  assign op_I_8_2_1 = I_8_2_1; // @[MapT.scala 14:10]
  assign op_I_8_2_2 = I_8_2_2; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_2 = I_9_0_2; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_9_1_2 = I_9_1_2; // @[MapT.scala 14:10]
  assign op_I_9_2_0 = I_9_2_0; // @[MapT.scala 14:10]
  assign op_I_9_2_1 = I_9_2_1; // @[MapT.scala 14:10]
  assign op_I_9_2_2 = I_9_2_2; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_2 = I_10_0_2; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_10_1_2 = I_10_1_2; // @[MapT.scala 14:10]
  assign op_I_10_2_0 = I_10_2_0; // @[MapT.scala 14:10]
  assign op_I_10_2_1 = I_10_2_1; // @[MapT.scala 14:10]
  assign op_I_10_2_2 = I_10_2_2; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_2 = I_11_0_2; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_11_1_2 = I_11_1_2; // @[MapT.scala 14:10]
  assign op_I_11_2_0 = I_11_2_0; // @[MapT.scala 14:10]
  assign op_I_11_2_1 = I_11_2_1; // @[MapT.scala 14:10]
  assign op_I_11_2_2 = I_11_2_2; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_2 = I_12_0_2; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_12_1_2 = I_12_1_2; // @[MapT.scala 14:10]
  assign op_I_12_2_0 = I_12_2_0; // @[MapT.scala 14:10]
  assign op_I_12_2_1 = I_12_2_1; // @[MapT.scala 14:10]
  assign op_I_12_2_2 = I_12_2_2; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_2 = I_13_0_2; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_13_1_2 = I_13_1_2; // @[MapT.scala 14:10]
  assign op_I_13_2_0 = I_13_2_0; // @[MapT.scala 14:10]
  assign op_I_13_2_1 = I_13_2_1; // @[MapT.scala 14:10]
  assign op_I_13_2_2 = I_13_2_2; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_2 = I_14_0_2; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_14_1_2 = I_14_1_2; // @[MapT.scala 14:10]
  assign op_I_14_2_0 = I_14_2_0; // @[MapT.scala 14:10]
  assign op_I_14_2_1 = I_14_2_1; // @[MapT.scala 14:10]
  assign op_I_14_2_2 = I_14_2_2; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_2 = I_15_0_2; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
  assign op_I_15_1_2 = I_15_1_2; // @[MapT.scala 14:10]
  assign op_I_15_2_0 = I_15_2_0; // @[MapT.scala 14:10]
  assign op_I_15_2_1 = I_15_2_1; // @[MapT.scala 14:10]
  assign op_I_15_2_2 = I_15_2_2; // @[MapT.scala 14:10]
endmodule
module Passthrough(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_1_0_0,
  input  [7:0] I_2_0_0,
  input  [7:0] I_3_0_0,
  input  [7:0] I_4_0_0,
  input  [7:0] I_5_0_0,
  input  [7:0] I_6_0_0,
  input  [7:0] I_7_0_0,
  input  [7:0] I_8_0_0,
  input  [7:0] I_9_0_0,
  input  [7:0] I_10_0_0,
  input  [7:0] I_11_0_0,
  input  [7:0] I_12_0_0,
  input  [7:0] I_13_0_0,
  input  [7:0] I_14_0_0,
  input  [7:0] I_15_0_0,
  output [7:0] O_0_0,
  output [7:0] O_1_0,
  output [7:0] O_2_0,
  output [7:0] O_3_0,
  output [7:0] O_4_0,
  output [7:0] O_5_0,
  output [7:0] O_6_0,
  output [7:0] O_7_0,
  output [7:0] O_8_0,
  output [7:0] O_9_0,
  output [7:0] O_10_0,
  output [7:0] O_11_0,
  output [7:0] O_12_0,
  output [7:0] O_13_0,
  output [7:0] O_14_0,
  output [7:0] O_15_0
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0_0 = I_0_0_0; // @[Passthrough.scala 17:68]
  assign O_1_0 = I_1_0_0; // @[Passthrough.scala 17:68]
  assign O_2_0 = I_2_0_0; // @[Passthrough.scala 17:68]
  assign O_3_0 = I_3_0_0; // @[Passthrough.scala 17:68]
  assign O_4_0 = I_4_0_0; // @[Passthrough.scala 17:68]
  assign O_5_0 = I_5_0_0; // @[Passthrough.scala 17:68]
  assign O_6_0 = I_6_0_0; // @[Passthrough.scala 17:68]
  assign O_7_0 = I_7_0_0; // @[Passthrough.scala 17:68]
  assign O_8_0 = I_8_0_0; // @[Passthrough.scala 17:68]
  assign O_9_0 = I_9_0_0; // @[Passthrough.scala 17:68]
  assign O_10_0 = I_10_0_0; // @[Passthrough.scala 17:68]
  assign O_11_0 = I_11_0_0; // @[Passthrough.scala 17:68]
  assign O_12_0 = I_12_0_0; // @[Passthrough.scala 17:68]
  assign O_13_0 = I_13_0_0; // @[Passthrough.scala 17:68]
  assign O_14_0 = I_14_0_0; // @[Passthrough.scala 17:68]
  assign O_15_0 = I_15_0_0; // @[Passthrough.scala 17:68]
endmodule
module Passthrough_1(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  input  [7:0] I_2_0,
  input  [7:0] I_3_0,
  input  [7:0] I_4_0,
  input  [7:0] I_5_0,
  input  [7:0] I_6_0,
  input  [7:0] I_7_0,
  input  [7:0] I_8_0,
  input  [7:0] I_9_0,
  input  [7:0] I_10_0,
  input  [7:0] I_11_0,
  input  [7:0] I_12_0,
  input  [7:0] I_13_0,
  input  [7:0] I_14_0,
  input  [7:0] I_15_0,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  assign valid_down = valid_up; // @[Passthrough.scala 18:14]
  assign O_0 = I_0_0; // @[Passthrough.scala 17:68]
  assign O_1 = I_1_0; // @[Passthrough.scala 17:68]
  assign O_2 = I_2_0; // @[Passthrough.scala 17:68]
  assign O_3 = I_3_0; // @[Passthrough.scala 17:68]
  assign O_4 = I_4_0; // @[Passthrough.scala 17:68]
  assign O_5 = I_5_0; // @[Passthrough.scala 17:68]
  assign O_6 = I_6_0; // @[Passthrough.scala 17:68]
  assign O_7 = I_7_0; // @[Passthrough.scala 17:68]
  assign O_8 = I_8_0; // @[Passthrough.scala 17:68]
  assign O_9 = I_9_0; // @[Passthrough.scala 17:68]
  assign O_10 = I_10_0; // @[Passthrough.scala 17:68]
  assign O_11 = I_11_0; // @[Passthrough.scala 17:68]
  assign O_12 = I_12_0; // @[Passthrough.scala 17:68]
  assign O_13 = I_13_0; // @[Passthrough.scala 17:68]
  assign O_14 = I_14_0; // @[Passthrough.scala 17:68]
  assign O_15 = I_15_0; // @[Passthrough.scala 17:68]
endmodule
module PartitionS_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_3_0,
  input  [7:0] I_3_1,
  input  [7:0] I_4_0,
  input  [7:0] I_4_1,
  input  [7:0] I_5_0,
  input  [7:0] I_5_1,
  input  [7:0] I_6_0,
  input  [7:0] I_6_1,
  input  [7:0] I_7_0,
  input  [7:0] I_7_1,
  input  [7:0] I_8_0,
  input  [7:0] I_8_1,
  input  [7:0] I_9_0,
  input  [7:0] I_9_1,
  input  [7:0] I_10_0,
  input  [7:0] I_10_1,
  input  [7:0] I_11_0,
  input  [7:0] I_11_1,
  input  [7:0] I_12_0,
  input  [7:0] I_12_1,
  input  [7:0] I_13_0,
  input  [7:0] I_13_1,
  input  [7:0] I_14_0,
  input  [7:0] I_14_1,
  input  [7:0] I_15_0,
  input  [7:0] I_15_1,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0 = I_0_0; // @[Partition.scala 15:39]
  assign O_0_0_1 = I_0_1; // @[Partition.scala 15:39]
  assign O_1_0_0 = I_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1 = I_1_1; // @[Partition.scala 15:39]
  assign O_2_0_0 = I_2_0; // @[Partition.scala 15:39]
  assign O_2_0_1 = I_2_1; // @[Partition.scala 15:39]
  assign O_3_0_0 = I_3_0; // @[Partition.scala 15:39]
  assign O_3_0_1 = I_3_1; // @[Partition.scala 15:39]
  assign O_4_0_0 = I_4_0; // @[Partition.scala 15:39]
  assign O_4_0_1 = I_4_1; // @[Partition.scala 15:39]
  assign O_5_0_0 = I_5_0; // @[Partition.scala 15:39]
  assign O_5_0_1 = I_5_1; // @[Partition.scala 15:39]
  assign O_6_0_0 = I_6_0; // @[Partition.scala 15:39]
  assign O_6_0_1 = I_6_1; // @[Partition.scala 15:39]
  assign O_7_0_0 = I_7_0; // @[Partition.scala 15:39]
  assign O_7_0_1 = I_7_1; // @[Partition.scala 15:39]
  assign O_8_0_0 = I_8_0; // @[Partition.scala 15:39]
  assign O_8_0_1 = I_8_1; // @[Partition.scala 15:39]
  assign O_9_0_0 = I_9_0; // @[Partition.scala 15:39]
  assign O_9_0_1 = I_9_1; // @[Partition.scala 15:39]
  assign O_10_0_0 = I_10_0; // @[Partition.scala 15:39]
  assign O_10_0_1 = I_10_1; // @[Partition.scala 15:39]
  assign O_11_0_0 = I_11_0; // @[Partition.scala 15:39]
  assign O_11_0_1 = I_11_1; // @[Partition.scala 15:39]
  assign O_12_0_0 = I_12_0; // @[Partition.scala 15:39]
  assign O_12_0_1 = I_12_1; // @[Partition.scala 15:39]
  assign O_13_0_0 = I_13_0; // @[Partition.scala 15:39]
  assign O_13_0_1 = I_13_1; // @[Partition.scala 15:39]
  assign O_14_0_0 = I_14_0; // @[Partition.scala 15:39]
  assign O_14_0_1 = I_14_1; // @[Partition.scala 15:39]
  assign O_15_0_0 = I_15_0; // @[Partition.scala 15:39]
  assign O_15_0_1 = I_15_1; // @[Partition.scala 15:39]
endmodule
module MapT_9(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  input  [7:0] I_2_0,
  input  [7:0] I_2_1,
  input  [7:0] I_3_0,
  input  [7:0] I_3_1,
  input  [7:0] I_4_0,
  input  [7:0] I_4_1,
  input  [7:0] I_5_0,
  input  [7:0] I_5_1,
  input  [7:0] I_6_0,
  input  [7:0] I_6_1,
  input  [7:0] I_7_0,
  input  [7:0] I_7_1,
  input  [7:0] I_8_0,
  input  [7:0] I_8_1,
  input  [7:0] I_9_0,
  input  [7:0] I_9_1,
  input  [7:0] I_10_0,
  input  [7:0] I_10_1,
  input  [7:0] I_11_0,
  input  [7:0] I_11_1,
  input  [7:0] I_12_0,
  input  [7:0] I_12_1,
  input  [7:0] I_13_0,
  input  [7:0] I_13_1,
  input  [7:0] I_14_0,
  input  [7:0] I_14_1,
  input  [7:0] I_15_0,
  input  [7:0] I_15_1,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[MapT.scala 8:20]
  PartitionS_4 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0(op_I_0_0),
    .I_0_1(op_I_0_1),
    .I_1_0(op_I_1_0),
    .I_1_1(op_I_1_1),
    .I_2_0(op_I_2_0),
    .I_2_1(op_I_2_1),
    .I_3_0(op_I_3_0),
    .I_3_1(op_I_3_1),
    .I_4_0(op_I_4_0),
    .I_4_1(op_I_4_1),
    .I_5_0(op_I_5_0),
    .I_5_1(op_I_5_1),
    .I_6_0(op_I_6_0),
    .I_6_1(op_I_6_1),
    .I_7_0(op_I_7_0),
    .I_7_1(op_I_7_1),
    .I_8_0(op_I_8_0),
    .I_8_1(op_I_8_1),
    .I_9_0(op_I_9_0),
    .I_9_1(op_I_9_1),
    .I_10_0(op_I_10_0),
    .I_10_1(op_I_10_1),
    .I_11_0(op_I_11_0),
    .I_11_1(op_I_11_1),
    .I_12_0(op_I_12_0),
    .I_12_1(op_I_12_1),
    .I_13_0(op_I_13_0),
    .I_13_1(op_I_13_1),
    .I_14_0(op_I_14_0),
    .I_14_1(op_I_14_1),
    .I_15_0(op_I_15_0),
    .I_15_1(op_I_15_1),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0 = I_0_0; // @[MapT.scala 14:10]
  assign op_I_0_1 = I_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0 = I_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1 = I_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0 = I_2_0; // @[MapT.scala 14:10]
  assign op_I_2_1 = I_2_1; // @[MapT.scala 14:10]
  assign op_I_3_0 = I_3_0; // @[MapT.scala 14:10]
  assign op_I_3_1 = I_3_1; // @[MapT.scala 14:10]
  assign op_I_4_0 = I_4_0; // @[MapT.scala 14:10]
  assign op_I_4_1 = I_4_1; // @[MapT.scala 14:10]
  assign op_I_5_0 = I_5_0; // @[MapT.scala 14:10]
  assign op_I_5_1 = I_5_1; // @[MapT.scala 14:10]
  assign op_I_6_0 = I_6_0; // @[MapT.scala 14:10]
  assign op_I_6_1 = I_6_1; // @[MapT.scala 14:10]
  assign op_I_7_0 = I_7_0; // @[MapT.scala 14:10]
  assign op_I_7_1 = I_7_1; // @[MapT.scala 14:10]
  assign op_I_8_0 = I_8_0; // @[MapT.scala 14:10]
  assign op_I_8_1 = I_8_1; // @[MapT.scala 14:10]
  assign op_I_9_0 = I_9_0; // @[MapT.scala 14:10]
  assign op_I_9_1 = I_9_1; // @[MapT.scala 14:10]
  assign op_I_10_0 = I_10_0; // @[MapT.scala 14:10]
  assign op_I_10_1 = I_10_1; // @[MapT.scala 14:10]
  assign op_I_11_0 = I_11_0; // @[MapT.scala 14:10]
  assign op_I_11_1 = I_11_1; // @[MapT.scala 14:10]
  assign op_I_12_0 = I_12_0; // @[MapT.scala 14:10]
  assign op_I_12_1 = I_12_1; // @[MapT.scala 14:10]
  assign op_I_13_0 = I_13_0; // @[MapT.scala 14:10]
  assign op_I_13_1 = I_13_1; // @[MapT.scala 14:10]
  assign op_I_14_0 = I_14_0; // @[MapT.scala 14:10]
  assign op_I_14_1 = I_14_1; // @[MapT.scala 14:10]
  assign op_I_15_0 = I_15_0; // @[MapT.scala 14:10]
  assign op_I_15_1 = I_15_1; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0 = I_0; // @[Tuple.scala 41:5]
  assign O_1 = I_1; // @[Tuple.scala 41:5]
endmodule
module Remove1S_4(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_4 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0(op_inst_I_0),
    .I_1(op_inst_I_1),
    .O_0(op_inst_O_0),
    .O_1(op_inst_O_1)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0 = op_inst_O_0; // @[Remove1S.scala 14:5]
  assign O_1 = op_inst_O_1; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0 = I_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1 = I_0_1; // @[Remove1S.scala 13:13]
endmodule
module MapS_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_15_0,
  output [7:0] O_15_1
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S_4 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  Remove1S_4 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  Remove1S_4 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .O_0(other_ops_1_O_0),
    .O_1(other_ops_1_O_1)
  );
  Remove1S_4 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .O_0(other_ops_2_O_0),
    .O_1(other_ops_2_O_1)
  );
  Remove1S_4 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .O_0(other_ops_3_O_0),
    .O_1(other_ops_3_O_1)
  );
  Remove1S_4 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .O_0(other_ops_4_O_0),
    .O_1(other_ops_4_O_1)
  );
  Remove1S_4 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .O_0(other_ops_5_O_0),
    .O_1(other_ops_5_O_1)
  );
  Remove1S_4 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .O_0(other_ops_6_O_0),
    .O_1(other_ops_6_O_1)
  );
  Remove1S_4 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .O_0(other_ops_7_O_0),
    .O_1(other_ops_7_O_1)
  );
  Remove1S_4 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .O_0(other_ops_8_O_0),
    .O_1(other_ops_8_O_1)
  );
  Remove1S_4 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .O_0(other_ops_9_O_0),
    .O_1(other_ops_9_O_1)
  );
  Remove1S_4 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .O_0(other_ops_10_O_0),
    .O_1(other_ops_10_O_1)
  );
  Remove1S_4 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .O_0(other_ops_11_O_0),
    .O_1(other_ops_11_O_1)
  );
  Remove1S_4 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .O_0(other_ops_12_O_0),
    .O_1(other_ops_12_O_1)
  );
  Remove1S_4 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .O_0(other_ops_13_O_0),
    .O_1(other_ops_13_O_1)
  );
  Remove1S_4 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .O_0(other_ops_14_O_0),
    .O_1(other_ops_14_O_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign O_2_0 = other_ops_1_O_0; // @[MapS.scala 21:12]
  assign O_2_1 = other_ops_1_O_1; // @[MapS.scala 21:12]
  assign O_3_0 = other_ops_2_O_0; // @[MapS.scala 21:12]
  assign O_3_1 = other_ops_2_O_1; // @[MapS.scala 21:12]
  assign O_4_0 = other_ops_3_O_0; // @[MapS.scala 21:12]
  assign O_4_1 = other_ops_3_O_1; // @[MapS.scala 21:12]
  assign O_5_0 = other_ops_4_O_0; // @[MapS.scala 21:12]
  assign O_5_1 = other_ops_4_O_1; // @[MapS.scala 21:12]
  assign O_6_0 = other_ops_5_O_0; // @[MapS.scala 21:12]
  assign O_6_1 = other_ops_5_O_1; // @[MapS.scala 21:12]
  assign O_7_0 = other_ops_6_O_0; // @[MapS.scala 21:12]
  assign O_7_1 = other_ops_6_O_1; // @[MapS.scala 21:12]
  assign O_8_0 = other_ops_7_O_0; // @[MapS.scala 21:12]
  assign O_8_1 = other_ops_7_O_1; // @[MapS.scala 21:12]
  assign O_9_0 = other_ops_8_O_0; // @[MapS.scala 21:12]
  assign O_9_1 = other_ops_8_O_1; // @[MapS.scala 21:12]
  assign O_10_0 = other_ops_9_O_0; // @[MapS.scala 21:12]
  assign O_10_1 = other_ops_9_O_1; // @[MapS.scala 21:12]
  assign O_11_0 = other_ops_10_O_0; // @[MapS.scala 21:12]
  assign O_11_1 = other_ops_10_O_1; // @[MapS.scala 21:12]
  assign O_12_0 = other_ops_11_O_0; // @[MapS.scala 21:12]
  assign O_12_1 = other_ops_11_O_1; // @[MapS.scala 21:12]
  assign O_13_0 = other_ops_12_O_0; // @[MapS.scala 21:12]
  assign O_13_1 = other_ops_12_O_1; // @[MapS.scala 21:12]
  assign O_14_0 = other_ops_13_O_0; // @[MapS.scala 21:12]
  assign O_14_1 = other_ops_13_O_1; // @[MapS.scala 21:12]
  assign O_15_0 = other_ops_14_O_0; // @[MapS.scala 21:12]
  assign O_15_1 = other_ops_14_O_1; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
endmodule
module MapT_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1,
  output [7:0] O_2_0,
  output [7:0] O_2_1,
  output [7:0] O_3_0,
  output [7:0] O_3_1,
  output [7:0] O_4_0,
  output [7:0] O_4_1,
  output [7:0] O_5_0,
  output [7:0] O_5_1,
  output [7:0] O_6_0,
  output [7:0] O_6_1,
  output [7:0] O_7_0,
  output [7:0] O_7_1,
  output [7:0] O_8_0,
  output [7:0] O_8_1,
  output [7:0] O_9_0,
  output [7:0] O_9_1,
  output [7:0] O_10_0,
  output [7:0] O_10_1,
  output [7:0] O_11_0,
  output [7:0] O_11_1,
  output [7:0] O_12_0,
  output [7:0] O_12_1,
  output [7:0] O_13_0,
  output [7:0] O_13_1,
  output [7:0] O_14_0,
  output [7:0] O_14_1,
  output [7:0] O_15_0,
  output [7:0] O_15_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1; // @[MapT.scala 8:20]
  MapS_10 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .O_0_0(op_O_0_0),
    .O_0_1(op_O_0_1),
    .O_1_0(op_O_1_0),
    .O_1_1(op_O_1_1),
    .O_2_0(op_O_2_0),
    .O_2_1(op_O_2_1),
    .O_3_0(op_O_3_0),
    .O_3_1(op_O_3_1),
    .O_4_0(op_O_4_0),
    .O_4_1(op_O_4_1),
    .O_5_0(op_O_5_0),
    .O_5_1(op_O_5_1),
    .O_6_0(op_O_6_0),
    .O_6_1(op_O_6_1),
    .O_7_0(op_O_7_0),
    .O_7_1(op_O_7_1),
    .O_8_0(op_O_8_0),
    .O_8_1(op_O_8_1),
    .O_9_0(op_O_9_0),
    .O_9_1(op_O_9_1),
    .O_10_0(op_O_10_0),
    .O_10_1(op_O_10_1),
    .O_11_0(op_O_11_0),
    .O_11_1(op_O_11_1),
    .O_12_0(op_O_12_0),
    .O_12_1(op_O_12_1),
    .O_13_0(op_O_13_0),
    .O_13_1(op_O_13_1),
    .O_14_0(op_O_14_0),
    .O_14_1(op_O_14_1),
    .O_15_0(op_O_15_0),
    .O_15_1(op_O_15_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0 = op_O_0_0; // @[MapT.scala 15:7]
  assign O_0_1 = op_O_0_1; // @[MapT.scala 15:7]
  assign O_1_0 = op_O_1_0; // @[MapT.scala 15:7]
  assign O_1_1 = op_O_1_1; // @[MapT.scala 15:7]
  assign O_2_0 = op_O_2_0; // @[MapT.scala 15:7]
  assign O_2_1 = op_O_2_1; // @[MapT.scala 15:7]
  assign O_3_0 = op_O_3_0; // @[MapT.scala 15:7]
  assign O_3_1 = op_O_3_1; // @[MapT.scala 15:7]
  assign O_4_0 = op_O_4_0; // @[MapT.scala 15:7]
  assign O_4_1 = op_O_4_1; // @[MapT.scala 15:7]
  assign O_5_0 = op_O_5_0; // @[MapT.scala 15:7]
  assign O_5_1 = op_O_5_1; // @[MapT.scala 15:7]
  assign O_6_0 = op_O_6_0; // @[MapT.scala 15:7]
  assign O_6_1 = op_O_6_1; // @[MapT.scala 15:7]
  assign O_7_0 = op_O_7_0; // @[MapT.scala 15:7]
  assign O_7_1 = op_O_7_1; // @[MapT.scala 15:7]
  assign O_8_0 = op_O_8_0; // @[MapT.scala 15:7]
  assign O_8_1 = op_O_8_1; // @[MapT.scala 15:7]
  assign O_9_0 = op_O_9_0; // @[MapT.scala 15:7]
  assign O_9_1 = op_O_9_1; // @[MapT.scala 15:7]
  assign O_10_0 = op_O_10_0; // @[MapT.scala 15:7]
  assign O_10_1 = op_O_10_1; // @[MapT.scala 15:7]
  assign O_11_0 = op_O_11_0; // @[MapT.scala 15:7]
  assign O_11_1 = op_O_11_1; // @[MapT.scala 15:7]
  assign O_12_0 = op_O_12_0; // @[MapT.scala 15:7]
  assign O_12_1 = op_O_12_1; // @[MapT.scala 15:7]
  assign O_13_0 = op_O_13_0; // @[MapT.scala 15:7]
  assign O_13_1 = op_O_13_1; // @[MapT.scala 15:7]
  assign O_14_0 = op_O_14_0; // @[MapT.scala 15:7]
  assign O_14_1 = op_O_14_1; // @[MapT.scala 15:7]
  assign O_15_0 = op_O_15_0; // @[MapT.scala 15:7]
  assign O_15_1 = op_O_15_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
endmodule
module SSeqTupleCreator_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1
);
  assign valid_down = valid_up; // @[Tuple.scala 15:14]
  assign O_0_0 = I0_0; // @[Tuple.scala 12:32]
  assign O_0_1 = I0_1; // @[Tuple.scala 12:32]
  assign O_1_0 = I1_0; // @[Tuple.scala 13:32]
  assign O_1_1 = I1_1; // @[Tuple.scala 13:32]
endmodule
module Map2S_14(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_3_0,
  input  [7:0] I0_3_1,
  input  [7:0] I0_4_0,
  input  [7:0] I0_4_1,
  input  [7:0] I0_5_0,
  input  [7:0] I0_5_1,
  input  [7:0] I0_6_0,
  input  [7:0] I0_6_1,
  input  [7:0] I0_7_0,
  input  [7:0] I0_7_1,
  input  [7:0] I0_8_0,
  input  [7:0] I0_8_1,
  input  [7:0] I0_9_0,
  input  [7:0] I0_9_1,
  input  [7:0] I0_10_0,
  input  [7:0] I0_10_1,
  input  [7:0] I0_11_0,
  input  [7:0] I0_11_1,
  input  [7:0] I0_12_0,
  input  [7:0] I0_12_1,
  input  [7:0] I0_13_0,
  input  [7:0] I0_13_1,
  input  [7:0] I0_14_0,
  input  [7:0] I0_14_1,
  input  [7:0] I0_15_0,
  input  [7:0] I0_15_1,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_2_0,
  input  [7:0] I1_2_1,
  input  [7:0] I1_3_0,
  input  [7:0] I1_3_1,
  input  [7:0] I1_4_0,
  input  [7:0] I1_4_1,
  input  [7:0] I1_5_0,
  input  [7:0] I1_5_1,
  input  [7:0] I1_6_0,
  input  [7:0] I1_6_1,
  input  [7:0] I1_7_0,
  input  [7:0] I1_7_1,
  input  [7:0] I1_8_0,
  input  [7:0] I1_8_1,
  input  [7:0] I1_9_0,
  input  [7:0] I1_9_1,
  input  [7:0] I1_10_0,
  input  [7:0] I1_10_1,
  input  [7:0] I1_11_0,
  input  [7:0] I1_11_1,
  input  [7:0] I1_12_0,
  input  [7:0] I1_12_1,
  input  [7:0] I1_13_0,
  input  [7:0] I1_13_1,
  input  [7:0] I1_14_0,
  input  [7:0] I1_14_1,
  input  [7:0] I1_15_0,
  input  [7:0] I1_15_1,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_1_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_2_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_3_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_4_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_5_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_6_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_7_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_8_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_9_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_10_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_11_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_12_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_13_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_14_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[Map2S.scala 10:86]
  wire  _T; // @[Map2S.scala 26:83]
  wire  _T_1; // @[Map2S.scala 26:83]
  wire  _T_2; // @[Map2S.scala 26:83]
  wire  _T_3; // @[Map2S.scala 26:83]
  wire  _T_4; // @[Map2S.scala 26:83]
  wire  _T_5; // @[Map2S.scala 26:83]
  wire  _T_6; // @[Map2S.scala 26:83]
  wire  _T_7; // @[Map2S.scala 26:83]
  wire  _T_8; // @[Map2S.scala 26:83]
  wire  _T_9; // @[Map2S.scala 26:83]
  wire  _T_10; // @[Map2S.scala 26:83]
  wire  _T_11; // @[Map2S.scala 26:83]
  wire  _T_12; // @[Map2S.scala 26:83]
  wire  _T_13; // @[Map2S.scala 26:83]
  SSeqTupleCreator_6 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_1 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I0_0(other_ops_1_I0_0),
    .I0_1(other_ops_1_I0_1),
    .I1_0(other_ops_1_I1_0),
    .I1_1(other_ops_1_I1_1),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_2 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I0_0(other_ops_2_I0_0),
    .I0_1(other_ops_2_I0_1),
    .I1_0(other_ops_2_I1_0),
    .I1_1(other_ops_2_I1_1),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_3 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I0_0(other_ops_3_I0_0),
    .I0_1(other_ops_3_I0_1),
    .I1_0(other_ops_3_I1_0),
    .I1_1(other_ops_3_I1_1),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_4 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I0_0(other_ops_4_I0_0),
    .I0_1(other_ops_4_I0_1),
    .I1_0(other_ops_4_I1_0),
    .I1_1(other_ops_4_I1_1),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_5 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I0_0(other_ops_5_I0_0),
    .I0_1(other_ops_5_I0_1),
    .I1_0(other_ops_5_I1_0),
    .I1_1(other_ops_5_I1_1),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_6 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I0_0(other_ops_6_I0_0),
    .I0_1(other_ops_6_I0_1),
    .I1_0(other_ops_6_I1_0),
    .I1_1(other_ops_6_I1_1),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_7 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I0_0(other_ops_7_I0_0),
    .I0_1(other_ops_7_I0_1),
    .I1_0(other_ops_7_I1_0),
    .I1_1(other_ops_7_I1_1),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_8 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I0_0(other_ops_8_I0_0),
    .I0_1(other_ops_8_I0_1),
    .I1_0(other_ops_8_I1_0),
    .I1_1(other_ops_8_I1_1),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_9 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I0_0(other_ops_9_I0_0),
    .I0_1(other_ops_9_I0_1),
    .I1_0(other_ops_9_I1_0),
    .I1_1(other_ops_9_I1_1),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_10 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I0_0(other_ops_10_I0_0),
    .I0_1(other_ops_10_I0_1),
    .I1_0(other_ops_10_I1_0),
    .I1_1(other_ops_10_I1_1),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_11 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I0_0(other_ops_11_I0_0),
    .I0_1(other_ops_11_I0_1),
    .I1_0(other_ops_11_I1_0),
    .I1_1(other_ops_11_I1_1),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_12 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I0_0(other_ops_12_I0_0),
    .I0_1(other_ops_12_I0_1),
    .I1_0(other_ops_12_I1_0),
    .I1_1(other_ops_12_I1_1),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_13 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I0_0(other_ops_13_I0_0),
    .I0_1(other_ops_13_I0_1),
    .I1_0(other_ops_13_I1_0),
    .I1_1(other_ops_13_I1_1),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1)
  );
  SSeqTupleCreator_6 other_ops_14 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I0_0(other_ops_14_I0_0),
    .I0_1(other_ops_14_I0_1),
    .I1_0(other_ops_14_I1_0),
    .I1_1(other_ops_14_I1_1),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[Map2S.scala 26:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[Map2S.scala 26:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[Map2S.scala 26:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[Map2S.scala 26:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[Map2S.scala 26:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[Map2S.scala 26:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[Map2S.scala 26:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[Map2S.scala 26:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[Map2S.scala 26:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[Map2S.scala 26:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[Map2S.scala 26:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[Map2S.scala 26:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[Map2S.scala 26:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[Map2S.scala 19:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[Map2S.scala 19:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[Map2S.scala 19:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[Map2S.scala 19:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[Map2S.scala 24:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[Map2S.scala 24:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[Map2S.scala 24:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[Map2S.scala 24:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[Map2S.scala 24:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[Map2S.scala 24:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[Map2S.scala 24:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[Map2S.scala 24:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[Map2S.scala 24:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[Map2S.scala 24:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[Map2S.scala 24:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[Map2S.scala 24:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[Map2S.scala 24:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[Map2S.scala 24:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[Map2S.scala 24:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[Map2S.scala 24:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[Map2S.scala 24:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[Map2S.scala 24:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[Map2S.scala 24:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[Map2S.scala 24:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[Map2S.scala 24:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[Map2S.scala 24:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[Map2S.scala 24:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[Map2S.scala 24:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[Map2S.scala 24:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[Map2S.scala 24:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[Map2S.scala 24:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[Map2S.scala 24:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[Map2S.scala 24:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[Map2S.scala 24:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[Map2S.scala 24:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[Map2S.scala 24:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[Map2S.scala 24:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[Map2S.scala 24:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[Map2S.scala 24:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[Map2S.scala 24:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[Map2S.scala 24:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[Map2S.scala 24:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[Map2S.scala 24:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[Map2S.scala 24:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[Map2S.scala 24:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[Map2S.scala 24:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[Map2S.scala 24:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[Map2S.scala 24:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[Map2S.scala 24:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[Map2S.scala 24:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[Map2S.scala 24:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[Map2S.scala 24:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[Map2S.scala 24:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[Map2S.scala 24:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[Map2S.scala 24:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[Map2S.scala 24:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[Map2S.scala 24:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[Map2S.scala 24:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[Map2S.scala 24:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[Map2S.scala 24:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[Map2S.scala 24:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[Map2S.scala 24:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[Map2S.scala 24:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = I1_0_0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = I1_0_1; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = I1_1_0; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = I1_1_1; // @[Map2S.scala 23:43]
  assign other_ops_1_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_1_I0_0 = I0_2_0; // @[Map2S.scala 22:43]
  assign other_ops_1_I0_1 = I0_2_1; // @[Map2S.scala 22:43]
  assign other_ops_1_I1_0 = I1_2_0; // @[Map2S.scala 23:43]
  assign other_ops_1_I1_1 = I1_2_1; // @[Map2S.scala 23:43]
  assign other_ops_2_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_2_I0_0 = I0_3_0; // @[Map2S.scala 22:43]
  assign other_ops_2_I0_1 = I0_3_1; // @[Map2S.scala 22:43]
  assign other_ops_2_I1_0 = I1_3_0; // @[Map2S.scala 23:43]
  assign other_ops_2_I1_1 = I1_3_1; // @[Map2S.scala 23:43]
  assign other_ops_3_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_3_I0_0 = I0_4_0; // @[Map2S.scala 22:43]
  assign other_ops_3_I0_1 = I0_4_1; // @[Map2S.scala 22:43]
  assign other_ops_3_I1_0 = I1_4_0; // @[Map2S.scala 23:43]
  assign other_ops_3_I1_1 = I1_4_1; // @[Map2S.scala 23:43]
  assign other_ops_4_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_4_I0_0 = I0_5_0; // @[Map2S.scala 22:43]
  assign other_ops_4_I0_1 = I0_5_1; // @[Map2S.scala 22:43]
  assign other_ops_4_I1_0 = I1_5_0; // @[Map2S.scala 23:43]
  assign other_ops_4_I1_1 = I1_5_1; // @[Map2S.scala 23:43]
  assign other_ops_5_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_5_I0_0 = I0_6_0; // @[Map2S.scala 22:43]
  assign other_ops_5_I0_1 = I0_6_1; // @[Map2S.scala 22:43]
  assign other_ops_5_I1_0 = I1_6_0; // @[Map2S.scala 23:43]
  assign other_ops_5_I1_1 = I1_6_1; // @[Map2S.scala 23:43]
  assign other_ops_6_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_6_I0_0 = I0_7_0; // @[Map2S.scala 22:43]
  assign other_ops_6_I0_1 = I0_7_1; // @[Map2S.scala 22:43]
  assign other_ops_6_I1_0 = I1_7_0; // @[Map2S.scala 23:43]
  assign other_ops_6_I1_1 = I1_7_1; // @[Map2S.scala 23:43]
  assign other_ops_7_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_7_I0_0 = I0_8_0; // @[Map2S.scala 22:43]
  assign other_ops_7_I0_1 = I0_8_1; // @[Map2S.scala 22:43]
  assign other_ops_7_I1_0 = I1_8_0; // @[Map2S.scala 23:43]
  assign other_ops_7_I1_1 = I1_8_1; // @[Map2S.scala 23:43]
  assign other_ops_8_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_8_I0_0 = I0_9_0; // @[Map2S.scala 22:43]
  assign other_ops_8_I0_1 = I0_9_1; // @[Map2S.scala 22:43]
  assign other_ops_8_I1_0 = I1_9_0; // @[Map2S.scala 23:43]
  assign other_ops_8_I1_1 = I1_9_1; // @[Map2S.scala 23:43]
  assign other_ops_9_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_9_I0_0 = I0_10_0; // @[Map2S.scala 22:43]
  assign other_ops_9_I0_1 = I0_10_1; // @[Map2S.scala 22:43]
  assign other_ops_9_I1_0 = I1_10_0; // @[Map2S.scala 23:43]
  assign other_ops_9_I1_1 = I1_10_1; // @[Map2S.scala 23:43]
  assign other_ops_10_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_10_I0_0 = I0_11_0; // @[Map2S.scala 22:43]
  assign other_ops_10_I0_1 = I0_11_1; // @[Map2S.scala 22:43]
  assign other_ops_10_I1_0 = I1_11_0; // @[Map2S.scala 23:43]
  assign other_ops_10_I1_1 = I1_11_1; // @[Map2S.scala 23:43]
  assign other_ops_11_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_11_I0_0 = I0_12_0; // @[Map2S.scala 22:43]
  assign other_ops_11_I0_1 = I0_12_1; // @[Map2S.scala 22:43]
  assign other_ops_11_I1_0 = I1_12_0; // @[Map2S.scala 23:43]
  assign other_ops_11_I1_1 = I1_12_1; // @[Map2S.scala 23:43]
  assign other_ops_12_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_12_I0_0 = I0_13_0; // @[Map2S.scala 22:43]
  assign other_ops_12_I0_1 = I0_13_1; // @[Map2S.scala 22:43]
  assign other_ops_12_I1_0 = I1_13_0; // @[Map2S.scala 23:43]
  assign other_ops_12_I1_1 = I1_13_1; // @[Map2S.scala 23:43]
  assign other_ops_13_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_13_I0_0 = I0_14_0; // @[Map2S.scala 22:43]
  assign other_ops_13_I0_1 = I0_14_1; // @[Map2S.scala 22:43]
  assign other_ops_13_I1_0 = I1_14_0; // @[Map2S.scala 23:43]
  assign other_ops_13_I1_1 = I1_14_1; // @[Map2S.scala 23:43]
  assign other_ops_14_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_14_I0_0 = I0_15_0; // @[Map2S.scala 22:43]
  assign other_ops_14_I0_1 = I0_15_1; // @[Map2S.scala 22:43]
  assign other_ops_14_I1_0 = I1_15_0; // @[Map2S.scala 23:43]
  assign other_ops_14_I1_1 = I1_15_1; // @[Map2S.scala 23:43]
endmodule
module Map2T_10(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  input  [7:0] I0_2_0,
  input  [7:0] I0_2_1,
  input  [7:0] I0_3_0,
  input  [7:0] I0_3_1,
  input  [7:0] I0_4_0,
  input  [7:0] I0_4_1,
  input  [7:0] I0_5_0,
  input  [7:0] I0_5_1,
  input  [7:0] I0_6_0,
  input  [7:0] I0_6_1,
  input  [7:0] I0_7_0,
  input  [7:0] I0_7_1,
  input  [7:0] I0_8_0,
  input  [7:0] I0_8_1,
  input  [7:0] I0_9_0,
  input  [7:0] I0_9_1,
  input  [7:0] I0_10_0,
  input  [7:0] I0_10_1,
  input  [7:0] I0_11_0,
  input  [7:0] I0_11_1,
  input  [7:0] I0_12_0,
  input  [7:0] I0_12_1,
  input  [7:0] I0_13_0,
  input  [7:0] I0_13_1,
  input  [7:0] I0_14_0,
  input  [7:0] I0_14_1,
  input  [7:0] I0_15_0,
  input  [7:0] I0_15_1,
  input  [7:0] I1_0_0,
  input  [7:0] I1_0_1,
  input  [7:0] I1_1_0,
  input  [7:0] I1_1_1,
  input  [7:0] I1_2_0,
  input  [7:0] I1_2_1,
  input  [7:0] I1_3_0,
  input  [7:0] I1_3_1,
  input  [7:0] I1_4_0,
  input  [7:0] I1_4_1,
  input  [7:0] I1_5_0,
  input  [7:0] I1_5_1,
  input  [7:0] I1_6_0,
  input  [7:0] I1_6_1,
  input  [7:0] I1_7_0,
  input  [7:0] I1_7_1,
  input  [7:0] I1_8_0,
  input  [7:0] I1_8_1,
  input  [7:0] I1_9_0,
  input  [7:0] I1_9_1,
  input  [7:0] I1_10_0,
  input  [7:0] I1_10_1,
  input  [7:0] I1_11_0,
  input  [7:0] I1_11_1,
  input  [7:0] I1_12_0,
  input  [7:0] I1_12_1,
  input  [7:0] I1_13_0,
  input  [7:0] I1_13_1,
  input  [7:0] I1_14_0,
  input  [7:0] I1_14_1,
  input  [7:0] I1_15_0,
  input  [7:0] I1_15_1,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1
);
  wire  op_valid_up; // @[Map2T.scala 8:20]
  wire  op_valid_down; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_3_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_4_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_5_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_6_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_7_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_8_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_9_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_10_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_11_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_12_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_13_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_14_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I0_15_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_2_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_3_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_4_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_5_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_6_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_7_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_8_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_9_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_10_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_11_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_12_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_13_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_14_1; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_0; // @[Map2T.scala 8:20]
  wire [7:0] op_I1_15_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_2_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_3_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_4_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_5_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_6_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_7_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_8_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_9_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_10_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_11_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_12_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_13_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_14_1_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1_0; // @[Map2T.scala 8:20]
  wire [7:0] op_O_15_1_1; // @[Map2T.scala 8:20]
  Map2S_14 op ( // @[Map2T.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I0_0_0(op_I0_0_0),
    .I0_0_1(op_I0_0_1),
    .I0_1_0(op_I0_1_0),
    .I0_1_1(op_I0_1_1),
    .I0_2_0(op_I0_2_0),
    .I0_2_1(op_I0_2_1),
    .I0_3_0(op_I0_3_0),
    .I0_3_1(op_I0_3_1),
    .I0_4_0(op_I0_4_0),
    .I0_4_1(op_I0_4_1),
    .I0_5_0(op_I0_5_0),
    .I0_5_1(op_I0_5_1),
    .I0_6_0(op_I0_6_0),
    .I0_6_1(op_I0_6_1),
    .I0_7_0(op_I0_7_0),
    .I0_7_1(op_I0_7_1),
    .I0_8_0(op_I0_8_0),
    .I0_8_1(op_I0_8_1),
    .I0_9_0(op_I0_9_0),
    .I0_9_1(op_I0_9_1),
    .I0_10_0(op_I0_10_0),
    .I0_10_1(op_I0_10_1),
    .I0_11_0(op_I0_11_0),
    .I0_11_1(op_I0_11_1),
    .I0_12_0(op_I0_12_0),
    .I0_12_1(op_I0_12_1),
    .I0_13_0(op_I0_13_0),
    .I0_13_1(op_I0_13_1),
    .I0_14_0(op_I0_14_0),
    .I0_14_1(op_I0_14_1),
    .I0_15_0(op_I0_15_0),
    .I0_15_1(op_I0_15_1),
    .I1_0_0(op_I1_0_0),
    .I1_0_1(op_I1_0_1),
    .I1_1_0(op_I1_1_0),
    .I1_1_1(op_I1_1_1),
    .I1_2_0(op_I1_2_0),
    .I1_2_1(op_I1_2_1),
    .I1_3_0(op_I1_3_0),
    .I1_3_1(op_I1_3_1),
    .I1_4_0(op_I1_4_0),
    .I1_4_1(op_I1_4_1),
    .I1_5_0(op_I1_5_0),
    .I1_5_1(op_I1_5_1),
    .I1_6_0(op_I1_6_0),
    .I1_6_1(op_I1_6_1),
    .I1_7_0(op_I1_7_0),
    .I1_7_1(op_I1_7_1),
    .I1_8_0(op_I1_8_0),
    .I1_8_1(op_I1_8_1),
    .I1_9_0(op_I1_9_0),
    .I1_9_1(op_I1_9_1),
    .I1_10_0(op_I1_10_0),
    .I1_10_1(op_I1_10_1),
    .I1_11_0(op_I1_11_0),
    .I1_11_1(op_I1_11_1),
    .I1_12_0(op_I1_12_0),
    .I1_12_1(op_I1_12_1),
    .I1_13_0(op_I1_13_0),
    .I1_13_1(op_I1_13_1),
    .I1_14_0(op_I1_14_0),
    .I1_14_1(op_I1_14_1),
    .I1_15_0(op_I1_15_0),
    .I1_15_1(op_I1_15_1),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1)
  );
  assign valid_down = op_valid_down; // @[Map2T.scala 18:16]
  assign O_0_0_0 = op_O_0_0_0; // @[Map2T.scala 17:7]
  assign O_0_0_1 = op_O_0_0_1; // @[Map2T.scala 17:7]
  assign O_0_1_0 = op_O_0_1_0; // @[Map2T.scala 17:7]
  assign O_0_1_1 = op_O_0_1_1; // @[Map2T.scala 17:7]
  assign O_1_0_0 = op_O_1_0_0; // @[Map2T.scala 17:7]
  assign O_1_0_1 = op_O_1_0_1; // @[Map2T.scala 17:7]
  assign O_1_1_0 = op_O_1_1_0; // @[Map2T.scala 17:7]
  assign O_1_1_1 = op_O_1_1_1; // @[Map2T.scala 17:7]
  assign O_2_0_0 = op_O_2_0_0; // @[Map2T.scala 17:7]
  assign O_2_0_1 = op_O_2_0_1; // @[Map2T.scala 17:7]
  assign O_2_1_0 = op_O_2_1_0; // @[Map2T.scala 17:7]
  assign O_2_1_1 = op_O_2_1_1; // @[Map2T.scala 17:7]
  assign O_3_0_0 = op_O_3_0_0; // @[Map2T.scala 17:7]
  assign O_3_0_1 = op_O_3_0_1; // @[Map2T.scala 17:7]
  assign O_3_1_0 = op_O_3_1_0; // @[Map2T.scala 17:7]
  assign O_3_1_1 = op_O_3_1_1; // @[Map2T.scala 17:7]
  assign O_4_0_0 = op_O_4_0_0; // @[Map2T.scala 17:7]
  assign O_4_0_1 = op_O_4_0_1; // @[Map2T.scala 17:7]
  assign O_4_1_0 = op_O_4_1_0; // @[Map2T.scala 17:7]
  assign O_4_1_1 = op_O_4_1_1; // @[Map2T.scala 17:7]
  assign O_5_0_0 = op_O_5_0_0; // @[Map2T.scala 17:7]
  assign O_5_0_1 = op_O_5_0_1; // @[Map2T.scala 17:7]
  assign O_5_1_0 = op_O_5_1_0; // @[Map2T.scala 17:7]
  assign O_5_1_1 = op_O_5_1_1; // @[Map2T.scala 17:7]
  assign O_6_0_0 = op_O_6_0_0; // @[Map2T.scala 17:7]
  assign O_6_0_1 = op_O_6_0_1; // @[Map2T.scala 17:7]
  assign O_6_1_0 = op_O_6_1_0; // @[Map2T.scala 17:7]
  assign O_6_1_1 = op_O_6_1_1; // @[Map2T.scala 17:7]
  assign O_7_0_0 = op_O_7_0_0; // @[Map2T.scala 17:7]
  assign O_7_0_1 = op_O_7_0_1; // @[Map2T.scala 17:7]
  assign O_7_1_0 = op_O_7_1_0; // @[Map2T.scala 17:7]
  assign O_7_1_1 = op_O_7_1_1; // @[Map2T.scala 17:7]
  assign O_8_0_0 = op_O_8_0_0; // @[Map2T.scala 17:7]
  assign O_8_0_1 = op_O_8_0_1; // @[Map2T.scala 17:7]
  assign O_8_1_0 = op_O_8_1_0; // @[Map2T.scala 17:7]
  assign O_8_1_1 = op_O_8_1_1; // @[Map2T.scala 17:7]
  assign O_9_0_0 = op_O_9_0_0; // @[Map2T.scala 17:7]
  assign O_9_0_1 = op_O_9_0_1; // @[Map2T.scala 17:7]
  assign O_9_1_0 = op_O_9_1_0; // @[Map2T.scala 17:7]
  assign O_9_1_1 = op_O_9_1_1; // @[Map2T.scala 17:7]
  assign O_10_0_0 = op_O_10_0_0; // @[Map2T.scala 17:7]
  assign O_10_0_1 = op_O_10_0_1; // @[Map2T.scala 17:7]
  assign O_10_1_0 = op_O_10_1_0; // @[Map2T.scala 17:7]
  assign O_10_1_1 = op_O_10_1_1; // @[Map2T.scala 17:7]
  assign O_11_0_0 = op_O_11_0_0; // @[Map2T.scala 17:7]
  assign O_11_0_1 = op_O_11_0_1; // @[Map2T.scala 17:7]
  assign O_11_1_0 = op_O_11_1_0; // @[Map2T.scala 17:7]
  assign O_11_1_1 = op_O_11_1_1; // @[Map2T.scala 17:7]
  assign O_12_0_0 = op_O_12_0_0; // @[Map2T.scala 17:7]
  assign O_12_0_1 = op_O_12_0_1; // @[Map2T.scala 17:7]
  assign O_12_1_0 = op_O_12_1_0; // @[Map2T.scala 17:7]
  assign O_12_1_1 = op_O_12_1_1; // @[Map2T.scala 17:7]
  assign O_13_0_0 = op_O_13_0_0; // @[Map2T.scala 17:7]
  assign O_13_0_1 = op_O_13_0_1; // @[Map2T.scala 17:7]
  assign O_13_1_0 = op_O_13_1_0; // @[Map2T.scala 17:7]
  assign O_13_1_1 = op_O_13_1_1; // @[Map2T.scala 17:7]
  assign O_14_0_0 = op_O_14_0_0; // @[Map2T.scala 17:7]
  assign O_14_0_1 = op_O_14_0_1; // @[Map2T.scala 17:7]
  assign O_14_1_0 = op_O_14_1_0; // @[Map2T.scala 17:7]
  assign O_14_1_1 = op_O_14_1_1; // @[Map2T.scala 17:7]
  assign O_15_0_0 = op_O_15_0_0; // @[Map2T.scala 17:7]
  assign O_15_0_1 = op_O_15_0_1; // @[Map2T.scala 17:7]
  assign O_15_1_0 = op_O_15_1_0; // @[Map2T.scala 17:7]
  assign O_15_1_1 = op_O_15_1_1; // @[Map2T.scala 17:7]
  assign op_valid_up = valid_up; // @[Map2T.scala 14:17]
  assign op_I0_0_0 = I0_0_0; // @[Map2T.scala 15:11]
  assign op_I0_0_1 = I0_0_1; // @[Map2T.scala 15:11]
  assign op_I0_1_0 = I0_1_0; // @[Map2T.scala 15:11]
  assign op_I0_1_1 = I0_1_1; // @[Map2T.scala 15:11]
  assign op_I0_2_0 = I0_2_0; // @[Map2T.scala 15:11]
  assign op_I0_2_1 = I0_2_1; // @[Map2T.scala 15:11]
  assign op_I0_3_0 = I0_3_0; // @[Map2T.scala 15:11]
  assign op_I0_3_1 = I0_3_1; // @[Map2T.scala 15:11]
  assign op_I0_4_0 = I0_4_0; // @[Map2T.scala 15:11]
  assign op_I0_4_1 = I0_4_1; // @[Map2T.scala 15:11]
  assign op_I0_5_0 = I0_5_0; // @[Map2T.scala 15:11]
  assign op_I0_5_1 = I0_5_1; // @[Map2T.scala 15:11]
  assign op_I0_6_0 = I0_6_0; // @[Map2T.scala 15:11]
  assign op_I0_6_1 = I0_6_1; // @[Map2T.scala 15:11]
  assign op_I0_7_0 = I0_7_0; // @[Map2T.scala 15:11]
  assign op_I0_7_1 = I0_7_1; // @[Map2T.scala 15:11]
  assign op_I0_8_0 = I0_8_0; // @[Map2T.scala 15:11]
  assign op_I0_8_1 = I0_8_1; // @[Map2T.scala 15:11]
  assign op_I0_9_0 = I0_9_0; // @[Map2T.scala 15:11]
  assign op_I0_9_1 = I0_9_1; // @[Map2T.scala 15:11]
  assign op_I0_10_0 = I0_10_0; // @[Map2T.scala 15:11]
  assign op_I0_10_1 = I0_10_1; // @[Map2T.scala 15:11]
  assign op_I0_11_0 = I0_11_0; // @[Map2T.scala 15:11]
  assign op_I0_11_1 = I0_11_1; // @[Map2T.scala 15:11]
  assign op_I0_12_0 = I0_12_0; // @[Map2T.scala 15:11]
  assign op_I0_12_1 = I0_12_1; // @[Map2T.scala 15:11]
  assign op_I0_13_0 = I0_13_0; // @[Map2T.scala 15:11]
  assign op_I0_13_1 = I0_13_1; // @[Map2T.scala 15:11]
  assign op_I0_14_0 = I0_14_0; // @[Map2T.scala 15:11]
  assign op_I0_14_1 = I0_14_1; // @[Map2T.scala 15:11]
  assign op_I0_15_0 = I0_15_0; // @[Map2T.scala 15:11]
  assign op_I0_15_1 = I0_15_1; // @[Map2T.scala 15:11]
  assign op_I1_0_0 = I1_0_0; // @[Map2T.scala 16:11]
  assign op_I1_0_1 = I1_0_1; // @[Map2T.scala 16:11]
  assign op_I1_1_0 = I1_1_0; // @[Map2T.scala 16:11]
  assign op_I1_1_1 = I1_1_1; // @[Map2T.scala 16:11]
  assign op_I1_2_0 = I1_2_0; // @[Map2T.scala 16:11]
  assign op_I1_2_1 = I1_2_1; // @[Map2T.scala 16:11]
  assign op_I1_3_0 = I1_3_0; // @[Map2T.scala 16:11]
  assign op_I1_3_1 = I1_3_1; // @[Map2T.scala 16:11]
  assign op_I1_4_0 = I1_4_0; // @[Map2T.scala 16:11]
  assign op_I1_4_1 = I1_4_1; // @[Map2T.scala 16:11]
  assign op_I1_5_0 = I1_5_0; // @[Map2T.scala 16:11]
  assign op_I1_5_1 = I1_5_1; // @[Map2T.scala 16:11]
  assign op_I1_6_0 = I1_6_0; // @[Map2T.scala 16:11]
  assign op_I1_6_1 = I1_6_1; // @[Map2T.scala 16:11]
  assign op_I1_7_0 = I1_7_0; // @[Map2T.scala 16:11]
  assign op_I1_7_1 = I1_7_1; // @[Map2T.scala 16:11]
  assign op_I1_8_0 = I1_8_0; // @[Map2T.scala 16:11]
  assign op_I1_8_1 = I1_8_1; // @[Map2T.scala 16:11]
  assign op_I1_9_0 = I1_9_0; // @[Map2T.scala 16:11]
  assign op_I1_9_1 = I1_9_1; // @[Map2T.scala 16:11]
  assign op_I1_10_0 = I1_10_0; // @[Map2T.scala 16:11]
  assign op_I1_10_1 = I1_10_1; // @[Map2T.scala 16:11]
  assign op_I1_11_0 = I1_11_0; // @[Map2T.scala 16:11]
  assign op_I1_11_1 = I1_11_1; // @[Map2T.scala 16:11]
  assign op_I1_12_0 = I1_12_0; // @[Map2T.scala 16:11]
  assign op_I1_12_1 = I1_12_1; // @[Map2T.scala 16:11]
  assign op_I1_13_0 = I1_13_0; // @[Map2T.scala 16:11]
  assign op_I1_13_1 = I1_13_1; // @[Map2T.scala 16:11]
  assign op_I1_14_0 = I1_14_0; // @[Map2T.scala 16:11]
  assign op_I1_14_1 = I1_14_1; // @[Map2T.scala 16:11]
  assign op_I1_15_0 = I1_15_0; // @[Map2T.scala 16:11]
  assign op_I1_15_1 = I1_15_1; // @[Map2T.scala 16:11]
endmodule
module PartitionS_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1
);
  assign valid_down = valid_up; // @[Partition.scala 18:14]
  assign O_0_0_0_0 = I_0_0_0; // @[Partition.scala 15:39]
  assign O_0_0_0_1 = I_0_0_1; // @[Partition.scala 15:39]
  assign O_0_0_1_0 = I_0_1_0; // @[Partition.scala 15:39]
  assign O_0_0_1_1 = I_0_1_1; // @[Partition.scala 15:39]
  assign O_1_0_0_0 = I_1_0_0; // @[Partition.scala 15:39]
  assign O_1_0_0_1 = I_1_0_1; // @[Partition.scala 15:39]
  assign O_1_0_1_0 = I_1_1_0; // @[Partition.scala 15:39]
  assign O_1_0_1_1 = I_1_1_1; // @[Partition.scala 15:39]
  assign O_2_0_0_0 = I_2_0_0; // @[Partition.scala 15:39]
  assign O_2_0_0_1 = I_2_0_1; // @[Partition.scala 15:39]
  assign O_2_0_1_0 = I_2_1_0; // @[Partition.scala 15:39]
  assign O_2_0_1_1 = I_2_1_1; // @[Partition.scala 15:39]
  assign O_3_0_0_0 = I_3_0_0; // @[Partition.scala 15:39]
  assign O_3_0_0_1 = I_3_0_1; // @[Partition.scala 15:39]
  assign O_3_0_1_0 = I_3_1_0; // @[Partition.scala 15:39]
  assign O_3_0_1_1 = I_3_1_1; // @[Partition.scala 15:39]
  assign O_4_0_0_0 = I_4_0_0; // @[Partition.scala 15:39]
  assign O_4_0_0_1 = I_4_0_1; // @[Partition.scala 15:39]
  assign O_4_0_1_0 = I_4_1_0; // @[Partition.scala 15:39]
  assign O_4_0_1_1 = I_4_1_1; // @[Partition.scala 15:39]
  assign O_5_0_0_0 = I_5_0_0; // @[Partition.scala 15:39]
  assign O_5_0_0_1 = I_5_0_1; // @[Partition.scala 15:39]
  assign O_5_0_1_0 = I_5_1_0; // @[Partition.scala 15:39]
  assign O_5_0_1_1 = I_5_1_1; // @[Partition.scala 15:39]
  assign O_6_0_0_0 = I_6_0_0; // @[Partition.scala 15:39]
  assign O_6_0_0_1 = I_6_0_1; // @[Partition.scala 15:39]
  assign O_6_0_1_0 = I_6_1_0; // @[Partition.scala 15:39]
  assign O_6_0_1_1 = I_6_1_1; // @[Partition.scala 15:39]
  assign O_7_0_0_0 = I_7_0_0; // @[Partition.scala 15:39]
  assign O_7_0_0_1 = I_7_0_1; // @[Partition.scala 15:39]
  assign O_7_0_1_0 = I_7_1_0; // @[Partition.scala 15:39]
  assign O_7_0_1_1 = I_7_1_1; // @[Partition.scala 15:39]
  assign O_8_0_0_0 = I_8_0_0; // @[Partition.scala 15:39]
  assign O_8_0_0_1 = I_8_0_1; // @[Partition.scala 15:39]
  assign O_8_0_1_0 = I_8_1_0; // @[Partition.scala 15:39]
  assign O_8_0_1_1 = I_8_1_1; // @[Partition.scala 15:39]
  assign O_9_0_0_0 = I_9_0_0; // @[Partition.scala 15:39]
  assign O_9_0_0_1 = I_9_0_1; // @[Partition.scala 15:39]
  assign O_9_0_1_0 = I_9_1_0; // @[Partition.scala 15:39]
  assign O_9_0_1_1 = I_9_1_1; // @[Partition.scala 15:39]
  assign O_10_0_0_0 = I_10_0_0; // @[Partition.scala 15:39]
  assign O_10_0_0_1 = I_10_0_1; // @[Partition.scala 15:39]
  assign O_10_0_1_0 = I_10_1_0; // @[Partition.scala 15:39]
  assign O_10_0_1_1 = I_10_1_1; // @[Partition.scala 15:39]
  assign O_11_0_0_0 = I_11_0_0; // @[Partition.scala 15:39]
  assign O_11_0_0_1 = I_11_0_1; // @[Partition.scala 15:39]
  assign O_11_0_1_0 = I_11_1_0; // @[Partition.scala 15:39]
  assign O_11_0_1_1 = I_11_1_1; // @[Partition.scala 15:39]
  assign O_12_0_0_0 = I_12_0_0; // @[Partition.scala 15:39]
  assign O_12_0_0_1 = I_12_0_1; // @[Partition.scala 15:39]
  assign O_12_0_1_0 = I_12_1_0; // @[Partition.scala 15:39]
  assign O_12_0_1_1 = I_12_1_1; // @[Partition.scala 15:39]
  assign O_13_0_0_0 = I_13_0_0; // @[Partition.scala 15:39]
  assign O_13_0_0_1 = I_13_0_1; // @[Partition.scala 15:39]
  assign O_13_0_1_0 = I_13_1_0; // @[Partition.scala 15:39]
  assign O_13_0_1_1 = I_13_1_1; // @[Partition.scala 15:39]
  assign O_14_0_0_0 = I_14_0_0; // @[Partition.scala 15:39]
  assign O_14_0_0_1 = I_14_0_1; // @[Partition.scala 15:39]
  assign O_14_0_1_0 = I_14_1_0; // @[Partition.scala 15:39]
  assign O_14_0_1_1 = I_14_1_1; // @[Partition.scala 15:39]
  assign O_15_0_0_0 = I_15_0_0; // @[Partition.scala 15:39]
  assign O_15_0_0_1 = I_15_0_1; // @[Partition.scala 15:39]
  assign O_15_0_1_0 = I_15_1_0; // @[Partition.scala 15:39]
  assign O_15_0_1_1 = I_15_1_1; // @[Partition.scala 15:39]
endmodule
module MapT_13(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  output [7:0] O_0_0_0_0,
  output [7:0] O_0_0_0_1,
  output [7:0] O_0_0_1_0,
  output [7:0] O_0_0_1_1,
  output [7:0] O_1_0_0_0,
  output [7:0] O_1_0_0_1,
  output [7:0] O_1_0_1_0,
  output [7:0] O_1_0_1_1,
  output [7:0] O_2_0_0_0,
  output [7:0] O_2_0_0_1,
  output [7:0] O_2_0_1_0,
  output [7:0] O_2_0_1_1,
  output [7:0] O_3_0_0_0,
  output [7:0] O_3_0_0_1,
  output [7:0] O_3_0_1_0,
  output [7:0] O_3_0_1_1,
  output [7:0] O_4_0_0_0,
  output [7:0] O_4_0_0_1,
  output [7:0] O_4_0_1_0,
  output [7:0] O_4_0_1_1,
  output [7:0] O_5_0_0_0,
  output [7:0] O_5_0_0_1,
  output [7:0] O_5_0_1_0,
  output [7:0] O_5_0_1_1,
  output [7:0] O_6_0_0_0,
  output [7:0] O_6_0_0_1,
  output [7:0] O_6_0_1_0,
  output [7:0] O_6_0_1_1,
  output [7:0] O_7_0_0_0,
  output [7:0] O_7_0_0_1,
  output [7:0] O_7_0_1_0,
  output [7:0] O_7_0_1_1,
  output [7:0] O_8_0_0_0,
  output [7:0] O_8_0_0_1,
  output [7:0] O_8_0_1_0,
  output [7:0] O_8_0_1_1,
  output [7:0] O_9_0_0_0,
  output [7:0] O_9_0_0_1,
  output [7:0] O_9_0_1_0,
  output [7:0] O_9_0_1_1,
  output [7:0] O_10_0_0_0,
  output [7:0] O_10_0_0_1,
  output [7:0] O_10_0_1_0,
  output [7:0] O_10_0_1_1,
  output [7:0] O_11_0_0_0,
  output [7:0] O_11_0_0_1,
  output [7:0] O_11_0_1_0,
  output [7:0] O_11_0_1_1,
  output [7:0] O_12_0_0_0,
  output [7:0] O_12_0_0_1,
  output [7:0] O_12_0_1_0,
  output [7:0] O_12_0_1_1,
  output [7:0] O_13_0_0_0,
  output [7:0] O_13_0_0_1,
  output [7:0] O_13_0_1_0,
  output [7:0] O_13_0_1_1,
  output [7:0] O_14_0_0_0,
  output [7:0] O_14_0_0_1,
  output [7:0] O_14_0_1_0,
  output [7:0] O_14_0_1_1,
  output [7:0] O_15_0_0_0,
  output [7:0] O_15_0_0_1,
  output [7:0] O_15_0_1_0,
  output [7:0] O_15_0_1_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1_1; // @[MapT.scala 8:20]
  PartitionS_6 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .O_0_0_0_0(op_O_0_0_0_0),
    .O_0_0_0_1(op_O_0_0_0_1),
    .O_0_0_1_0(op_O_0_0_1_0),
    .O_0_0_1_1(op_O_0_0_1_1),
    .O_1_0_0_0(op_O_1_0_0_0),
    .O_1_0_0_1(op_O_1_0_0_1),
    .O_1_0_1_0(op_O_1_0_1_0),
    .O_1_0_1_1(op_O_1_0_1_1),
    .O_2_0_0_0(op_O_2_0_0_0),
    .O_2_0_0_1(op_O_2_0_0_1),
    .O_2_0_1_0(op_O_2_0_1_0),
    .O_2_0_1_1(op_O_2_0_1_1),
    .O_3_0_0_0(op_O_3_0_0_0),
    .O_3_0_0_1(op_O_3_0_0_1),
    .O_3_0_1_0(op_O_3_0_1_0),
    .O_3_0_1_1(op_O_3_0_1_1),
    .O_4_0_0_0(op_O_4_0_0_0),
    .O_4_0_0_1(op_O_4_0_0_1),
    .O_4_0_1_0(op_O_4_0_1_0),
    .O_4_0_1_1(op_O_4_0_1_1),
    .O_5_0_0_0(op_O_5_0_0_0),
    .O_5_0_0_1(op_O_5_0_0_1),
    .O_5_0_1_0(op_O_5_0_1_0),
    .O_5_0_1_1(op_O_5_0_1_1),
    .O_6_0_0_0(op_O_6_0_0_0),
    .O_6_0_0_1(op_O_6_0_0_1),
    .O_6_0_1_0(op_O_6_0_1_0),
    .O_6_0_1_1(op_O_6_0_1_1),
    .O_7_0_0_0(op_O_7_0_0_0),
    .O_7_0_0_1(op_O_7_0_0_1),
    .O_7_0_1_0(op_O_7_0_1_0),
    .O_7_0_1_1(op_O_7_0_1_1),
    .O_8_0_0_0(op_O_8_0_0_0),
    .O_8_0_0_1(op_O_8_0_0_1),
    .O_8_0_1_0(op_O_8_0_1_0),
    .O_8_0_1_1(op_O_8_0_1_1),
    .O_9_0_0_0(op_O_9_0_0_0),
    .O_9_0_0_1(op_O_9_0_0_1),
    .O_9_0_1_0(op_O_9_0_1_0),
    .O_9_0_1_1(op_O_9_0_1_1),
    .O_10_0_0_0(op_O_10_0_0_0),
    .O_10_0_0_1(op_O_10_0_0_1),
    .O_10_0_1_0(op_O_10_0_1_0),
    .O_10_0_1_1(op_O_10_0_1_1),
    .O_11_0_0_0(op_O_11_0_0_0),
    .O_11_0_0_1(op_O_11_0_0_1),
    .O_11_0_1_0(op_O_11_0_1_0),
    .O_11_0_1_1(op_O_11_0_1_1),
    .O_12_0_0_0(op_O_12_0_0_0),
    .O_12_0_0_1(op_O_12_0_0_1),
    .O_12_0_1_0(op_O_12_0_1_0),
    .O_12_0_1_1(op_O_12_0_1_1),
    .O_13_0_0_0(op_O_13_0_0_0),
    .O_13_0_0_1(op_O_13_0_0_1),
    .O_13_0_1_0(op_O_13_0_1_0),
    .O_13_0_1_1(op_O_13_0_1_1),
    .O_14_0_0_0(op_O_14_0_0_0),
    .O_14_0_0_1(op_O_14_0_0_1),
    .O_14_0_1_0(op_O_14_0_1_0),
    .O_14_0_1_1(op_O_14_0_1_1),
    .O_15_0_0_0(op_O_15_0_0_0),
    .O_15_0_0_1(op_O_15_0_0_1),
    .O_15_0_1_0(op_O_15_0_1_0),
    .O_15_0_1_1(op_O_15_0_1_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0_0 = op_O_0_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_0_1 = op_O_0_0_0_1; // @[MapT.scala 15:7]
  assign O_0_0_1_0 = op_O_0_0_1_0; // @[MapT.scala 15:7]
  assign O_0_0_1_1 = op_O_0_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_0_0 = op_O_1_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0_1 = op_O_1_0_0_1; // @[MapT.scala 15:7]
  assign O_1_0_1_0 = op_O_1_0_1_0; // @[MapT.scala 15:7]
  assign O_1_0_1_1 = op_O_1_0_1_1; // @[MapT.scala 15:7]
  assign O_2_0_0_0 = op_O_2_0_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0_1 = op_O_2_0_0_1; // @[MapT.scala 15:7]
  assign O_2_0_1_0 = op_O_2_0_1_0; // @[MapT.scala 15:7]
  assign O_2_0_1_1 = op_O_2_0_1_1; // @[MapT.scala 15:7]
  assign O_3_0_0_0 = op_O_3_0_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0_1 = op_O_3_0_0_1; // @[MapT.scala 15:7]
  assign O_3_0_1_0 = op_O_3_0_1_0; // @[MapT.scala 15:7]
  assign O_3_0_1_1 = op_O_3_0_1_1; // @[MapT.scala 15:7]
  assign O_4_0_0_0 = op_O_4_0_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0_1 = op_O_4_0_0_1; // @[MapT.scala 15:7]
  assign O_4_0_1_0 = op_O_4_0_1_0; // @[MapT.scala 15:7]
  assign O_4_0_1_1 = op_O_4_0_1_1; // @[MapT.scala 15:7]
  assign O_5_0_0_0 = op_O_5_0_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0_1 = op_O_5_0_0_1; // @[MapT.scala 15:7]
  assign O_5_0_1_0 = op_O_5_0_1_0; // @[MapT.scala 15:7]
  assign O_5_0_1_1 = op_O_5_0_1_1; // @[MapT.scala 15:7]
  assign O_6_0_0_0 = op_O_6_0_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0_1 = op_O_6_0_0_1; // @[MapT.scala 15:7]
  assign O_6_0_1_0 = op_O_6_0_1_0; // @[MapT.scala 15:7]
  assign O_6_0_1_1 = op_O_6_0_1_1; // @[MapT.scala 15:7]
  assign O_7_0_0_0 = op_O_7_0_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0_1 = op_O_7_0_0_1; // @[MapT.scala 15:7]
  assign O_7_0_1_0 = op_O_7_0_1_0; // @[MapT.scala 15:7]
  assign O_7_0_1_1 = op_O_7_0_1_1; // @[MapT.scala 15:7]
  assign O_8_0_0_0 = op_O_8_0_0_0; // @[MapT.scala 15:7]
  assign O_8_0_0_1 = op_O_8_0_0_1; // @[MapT.scala 15:7]
  assign O_8_0_1_0 = op_O_8_0_1_0; // @[MapT.scala 15:7]
  assign O_8_0_1_1 = op_O_8_0_1_1; // @[MapT.scala 15:7]
  assign O_9_0_0_0 = op_O_9_0_0_0; // @[MapT.scala 15:7]
  assign O_9_0_0_1 = op_O_9_0_0_1; // @[MapT.scala 15:7]
  assign O_9_0_1_0 = op_O_9_0_1_0; // @[MapT.scala 15:7]
  assign O_9_0_1_1 = op_O_9_0_1_1; // @[MapT.scala 15:7]
  assign O_10_0_0_0 = op_O_10_0_0_0; // @[MapT.scala 15:7]
  assign O_10_0_0_1 = op_O_10_0_0_1; // @[MapT.scala 15:7]
  assign O_10_0_1_0 = op_O_10_0_1_0; // @[MapT.scala 15:7]
  assign O_10_0_1_1 = op_O_10_0_1_1; // @[MapT.scala 15:7]
  assign O_11_0_0_0 = op_O_11_0_0_0; // @[MapT.scala 15:7]
  assign O_11_0_0_1 = op_O_11_0_0_1; // @[MapT.scala 15:7]
  assign O_11_0_1_0 = op_O_11_0_1_0; // @[MapT.scala 15:7]
  assign O_11_0_1_1 = op_O_11_0_1_1; // @[MapT.scala 15:7]
  assign O_12_0_0_0 = op_O_12_0_0_0; // @[MapT.scala 15:7]
  assign O_12_0_0_1 = op_O_12_0_0_1; // @[MapT.scala 15:7]
  assign O_12_0_1_0 = op_O_12_0_1_0; // @[MapT.scala 15:7]
  assign O_12_0_1_1 = op_O_12_0_1_1; // @[MapT.scala 15:7]
  assign O_13_0_0_0 = op_O_13_0_0_0; // @[MapT.scala 15:7]
  assign O_13_0_0_1 = op_O_13_0_0_1; // @[MapT.scala 15:7]
  assign O_13_0_1_0 = op_O_13_0_1_0; // @[MapT.scala 15:7]
  assign O_13_0_1_1 = op_O_13_0_1_1; // @[MapT.scala 15:7]
  assign O_14_0_0_0 = op_O_14_0_0_0; // @[MapT.scala 15:7]
  assign O_14_0_0_1 = op_O_14_0_0_1; // @[MapT.scala 15:7]
  assign O_14_0_1_0 = op_O_14_0_1_0; // @[MapT.scala 15:7]
  assign O_14_0_1_1 = op_O_14_0_1_1; // @[MapT.scala 15:7]
  assign O_15_0_0_0 = op_O_15_0_0_0; // @[MapT.scala 15:7]
  assign O_15_0_0_1 = op_O_15_0_0_1; // @[MapT.scala 15:7]
  assign O_15_0_1_0 = op_O_15_0_1_0; // @[MapT.scala 15:7]
  assign O_15_0_1_1 = op_O_15_0_1_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
endmodule
module SSeqTupleToSSeq_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1
);
  assign valid_down = valid_up; // @[Tuple.scala 42:14]
  assign O_0_0 = I_0_0; // @[Tuple.scala 41:5]
  assign O_0_1 = I_0_1; // @[Tuple.scala 41:5]
  assign O_1_0 = I_1_0; // @[Tuple.scala 41:5]
  assign O_1_1 = I_1_1; // @[Tuple.scala 41:5]
endmodule
module Remove1S_6(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1
);
  wire  op_inst_valid_up; // @[Remove1S.scala 9:23]
  wire  op_inst_valid_down; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_I_1_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_0_1; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_0; // @[Remove1S.scala 9:23]
  wire [7:0] op_inst_O_1_1; // @[Remove1S.scala 9:23]
  SSeqTupleToSSeq_6 op_inst ( // @[Remove1S.scala 9:23]
    .valid_up(op_inst_valid_up),
    .valid_down(op_inst_valid_down),
    .I_0_0(op_inst_I_0_0),
    .I_0_1(op_inst_I_0_1),
    .I_1_0(op_inst_I_1_0),
    .I_1_1(op_inst_I_1_1),
    .O_0_0(op_inst_O_0_0),
    .O_0_1(op_inst_O_0_1),
    .O_1_0(op_inst_O_1_0),
    .O_1_1(op_inst_O_1_1)
  );
  assign valid_down = op_inst_valid_down; // @[Remove1S.scala 16:14]
  assign O_0_0 = op_inst_O_0_0; // @[Remove1S.scala 14:5]
  assign O_0_1 = op_inst_O_0_1; // @[Remove1S.scala 14:5]
  assign O_1_0 = op_inst_O_1_0; // @[Remove1S.scala 14:5]
  assign O_1_1 = op_inst_O_1_1; // @[Remove1S.scala 14:5]
  assign op_inst_valid_up = valid_up; // @[Remove1S.scala 15:20]
  assign op_inst_I_0_0 = I_0_0_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_0_1 = I_0_0_1; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_0 = I_0_1_0; // @[Remove1S.scala 13:13]
  assign op_inst_I_1_1 = I_0_1_1; // @[Remove1S.scala 13:13]
endmodule
module MapS_12(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_1_0,
  input  [7:0] I_8_0_1_1,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_1_0,
  input  [7:0] I_9_0_1_1,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_1_0,
  input  [7:0] I_10_0_1_1,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_1_0,
  input  [7:0] I_11_0_1_1,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_1_0,
  input  [7:0] I_12_0_1_1,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_1_0,
  input  [7:0] I_13_0_1_1,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_1_0,
  input  [7:0] I_14_0_1_1,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_1_0,
  input  [7:0] I_15_0_1_1,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1_1; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_1_1; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_1_1; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Remove1S_6 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0_0(fst_op_I_0_0_0),
    .I_0_0_1(fst_op_I_0_0_1),
    .I_0_1_0(fst_op_I_0_1_0),
    .I_0_1_1(fst_op_I_0_1_1),
    .O_0_0(fst_op_O_0_0),
    .O_0_1(fst_op_O_0_1),
    .O_1_0(fst_op_O_1_0),
    .O_1_1(fst_op_O_1_1)
  );
  Remove1S_6 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0_0(other_ops_0_I_0_0_0),
    .I_0_0_1(other_ops_0_I_0_0_1),
    .I_0_1_0(other_ops_0_I_0_1_0),
    .I_0_1_1(other_ops_0_I_0_1_1),
    .O_0_0(other_ops_0_O_0_0),
    .O_0_1(other_ops_0_O_0_1),
    .O_1_0(other_ops_0_O_1_0),
    .O_1_1(other_ops_0_O_1_1)
  );
  Remove1S_6 other_ops_1 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0_0(other_ops_1_I_0_0_0),
    .I_0_0_1(other_ops_1_I_0_0_1),
    .I_0_1_0(other_ops_1_I_0_1_0),
    .I_0_1_1(other_ops_1_I_0_1_1),
    .O_0_0(other_ops_1_O_0_0),
    .O_0_1(other_ops_1_O_0_1),
    .O_1_0(other_ops_1_O_1_0),
    .O_1_1(other_ops_1_O_1_1)
  );
  Remove1S_6 other_ops_2 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0_0(other_ops_2_I_0_0_0),
    .I_0_0_1(other_ops_2_I_0_0_1),
    .I_0_1_0(other_ops_2_I_0_1_0),
    .I_0_1_1(other_ops_2_I_0_1_1),
    .O_0_0(other_ops_2_O_0_0),
    .O_0_1(other_ops_2_O_0_1),
    .O_1_0(other_ops_2_O_1_0),
    .O_1_1(other_ops_2_O_1_1)
  );
  Remove1S_6 other_ops_3 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0_0(other_ops_3_I_0_0_0),
    .I_0_0_1(other_ops_3_I_0_0_1),
    .I_0_1_0(other_ops_3_I_0_1_0),
    .I_0_1_1(other_ops_3_I_0_1_1),
    .O_0_0(other_ops_3_O_0_0),
    .O_0_1(other_ops_3_O_0_1),
    .O_1_0(other_ops_3_O_1_0),
    .O_1_1(other_ops_3_O_1_1)
  );
  Remove1S_6 other_ops_4 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0_0(other_ops_4_I_0_0_0),
    .I_0_0_1(other_ops_4_I_0_0_1),
    .I_0_1_0(other_ops_4_I_0_1_0),
    .I_0_1_1(other_ops_4_I_0_1_1),
    .O_0_0(other_ops_4_O_0_0),
    .O_0_1(other_ops_4_O_0_1),
    .O_1_0(other_ops_4_O_1_0),
    .O_1_1(other_ops_4_O_1_1)
  );
  Remove1S_6 other_ops_5 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0_0(other_ops_5_I_0_0_0),
    .I_0_0_1(other_ops_5_I_0_0_1),
    .I_0_1_0(other_ops_5_I_0_1_0),
    .I_0_1_1(other_ops_5_I_0_1_1),
    .O_0_0(other_ops_5_O_0_0),
    .O_0_1(other_ops_5_O_0_1),
    .O_1_0(other_ops_5_O_1_0),
    .O_1_1(other_ops_5_O_1_1)
  );
  Remove1S_6 other_ops_6 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0_0(other_ops_6_I_0_0_0),
    .I_0_0_1(other_ops_6_I_0_0_1),
    .I_0_1_0(other_ops_6_I_0_1_0),
    .I_0_1_1(other_ops_6_I_0_1_1),
    .O_0_0(other_ops_6_O_0_0),
    .O_0_1(other_ops_6_O_0_1),
    .O_1_0(other_ops_6_O_1_0),
    .O_1_1(other_ops_6_O_1_1)
  );
  Remove1S_6 other_ops_7 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0_0(other_ops_7_I_0_0_0),
    .I_0_0_1(other_ops_7_I_0_0_1),
    .I_0_1_0(other_ops_7_I_0_1_0),
    .I_0_1_1(other_ops_7_I_0_1_1),
    .O_0_0(other_ops_7_O_0_0),
    .O_0_1(other_ops_7_O_0_1),
    .O_1_0(other_ops_7_O_1_0),
    .O_1_1(other_ops_7_O_1_1)
  );
  Remove1S_6 other_ops_8 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0_0(other_ops_8_I_0_0_0),
    .I_0_0_1(other_ops_8_I_0_0_1),
    .I_0_1_0(other_ops_8_I_0_1_0),
    .I_0_1_1(other_ops_8_I_0_1_1),
    .O_0_0(other_ops_8_O_0_0),
    .O_0_1(other_ops_8_O_0_1),
    .O_1_0(other_ops_8_O_1_0),
    .O_1_1(other_ops_8_O_1_1)
  );
  Remove1S_6 other_ops_9 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0_0(other_ops_9_I_0_0_0),
    .I_0_0_1(other_ops_9_I_0_0_1),
    .I_0_1_0(other_ops_9_I_0_1_0),
    .I_0_1_1(other_ops_9_I_0_1_1),
    .O_0_0(other_ops_9_O_0_0),
    .O_0_1(other_ops_9_O_0_1),
    .O_1_0(other_ops_9_O_1_0),
    .O_1_1(other_ops_9_O_1_1)
  );
  Remove1S_6 other_ops_10 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0_0(other_ops_10_I_0_0_0),
    .I_0_0_1(other_ops_10_I_0_0_1),
    .I_0_1_0(other_ops_10_I_0_1_0),
    .I_0_1_1(other_ops_10_I_0_1_1),
    .O_0_0(other_ops_10_O_0_0),
    .O_0_1(other_ops_10_O_0_1),
    .O_1_0(other_ops_10_O_1_0),
    .O_1_1(other_ops_10_O_1_1)
  );
  Remove1S_6 other_ops_11 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0_0(other_ops_11_I_0_0_0),
    .I_0_0_1(other_ops_11_I_0_0_1),
    .I_0_1_0(other_ops_11_I_0_1_0),
    .I_0_1_1(other_ops_11_I_0_1_1),
    .O_0_0(other_ops_11_O_0_0),
    .O_0_1(other_ops_11_O_0_1),
    .O_1_0(other_ops_11_O_1_0),
    .O_1_1(other_ops_11_O_1_1)
  );
  Remove1S_6 other_ops_12 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0_0(other_ops_12_I_0_0_0),
    .I_0_0_1(other_ops_12_I_0_0_1),
    .I_0_1_0(other_ops_12_I_0_1_0),
    .I_0_1_1(other_ops_12_I_0_1_1),
    .O_0_0(other_ops_12_O_0_0),
    .O_0_1(other_ops_12_O_0_1),
    .O_1_0(other_ops_12_O_1_0),
    .O_1_1(other_ops_12_O_1_1)
  );
  Remove1S_6 other_ops_13 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0_0(other_ops_13_I_0_0_0),
    .I_0_0_1(other_ops_13_I_0_0_1),
    .I_0_1_0(other_ops_13_I_0_1_0),
    .I_0_1_1(other_ops_13_I_0_1_1),
    .O_0_0(other_ops_13_O_0_0),
    .O_0_1(other_ops_13_O_0_1),
    .O_1_0(other_ops_13_O_1_0),
    .O_1_1(other_ops_13_O_1_1)
  );
  Remove1S_6 other_ops_14 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0_0(other_ops_14_I_0_0_0),
    .I_0_0_1(other_ops_14_I_0_0_1),
    .I_0_1_0(other_ops_14_I_0_1_0),
    .I_0_1_1(other_ops_14_I_0_1_1),
    .O_0_0(other_ops_14_O_0_0),
    .O_0_1(other_ops_14_O_0_1),
    .O_1_0(other_ops_14_O_1_0),
    .O_1_1(other_ops_14_O_1_1)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_0_0_1 = fst_op_O_0_1; // @[MapS.scala 17:8]
  assign O_0_1_0 = fst_op_O_1_0; // @[MapS.scala 17:8]
  assign O_0_1_1 = fst_op_O_1_1; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_1_0_1 = other_ops_0_O_0_1; // @[MapS.scala 21:12]
  assign O_1_1_0 = other_ops_0_O_1_0; // @[MapS.scala 21:12]
  assign O_1_1_1 = other_ops_0_O_1_1; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_1 = other_ops_1_O_0_1; // @[MapS.scala 21:12]
  assign O_2_1_0 = other_ops_1_O_1_0; // @[MapS.scala 21:12]
  assign O_2_1_1 = other_ops_1_O_1_1; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_1 = other_ops_2_O_0_1; // @[MapS.scala 21:12]
  assign O_3_1_0 = other_ops_2_O_1_0; // @[MapS.scala 21:12]
  assign O_3_1_1 = other_ops_2_O_1_1; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_1 = other_ops_3_O_0_1; // @[MapS.scala 21:12]
  assign O_4_1_0 = other_ops_3_O_1_0; // @[MapS.scala 21:12]
  assign O_4_1_1 = other_ops_3_O_1_1; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_1 = other_ops_4_O_0_1; // @[MapS.scala 21:12]
  assign O_5_1_0 = other_ops_4_O_1_0; // @[MapS.scala 21:12]
  assign O_5_1_1 = other_ops_4_O_1_1; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_1 = other_ops_5_O_0_1; // @[MapS.scala 21:12]
  assign O_6_1_0 = other_ops_5_O_1_0; // @[MapS.scala 21:12]
  assign O_6_1_1 = other_ops_5_O_1_1; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_1 = other_ops_6_O_0_1; // @[MapS.scala 21:12]
  assign O_7_1_0 = other_ops_6_O_1_0; // @[MapS.scala 21:12]
  assign O_7_1_1 = other_ops_6_O_1_1; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_1 = other_ops_7_O_0_1; // @[MapS.scala 21:12]
  assign O_8_1_0 = other_ops_7_O_1_0; // @[MapS.scala 21:12]
  assign O_8_1_1 = other_ops_7_O_1_1; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_1 = other_ops_8_O_0_1; // @[MapS.scala 21:12]
  assign O_9_1_0 = other_ops_8_O_1_0; // @[MapS.scala 21:12]
  assign O_9_1_1 = other_ops_8_O_1_1; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_1 = other_ops_9_O_0_1; // @[MapS.scala 21:12]
  assign O_10_1_0 = other_ops_9_O_1_0; // @[MapS.scala 21:12]
  assign O_10_1_1 = other_ops_9_O_1_1; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_1 = other_ops_10_O_0_1; // @[MapS.scala 21:12]
  assign O_11_1_0 = other_ops_10_O_1_0; // @[MapS.scala 21:12]
  assign O_11_1_1 = other_ops_10_O_1_1; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_1 = other_ops_11_O_0_1; // @[MapS.scala 21:12]
  assign O_12_1_0 = other_ops_11_O_1_0; // @[MapS.scala 21:12]
  assign O_12_1_1 = other_ops_11_O_1_1; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_1 = other_ops_12_O_0_1; // @[MapS.scala 21:12]
  assign O_13_1_0 = other_ops_12_O_1_0; // @[MapS.scala 21:12]
  assign O_13_1_1 = other_ops_12_O_1_1; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_1 = other_ops_13_O_0_1; // @[MapS.scala 21:12]
  assign O_14_1_0 = other_ops_13_O_1_0; // @[MapS.scala 21:12]
  assign O_14_1_1 = other_ops_13_O_1_1; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_1 = other_ops_14_O_0_1; // @[MapS.scala 21:12]
  assign O_15_1_0 = other_ops_14_O_1_0; // @[MapS.scala 21:12]
  assign O_15_1_1 = other_ops_14_O_1_1; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0_0 = I_0_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_0_1 = I_0_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_0 = I_0_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1_1 = I_0_0_1_1; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0_0 = I_1_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_0_1 = I_1_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_0 = I_1_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1_1 = I_1_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0_0 = I_2_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_0_1 = I_2_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_0 = I_2_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1_1 = I_2_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0_0 = I_3_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_0_1 = I_3_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_0 = I_3_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1_1 = I_3_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0_0 = I_4_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_0_1 = I_4_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_0 = I_4_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1_1 = I_4_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0_0 = I_5_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_0_1 = I_5_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_0 = I_5_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1_1 = I_5_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0_0 = I_6_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_0_1 = I_6_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_0 = I_6_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1_1 = I_6_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0_0 = I_7_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_0_1 = I_7_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_0 = I_7_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1_1 = I_7_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0_0 = I_8_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_0_1 = I_8_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_0 = I_8_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1_1 = I_8_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0_0 = I_9_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_0_1 = I_9_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_0 = I_9_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1_1 = I_9_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0_0 = I_10_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_0_1 = I_10_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_0 = I_10_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1_1 = I_10_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0_0 = I_11_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_0_1 = I_11_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_0 = I_11_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1_1 = I_11_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0_0 = I_12_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_0_1 = I_12_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_0 = I_12_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1_1 = I_12_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0_0 = I_13_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_0_1 = I_13_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_0 = I_13_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1_1 = I_13_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0_0 = I_14_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_0_1 = I_14_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_0 = I_14_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1_1 = I_14_0_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0_0 = I_15_0_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_0_1 = I_15_0_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_0 = I_15_0_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1_1 = I_15_0_1_1; // @[MapS.scala 20:41]
endmodule
module MapT_14(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0_0,
  input  [7:0] I_0_0_0_1,
  input  [7:0] I_0_0_1_0,
  input  [7:0] I_0_0_1_1,
  input  [7:0] I_1_0_0_0,
  input  [7:0] I_1_0_0_1,
  input  [7:0] I_1_0_1_0,
  input  [7:0] I_1_0_1_1,
  input  [7:0] I_2_0_0_0,
  input  [7:0] I_2_0_0_1,
  input  [7:0] I_2_0_1_0,
  input  [7:0] I_2_0_1_1,
  input  [7:0] I_3_0_0_0,
  input  [7:0] I_3_0_0_1,
  input  [7:0] I_3_0_1_0,
  input  [7:0] I_3_0_1_1,
  input  [7:0] I_4_0_0_0,
  input  [7:0] I_4_0_0_1,
  input  [7:0] I_4_0_1_0,
  input  [7:0] I_4_0_1_1,
  input  [7:0] I_5_0_0_0,
  input  [7:0] I_5_0_0_1,
  input  [7:0] I_5_0_1_0,
  input  [7:0] I_5_0_1_1,
  input  [7:0] I_6_0_0_0,
  input  [7:0] I_6_0_0_1,
  input  [7:0] I_6_0_1_0,
  input  [7:0] I_6_0_1_1,
  input  [7:0] I_7_0_0_0,
  input  [7:0] I_7_0_0_1,
  input  [7:0] I_7_0_1_0,
  input  [7:0] I_7_0_1_1,
  input  [7:0] I_8_0_0_0,
  input  [7:0] I_8_0_0_1,
  input  [7:0] I_8_0_1_0,
  input  [7:0] I_8_0_1_1,
  input  [7:0] I_9_0_0_0,
  input  [7:0] I_9_0_0_1,
  input  [7:0] I_9_0_1_0,
  input  [7:0] I_9_0_1_1,
  input  [7:0] I_10_0_0_0,
  input  [7:0] I_10_0_0_1,
  input  [7:0] I_10_0_1_0,
  input  [7:0] I_10_0_1_1,
  input  [7:0] I_11_0_0_0,
  input  [7:0] I_11_0_0_1,
  input  [7:0] I_11_0_1_0,
  input  [7:0] I_11_0_1_1,
  input  [7:0] I_12_0_0_0,
  input  [7:0] I_12_0_0_1,
  input  [7:0] I_12_0_1_0,
  input  [7:0] I_12_0_1_1,
  input  [7:0] I_13_0_0_0,
  input  [7:0] I_13_0_0_1,
  input  [7:0] I_13_0_1_0,
  input  [7:0] I_13_0_1_1,
  input  [7:0] I_14_0_0_0,
  input  [7:0] I_14_0_0_1,
  input  [7:0] I_14_0_1_0,
  input  [7:0] I_14_0_1_1,
  input  [7:0] I_15_0_0_0,
  input  [7:0] I_15_0_0_1,
  input  [7:0] I_15_0_1_0,
  input  [7:0] I_15_0_1_1,
  output [7:0] O_0_0_0,
  output [7:0] O_0_0_1,
  output [7:0] O_0_1_0,
  output [7:0] O_0_1_1,
  output [7:0] O_1_0_0,
  output [7:0] O_1_0_1,
  output [7:0] O_1_1_0,
  output [7:0] O_1_1_1,
  output [7:0] O_2_0_0,
  output [7:0] O_2_0_1,
  output [7:0] O_2_1_0,
  output [7:0] O_2_1_1,
  output [7:0] O_3_0_0,
  output [7:0] O_3_0_1,
  output [7:0] O_3_1_0,
  output [7:0] O_3_1_1,
  output [7:0] O_4_0_0,
  output [7:0] O_4_0_1,
  output [7:0] O_4_1_0,
  output [7:0] O_4_1_1,
  output [7:0] O_5_0_0,
  output [7:0] O_5_0_1,
  output [7:0] O_5_1_0,
  output [7:0] O_5_1_1,
  output [7:0] O_6_0_0,
  output [7:0] O_6_0_1,
  output [7:0] O_6_1_0,
  output [7:0] O_6_1_1,
  output [7:0] O_7_0_0,
  output [7:0] O_7_0_1,
  output [7:0] O_7_1_0,
  output [7:0] O_7_1_1,
  output [7:0] O_8_0_0,
  output [7:0] O_8_0_1,
  output [7:0] O_8_1_0,
  output [7:0] O_8_1_1,
  output [7:0] O_9_0_0,
  output [7:0] O_9_0_1,
  output [7:0] O_9_1_0,
  output [7:0] O_9_1_1,
  output [7:0] O_10_0_0,
  output [7:0] O_10_0_1,
  output [7:0] O_10_1_0,
  output [7:0] O_10_1_1,
  output [7:0] O_11_0_0,
  output [7:0] O_11_0_1,
  output [7:0] O_11_1_0,
  output [7:0] O_11_1_1,
  output [7:0] O_12_0_0,
  output [7:0] O_12_0_1,
  output [7:0] O_12_1_0,
  output [7:0] O_12_1_1,
  output [7:0] O_13_0_0,
  output [7:0] O_13_0_1,
  output [7:0] O_13_1_0,
  output [7:0] O_13_1_1,
  output [7:0] O_14_0_0,
  output [7:0] O_14_0_1,
  output [7:0] O_14_1_0,
  output [7:0] O_14_1_1,
  output [7:0] O_15_0_0,
  output [7:0] O_15_0_1,
  output [7:0] O_15_1_0,
  output [7:0] O_15_1_1
);
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_1_1; // @[MapT.scala 8:20]
  MapS_12 op ( // @[MapT.scala 8:20]
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0_0(op_I_0_0_0_0),
    .I_0_0_0_1(op_I_0_0_0_1),
    .I_0_0_1_0(op_I_0_0_1_0),
    .I_0_0_1_1(op_I_0_0_1_1),
    .I_1_0_0_0(op_I_1_0_0_0),
    .I_1_0_0_1(op_I_1_0_0_1),
    .I_1_0_1_0(op_I_1_0_1_0),
    .I_1_0_1_1(op_I_1_0_1_1),
    .I_2_0_0_0(op_I_2_0_0_0),
    .I_2_0_0_1(op_I_2_0_0_1),
    .I_2_0_1_0(op_I_2_0_1_0),
    .I_2_0_1_1(op_I_2_0_1_1),
    .I_3_0_0_0(op_I_3_0_0_0),
    .I_3_0_0_1(op_I_3_0_0_1),
    .I_3_0_1_0(op_I_3_0_1_0),
    .I_3_0_1_1(op_I_3_0_1_1),
    .I_4_0_0_0(op_I_4_0_0_0),
    .I_4_0_0_1(op_I_4_0_0_1),
    .I_4_0_1_0(op_I_4_0_1_0),
    .I_4_0_1_1(op_I_4_0_1_1),
    .I_5_0_0_0(op_I_5_0_0_0),
    .I_5_0_0_1(op_I_5_0_0_1),
    .I_5_0_1_0(op_I_5_0_1_0),
    .I_5_0_1_1(op_I_5_0_1_1),
    .I_6_0_0_0(op_I_6_0_0_0),
    .I_6_0_0_1(op_I_6_0_0_1),
    .I_6_0_1_0(op_I_6_0_1_0),
    .I_6_0_1_1(op_I_6_0_1_1),
    .I_7_0_0_0(op_I_7_0_0_0),
    .I_7_0_0_1(op_I_7_0_0_1),
    .I_7_0_1_0(op_I_7_0_1_0),
    .I_7_0_1_1(op_I_7_0_1_1),
    .I_8_0_0_0(op_I_8_0_0_0),
    .I_8_0_0_1(op_I_8_0_0_1),
    .I_8_0_1_0(op_I_8_0_1_0),
    .I_8_0_1_1(op_I_8_0_1_1),
    .I_9_0_0_0(op_I_9_0_0_0),
    .I_9_0_0_1(op_I_9_0_0_1),
    .I_9_0_1_0(op_I_9_0_1_0),
    .I_9_0_1_1(op_I_9_0_1_1),
    .I_10_0_0_0(op_I_10_0_0_0),
    .I_10_0_0_1(op_I_10_0_0_1),
    .I_10_0_1_0(op_I_10_0_1_0),
    .I_10_0_1_1(op_I_10_0_1_1),
    .I_11_0_0_0(op_I_11_0_0_0),
    .I_11_0_0_1(op_I_11_0_0_1),
    .I_11_0_1_0(op_I_11_0_1_0),
    .I_11_0_1_1(op_I_11_0_1_1),
    .I_12_0_0_0(op_I_12_0_0_0),
    .I_12_0_0_1(op_I_12_0_0_1),
    .I_12_0_1_0(op_I_12_0_1_0),
    .I_12_0_1_1(op_I_12_0_1_1),
    .I_13_0_0_0(op_I_13_0_0_0),
    .I_13_0_0_1(op_I_13_0_0_1),
    .I_13_0_1_0(op_I_13_0_1_0),
    .I_13_0_1_1(op_I_13_0_1_1),
    .I_14_0_0_0(op_I_14_0_0_0),
    .I_14_0_0_1(op_I_14_0_0_1),
    .I_14_0_1_0(op_I_14_0_1_0),
    .I_14_0_1_1(op_I_14_0_1_1),
    .I_15_0_0_0(op_I_15_0_0_0),
    .I_15_0_0_1(op_I_15_0_0_1),
    .I_15_0_1_0(op_I_15_0_1_0),
    .I_15_0_1_1(op_I_15_0_1_1),
    .O_0_0_0(op_O_0_0_0),
    .O_0_0_1(op_O_0_0_1),
    .O_0_1_0(op_O_0_1_0),
    .O_0_1_1(op_O_0_1_1),
    .O_1_0_0(op_O_1_0_0),
    .O_1_0_1(op_O_1_0_1),
    .O_1_1_0(op_O_1_1_0),
    .O_1_1_1(op_O_1_1_1),
    .O_2_0_0(op_O_2_0_0),
    .O_2_0_1(op_O_2_0_1),
    .O_2_1_0(op_O_2_1_0),
    .O_2_1_1(op_O_2_1_1),
    .O_3_0_0(op_O_3_0_0),
    .O_3_0_1(op_O_3_0_1),
    .O_3_1_0(op_O_3_1_0),
    .O_3_1_1(op_O_3_1_1),
    .O_4_0_0(op_O_4_0_0),
    .O_4_0_1(op_O_4_0_1),
    .O_4_1_0(op_O_4_1_0),
    .O_4_1_1(op_O_4_1_1),
    .O_5_0_0(op_O_5_0_0),
    .O_5_0_1(op_O_5_0_1),
    .O_5_1_0(op_O_5_1_0),
    .O_5_1_1(op_O_5_1_1),
    .O_6_0_0(op_O_6_0_0),
    .O_6_0_1(op_O_6_0_1),
    .O_6_1_0(op_O_6_1_0),
    .O_6_1_1(op_O_6_1_1),
    .O_7_0_0(op_O_7_0_0),
    .O_7_0_1(op_O_7_0_1),
    .O_7_1_0(op_O_7_1_0),
    .O_7_1_1(op_O_7_1_1),
    .O_8_0_0(op_O_8_0_0),
    .O_8_0_1(op_O_8_0_1),
    .O_8_1_0(op_O_8_1_0),
    .O_8_1_1(op_O_8_1_1),
    .O_9_0_0(op_O_9_0_0),
    .O_9_0_1(op_O_9_0_1),
    .O_9_1_0(op_O_9_1_0),
    .O_9_1_1(op_O_9_1_1),
    .O_10_0_0(op_O_10_0_0),
    .O_10_0_1(op_O_10_0_1),
    .O_10_1_0(op_O_10_1_0),
    .O_10_1_1(op_O_10_1_1),
    .O_11_0_0(op_O_11_0_0),
    .O_11_0_1(op_O_11_0_1),
    .O_11_1_0(op_O_11_1_0),
    .O_11_1_1(op_O_11_1_1),
    .O_12_0_0(op_O_12_0_0),
    .O_12_0_1(op_O_12_0_1),
    .O_12_1_0(op_O_12_1_0),
    .O_12_1_1(op_O_12_1_1),
    .O_13_0_0(op_O_13_0_0),
    .O_13_0_1(op_O_13_0_1),
    .O_13_1_0(op_O_13_1_0),
    .O_13_1_1(op_O_13_1_1),
    .O_14_0_0(op_O_14_0_0),
    .O_14_0_1(op_O_14_0_1),
    .O_14_1_0(op_O_14_1_0),
    .O_14_1_1(op_O_14_1_1),
    .O_15_0_0(op_O_15_0_0),
    .O_15_0_1(op_O_15_0_1),
    .O_15_1_0(op_O_15_1_0),
    .O_15_1_1(op_O_15_1_1)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_0_0_1 = op_O_0_0_1; // @[MapT.scala 15:7]
  assign O_0_1_0 = op_O_0_1_0; // @[MapT.scala 15:7]
  assign O_0_1_1 = op_O_0_1_1; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_1_0_1 = op_O_1_0_1; // @[MapT.scala 15:7]
  assign O_1_1_0 = op_O_1_1_0; // @[MapT.scala 15:7]
  assign O_1_1_1 = op_O_1_1_1; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_2_0_1 = op_O_2_0_1; // @[MapT.scala 15:7]
  assign O_2_1_0 = op_O_2_1_0; // @[MapT.scala 15:7]
  assign O_2_1_1 = op_O_2_1_1; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_3_0_1 = op_O_3_0_1; // @[MapT.scala 15:7]
  assign O_3_1_0 = op_O_3_1_0; // @[MapT.scala 15:7]
  assign O_3_1_1 = op_O_3_1_1; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_4_0_1 = op_O_4_0_1; // @[MapT.scala 15:7]
  assign O_4_1_0 = op_O_4_1_0; // @[MapT.scala 15:7]
  assign O_4_1_1 = op_O_4_1_1; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_5_0_1 = op_O_5_0_1; // @[MapT.scala 15:7]
  assign O_5_1_0 = op_O_5_1_0; // @[MapT.scala 15:7]
  assign O_5_1_1 = op_O_5_1_1; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_6_0_1 = op_O_6_0_1; // @[MapT.scala 15:7]
  assign O_6_1_0 = op_O_6_1_0; // @[MapT.scala 15:7]
  assign O_6_1_1 = op_O_6_1_1; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_7_0_1 = op_O_7_0_1; // @[MapT.scala 15:7]
  assign O_7_1_0 = op_O_7_1_0; // @[MapT.scala 15:7]
  assign O_7_1_1 = op_O_7_1_1; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_8_0_1 = op_O_8_0_1; // @[MapT.scala 15:7]
  assign O_8_1_0 = op_O_8_1_0; // @[MapT.scala 15:7]
  assign O_8_1_1 = op_O_8_1_1; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_9_0_1 = op_O_9_0_1; // @[MapT.scala 15:7]
  assign O_9_1_0 = op_O_9_1_0; // @[MapT.scala 15:7]
  assign O_9_1_1 = op_O_9_1_1; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_10_0_1 = op_O_10_0_1; // @[MapT.scala 15:7]
  assign O_10_1_0 = op_O_10_1_0; // @[MapT.scala 15:7]
  assign O_10_1_1 = op_O_10_1_1; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_11_0_1 = op_O_11_0_1; // @[MapT.scala 15:7]
  assign O_11_1_0 = op_O_11_1_0; // @[MapT.scala 15:7]
  assign O_11_1_1 = op_O_11_1_1; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_12_0_1 = op_O_12_0_1; // @[MapT.scala 15:7]
  assign O_12_1_0 = op_O_12_1_0; // @[MapT.scala 15:7]
  assign O_12_1_1 = op_O_12_1_1; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_13_0_1 = op_O_13_0_1; // @[MapT.scala 15:7]
  assign O_13_1_0 = op_O_13_1_0; // @[MapT.scala 15:7]
  assign O_13_1_1 = op_O_13_1_1; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_14_0_1 = op_O_14_0_1; // @[MapT.scala 15:7]
  assign O_14_1_0 = op_O_14_1_0; // @[MapT.scala 15:7]
  assign O_14_1_1 = op_O_14_1_1; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign O_15_0_1 = op_O_15_0_1; // @[MapT.scala 15:7]
  assign O_15_1_0 = op_O_15_1_0; // @[MapT.scala 15:7]
  assign O_15_1_1 = op_O_15_1_1; // @[MapT.scala 15:7]
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0_0 = I_0_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_0_1 = I_0_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_0_1_0 = I_0_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1_1 = I_0_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0_0 = I_1_0_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_0_1 = I_1_0_0_1; // @[MapT.scala 14:10]
  assign op_I_1_0_1_0 = I_1_0_1_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1_1 = I_1_0_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0_0 = I_2_0_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_0_1 = I_2_0_0_1; // @[MapT.scala 14:10]
  assign op_I_2_0_1_0 = I_2_0_1_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1_1 = I_2_0_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0_0 = I_3_0_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_0_1 = I_3_0_0_1; // @[MapT.scala 14:10]
  assign op_I_3_0_1_0 = I_3_0_1_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1_1 = I_3_0_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0_0 = I_4_0_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_0_1 = I_4_0_0_1; // @[MapT.scala 14:10]
  assign op_I_4_0_1_0 = I_4_0_1_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1_1 = I_4_0_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0_0 = I_5_0_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_0_1 = I_5_0_0_1; // @[MapT.scala 14:10]
  assign op_I_5_0_1_0 = I_5_0_1_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1_1 = I_5_0_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0_0 = I_6_0_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_0_1 = I_6_0_0_1; // @[MapT.scala 14:10]
  assign op_I_6_0_1_0 = I_6_0_1_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1_1 = I_6_0_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0_0 = I_7_0_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_0_1 = I_7_0_0_1; // @[MapT.scala 14:10]
  assign op_I_7_0_1_0 = I_7_0_1_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1_1 = I_7_0_1_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0_0 = I_8_0_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_0_1 = I_8_0_0_1; // @[MapT.scala 14:10]
  assign op_I_8_0_1_0 = I_8_0_1_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1_1 = I_8_0_1_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0_0 = I_9_0_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_0_1 = I_9_0_0_1; // @[MapT.scala 14:10]
  assign op_I_9_0_1_0 = I_9_0_1_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1_1 = I_9_0_1_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0_0 = I_10_0_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_0_1 = I_10_0_0_1; // @[MapT.scala 14:10]
  assign op_I_10_0_1_0 = I_10_0_1_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1_1 = I_10_0_1_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0_0 = I_11_0_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_0_1 = I_11_0_0_1; // @[MapT.scala 14:10]
  assign op_I_11_0_1_0 = I_11_0_1_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1_1 = I_11_0_1_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0_0 = I_12_0_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_0_1 = I_12_0_0_1; // @[MapT.scala 14:10]
  assign op_I_12_0_1_0 = I_12_0_1_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1_1 = I_12_0_1_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0_0 = I_13_0_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_0_1 = I_13_0_0_1; // @[MapT.scala 14:10]
  assign op_I_13_0_1_0 = I_13_0_1_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1_1 = I_13_0_1_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0_0 = I_14_0_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_0_1 = I_14_0_0_1; // @[MapT.scala 14:10]
  assign op_I_14_0_1_0 = I_14_0_1_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1_1 = I_14_0_1_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0_0 = I_15_0_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_0_1 = I_15_0_0_1; // @[MapT.scala 14:10]
  assign op_I_15_0_1_0 = I_15_0_1_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1_1 = I_15_0_1_1; // @[MapT.scala 14:10]
endmodule
module Map2S_15(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0,
  input  [7:0] I0_1,
  input  [7:0] I1_0,
  input  [7:0] I1_1,
  output [7:0] O_0_t0b,
  output [7:0] O_0_t1b,
  output [7:0] O_1_t0b,
  output [7:0] O_1_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_t1b; // @[Map2S.scala 10:86]
  AtomTuple fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0(fst_op_I0),
    .I1(fst_op_I1),
    .O_t0b(fst_op_O_t0b),
    .O_t1b(fst_op_O_t1b)
  );
  AtomTuple other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0(other_ops_0_I0),
    .I1(other_ops_0_I1),
    .O_t0b(other_ops_0_O_t0b),
    .O_t1b(other_ops_0_O_t1b)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_t0b = fst_op_O_t0b; // @[Map2S.scala 19:8]
  assign O_0_t1b = fst_op_O_t1b; // @[Map2S.scala 19:8]
  assign O_1_t0b = other_ops_0_O_t0b; // @[Map2S.scala 24:12]
  assign O_1_t1b = other_ops_0_O_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0 = I0_0; // @[Map2S.scala 17:13]
  assign fst_op_I1 = I1_0; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0 = I0_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1 = I1_1; // @[Map2S.scala 23:43]
endmodule
module Map2S_16(
  input        valid_up,
  output       valid_down,
  input  [7:0] I0_0_0,
  input  [7:0] I0_0_1,
  input  [7:0] I0_1_0,
  input  [7:0] I0_1_1,
  output [7:0] O_0_0_t0b,
  output [7:0] O_0_0_t1b,
  output [7:0] O_0_1_t0b,
  output [7:0] O_0_1_t1b,
  output [7:0] O_1_0_t0b,
  output [7:0] O_1_0_t1b,
  output [7:0] O_1_1_t0b,
  output [7:0] O_1_1_t1b
);
  wire  fst_op_valid_up; // @[Map2S.scala 9:22]
  wire  fst_op_valid_down; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I0_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_0; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_I1_1; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_0_t1b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t0b; // @[Map2S.scala 9:22]
  wire [7:0] fst_op_O_1_t1b; // @[Map2S.scala 9:22]
  wire  other_ops_0_valid_up; // @[Map2S.scala 10:86]
  wire  other_ops_0_valid_down; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I0_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_0; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_I1_1; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_0_t1b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t0b; // @[Map2S.scala 10:86]
  wire [7:0] other_ops_0_O_1_t1b; // @[Map2S.scala 10:86]
  Map2S_15 fst_op ( // @[Map2S.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I0_0(fst_op_I0_0),
    .I0_1(fst_op_I0_1),
    .I1_0(fst_op_I1_0),
    .I1_1(fst_op_I1_1),
    .O_0_t0b(fst_op_O_0_t0b),
    .O_0_t1b(fst_op_O_0_t1b),
    .O_1_t0b(fst_op_O_1_t0b),
    .O_1_t1b(fst_op_O_1_t1b)
  );
  Map2S_15 other_ops_0 ( // @[Map2S.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I0_0(other_ops_0_I0_0),
    .I0_1(other_ops_0_I0_1),
    .I1_0(other_ops_0_I1_0),
    .I1_1(other_ops_0_I1_1),
    .O_0_t0b(other_ops_0_O_0_t0b),
    .O_0_t1b(other_ops_0_O_0_t1b),
    .O_1_t0b(other_ops_0_O_1_t0b),
    .O_1_t1b(other_ops_0_O_1_t1b)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[Map2S.scala 26:14]
  assign O_0_0_t0b = fst_op_O_0_t0b; // @[Map2S.scala 19:8]
  assign O_0_0_t1b = fst_op_O_0_t1b; // @[Map2S.scala 19:8]
  assign O_0_1_t0b = fst_op_O_1_t0b; // @[Map2S.scala 19:8]
  assign O_0_1_t1b = fst_op_O_1_t1b; // @[Map2S.scala 19:8]
  assign O_1_0_t0b = other_ops_0_O_0_t0b; // @[Map2S.scala 24:12]
  assign O_1_0_t1b = other_ops_0_O_0_t1b; // @[Map2S.scala 24:12]
  assign O_1_1_t0b = other_ops_0_O_1_t0b; // @[Map2S.scala 24:12]
  assign O_1_1_t1b = other_ops_0_O_1_t1b; // @[Map2S.scala 24:12]
  assign fst_op_valid_up = valid_up; // @[Map2S.scala 16:19]
  assign fst_op_I0_0 = I0_0_0; // @[Map2S.scala 17:13]
  assign fst_op_I0_1 = I0_0_1; // @[Map2S.scala 17:13]
  assign fst_op_I1_0 = 8'h0; // @[Map2S.scala 18:13]
  assign fst_op_I1_1 = 8'h2; // @[Map2S.scala 18:13]
  assign other_ops_0_valid_up = valid_up; // @[Map2S.scala 21:39]
  assign other_ops_0_I0_0 = I0_1_0; // @[Map2S.scala 22:43]
  assign other_ops_0_I0_1 = I0_1_1; // @[Map2S.scala 22:43]
  assign other_ops_0_I1_0 = 8'h1; // @[Map2S.scala 23:43]
  assign other_ops_0_I1_1 = 8'h0; // @[Map2S.scala 23:43]
endmodule
module MapS_13(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_t0b,
  input  [7:0] I_0_t1b,
  input  [7:0] I_1_t0b,
  input  [7:0] I_1_t1b,
  output [7:0] O_0,
  output [7:0] O_1
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O; // @[MapS.scala 10:86]
  LShift fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_t0b(fst_op_I_t0b),
    .I_t1b(fst_op_I_t1b),
    .O(fst_op_O)
  );
  LShift other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_t0b(other_ops_0_I_t0b),
    .I_t1b(other_ops_0_I_t1b),
    .O(other_ops_0_O)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0 = fst_op_O; // @[MapS.scala 17:8]
  assign O_1 = other_ops_0_O; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_t0b = I_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_t1b = I_0_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_t0b = I_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_t1b = I_1_t1b; // @[MapS.scala 20:41]
endmodule
module MapS_14(
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_t0b,
  input  [7:0] I_0_0_t1b,
  input  [7:0] I_0_1_t0b,
  input  [7:0] I_0_1_t1b,
  input  [7:0] I_1_0_t0b,
  input  [7:0] I_1_0_t1b,
  input  [7:0] I_1_1_t0b,
  input  [7:0] I_1_1_t1b,
  output [7:0] O_0_0,
  output [7:0] O_0_1,
  output [7:0] O_1_0,
  output [7:0] O_1_1
);
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t0b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_t1b; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_1; // @[MapS.scala 9:22]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t0b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_t1b; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_1; // @[MapS.scala 10:86]
  MapS_13 fst_op ( // @[MapS.scala 9:22]
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_t0b(fst_op_I_0_t0b),
    .I_0_t1b(fst_op_I_0_t1b),
    .I_1_t0b(fst_op_I_1_t0b),
    .I_1_t1b(fst_op_I_1_t1b),
    .O_0(fst_op_O_0),
    .O_1(fst_op_O_1)
  );
  MapS_13 other_ops_0 ( // @[MapS.scala 10:86]
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_t0b(other_ops_0_I_0_t0b),
    .I_0_t1b(other_ops_0_I_0_t1b),
    .I_1_t0b(other_ops_0_I_1_t0b),
    .I_1_t1b(other_ops_0_I_1_t1b),
    .O_0(other_ops_0_O_0),
    .O_1(other_ops_0_O_1)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_0_1 = fst_op_O_1; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign O_1_1 = other_ops_0_O_1; // @[MapS.scala 21:12]
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_t0b = I_0_0_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_0_t1b = I_0_0_t1b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t0b = I_0_1_t0b; // @[MapS.scala 16:12]
  assign fst_op_I_1_t1b = I_0_1_t1b; // @[MapS.scala 16:12]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_t0b = I_1_0_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_t1b = I_1_0_t1b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t0b = I_1_1_t0b; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_t1b = I_1_1_t1b; // @[MapS.scala 20:41]
endmodule
module ReduceS_2(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  output [7:0] O_0
);
  wire [7:0] AddNoValid_I_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_I_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] AddNoValid_O; // @[ReduceS.scala 20:43]
  reg [7:0] _T; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  AddNoValid AddNoValid ( // @[ReduceS.scala 20:43]
    .I_t0b(AddNoValid_I_t0b),
    .I_t1b(AddNoValid_I_t1b),
    .O(AddNoValid_O)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0 = _T; // @[ReduceS.scala 27:14]
  assign AddNoValid_I_t0b = I_0; // @[ReduceS.scala 43:18]
  assign AddNoValid_I_t1b = I_1; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= AddNoValid_O;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module MapS_15(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  output [7:0] O_0_0,
  output [7:0] O_1_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0; // @[MapS.scala 10:86]
  ReduceS_2 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0(fst_op_I_0),
    .I_1(fst_op_I_1),
    .O_0(fst_op_O_0)
  );
  ReduceS_2 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0(other_ops_0_I_0),
    .I_1(other_ops_0_I_1),
    .O_0(other_ops_0_O_0)
  );
  assign valid_down = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:14]
  assign O_0_0 = fst_op_O_0; // @[MapS.scala 17:8]
  assign O_1_0 = other_ops_0_O_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0 = I_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_1 = I_0_1; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0 = I_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1 = I_1_1; // @[MapS.scala 20:41]
endmodule
module ReduceS_3(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_1_0,
  output [7:0] O_0_0
);
  wire [7:0] MapSNoValid_I_0_t0b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_I_0_t1b; // @[ReduceS.scala 20:43]
  wire [7:0] MapSNoValid_O_0; // @[ReduceS.scala 20:43]
  reg [7:0] _T_0; // @[ReduceS.scala 27:24]
  reg [31:0] _RAND_0;
  reg  _T_1; // @[ReduceS.scala 47:24]
  reg [31:0] _RAND_1;
  MapSNoValid MapSNoValid ( // @[ReduceS.scala 20:43]
    .I_0_t0b(MapSNoValid_I_0_t0b),
    .I_0_t1b(MapSNoValid_I_0_t1b),
    .O_0(MapSNoValid_O_0)
  );
  assign valid_down = _T_1; // @[ReduceS.scala 47:14]
  assign O_0_0 = _T_0; // @[ReduceS.scala 27:14]
  assign MapSNoValid_I_0_t0b = I_0_0; // @[ReduceS.scala 43:18]
  assign MapSNoValid_I_0_t1b = I_1_0; // @[ReduceS.scala 43:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_0 = _RAND_0[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_0 <= MapSNoValid_O_0;
    if (reset) begin
      _T_1 <= 1'h0;
    end else begin
      _T_1 <= valid_up;
    end
  end
endmodule
module InitialDelayCounter_3(
  input   clock,
  input   reset,
  output  valid_down
);
  reg [2:0] value; // @[InitialDelayCounter.scala 8:34]
  reg [31:0] _RAND_0;
  wire  _T_1; // @[InitialDelayCounter.scala 17:17]
  wire [2:0] _T_4; // @[InitialDelayCounter.scala 17:53]
  assign _T_1 = value < 3'h5; // @[InitialDelayCounter.scala 17:17]
  assign _T_4 = value + 3'h1; // @[InitialDelayCounter.scala 17:53]
  assign valid_down = value == 3'h5; // @[InitialDelayCounter.scala 16:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_1) begin
      value <= _T_4;
    end
  end
endmodule
module Module_1(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0,
  input  [7:0] I_0_1,
  input  [7:0] I_1_0,
  input  [7:0] I_1_1,
  output [7:0] O_0_0
);
  wire  InitialDelayCounter_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_valid_down; // @[Const.scala 11:33]
  wire  n208_valid_up; // @[Top.scala 46:22]
  wire  n208_valid_down; // @[Top.scala 46:22]
  wire [7:0] n208_I0_0_0; // @[Top.scala 46:22]
  wire [7:0] n208_I0_0_1; // @[Top.scala 46:22]
  wire [7:0] n208_I0_1_0; // @[Top.scala 46:22]
  wire [7:0] n208_I0_1_1; // @[Top.scala 46:22]
  wire [7:0] n208_O_0_0_t0b; // @[Top.scala 46:22]
  wire [7:0] n208_O_0_0_t1b; // @[Top.scala 46:22]
  wire [7:0] n208_O_0_1_t0b; // @[Top.scala 46:22]
  wire [7:0] n208_O_0_1_t1b; // @[Top.scala 46:22]
  wire [7:0] n208_O_1_0_t0b; // @[Top.scala 46:22]
  wire [7:0] n208_O_1_0_t1b; // @[Top.scala 46:22]
  wire [7:0] n208_O_1_1_t0b; // @[Top.scala 46:22]
  wire [7:0] n208_O_1_1_t1b; // @[Top.scala 46:22]
  wire  n219_valid_up; // @[Top.scala 50:22]
  wire  n219_valid_down; // @[Top.scala 50:22]
  wire [7:0] n219_I_0_0_t0b; // @[Top.scala 50:22]
  wire [7:0] n219_I_0_0_t1b; // @[Top.scala 50:22]
  wire [7:0] n219_I_0_1_t0b; // @[Top.scala 50:22]
  wire [7:0] n219_I_0_1_t1b; // @[Top.scala 50:22]
  wire [7:0] n219_I_1_0_t0b; // @[Top.scala 50:22]
  wire [7:0] n219_I_1_0_t1b; // @[Top.scala 50:22]
  wire [7:0] n219_I_1_1_t0b; // @[Top.scala 50:22]
  wire [7:0] n219_I_1_1_t1b; // @[Top.scala 50:22]
  wire [7:0] n219_O_0_0; // @[Top.scala 50:22]
  wire [7:0] n219_O_0_1; // @[Top.scala 50:22]
  wire [7:0] n219_O_1_0; // @[Top.scala 50:22]
  wire [7:0] n219_O_1_1; // @[Top.scala 50:22]
  wire  n224_clock; // @[Top.scala 53:22]
  wire  n224_reset; // @[Top.scala 53:22]
  wire  n224_valid_up; // @[Top.scala 53:22]
  wire  n224_valid_down; // @[Top.scala 53:22]
  wire [7:0] n224_I_0_0; // @[Top.scala 53:22]
  wire [7:0] n224_I_0_1; // @[Top.scala 53:22]
  wire [7:0] n224_I_1_0; // @[Top.scala 53:22]
  wire [7:0] n224_I_1_1; // @[Top.scala 53:22]
  wire [7:0] n224_O_0_0; // @[Top.scala 53:22]
  wire [7:0] n224_O_1_0; // @[Top.scala 53:22]
  wire  n229_clock; // @[Top.scala 56:22]
  wire  n229_reset; // @[Top.scala 56:22]
  wire  n229_valid_up; // @[Top.scala 56:22]
  wire  n229_valid_down; // @[Top.scala 56:22]
  wire [7:0] n229_I_0_0; // @[Top.scala 56:22]
  wire [7:0] n229_I_1_0; // @[Top.scala 56:22]
  wire [7:0] n229_O_0_0; // @[Top.scala 56:22]
  wire  InitialDelayCounter_1_clock; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_reset; // @[Const.scala 11:33]
  wire  InitialDelayCounter_1_valid_down; // @[Const.scala 11:33]
  wire  n232_valid_up; // @[Top.scala 60:22]
  wire  n232_valid_down; // @[Top.scala 60:22]
  wire [7:0] n232_I0_0_0; // @[Top.scala 60:22]
  wire [7:0] n232_I1_0_0; // @[Top.scala 60:22]
  wire [7:0] n232_O_0_0_t0b; // @[Top.scala 60:22]
  wire [7:0] n232_O_0_0_t1b; // @[Top.scala 60:22]
  wire  n243_valid_up; // @[Top.scala 64:22]
  wire  n243_valid_down; // @[Top.scala 64:22]
  wire [7:0] n243_I_0_0_t0b; // @[Top.scala 64:22]
  wire [7:0] n243_I_0_0_t1b; // @[Top.scala 64:22]
  wire [7:0] n243_O_0_0; // @[Top.scala 64:22]
  InitialDelayCounter_1 InitialDelayCounter ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_clock),
    .reset(InitialDelayCounter_reset),
    .valid_down(InitialDelayCounter_valid_down)
  );
  Map2S_16 n208 ( // @[Top.scala 46:22]
    .valid_up(n208_valid_up),
    .valid_down(n208_valid_down),
    .I0_0_0(n208_I0_0_0),
    .I0_0_1(n208_I0_0_1),
    .I0_1_0(n208_I0_1_0),
    .I0_1_1(n208_I0_1_1),
    .O_0_0_t0b(n208_O_0_0_t0b),
    .O_0_0_t1b(n208_O_0_0_t1b),
    .O_0_1_t0b(n208_O_0_1_t0b),
    .O_0_1_t1b(n208_O_0_1_t1b),
    .O_1_0_t0b(n208_O_1_0_t0b),
    .O_1_0_t1b(n208_O_1_0_t1b),
    .O_1_1_t0b(n208_O_1_1_t0b),
    .O_1_1_t1b(n208_O_1_1_t1b)
  );
  MapS_14 n219 ( // @[Top.scala 50:22]
    .valid_up(n219_valid_up),
    .valid_down(n219_valid_down),
    .I_0_0_t0b(n219_I_0_0_t0b),
    .I_0_0_t1b(n219_I_0_0_t1b),
    .I_0_1_t0b(n219_I_0_1_t0b),
    .I_0_1_t1b(n219_I_0_1_t1b),
    .I_1_0_t0b(n219_I_1_0_t0b),
    .I_1_0_t1b(n219_I_1_0_t1b),
    .I_1_1_t0b(n219_I_1_1_t0b),
    .I_1_1_t1b(n219_I_1_1_t1b),
    .O_0_0(n219_O_0_0),
    .O_0_1(n219_O_0_1),
    .O_1_0(n219_O_1_0),
    .O_1_1(n219_O_1_1)
  );
  MapS_15 n224 ( // @[Top.scala 53:22]
    .clock(n224_clock),
    .reset(n224_reset),
    .valid_up(n224_valid_up),
    .valid_down(n224_valid_down),
    .I_0_0(n224_I_0_0),
    .I_0_1(n224_I_0_1),
    .I_1_0(n224_I_1_0),
    .I_1_1(n224_I_1_1),
    .O_0_0(n224_O_0_0),
    .O_1_0(n224_O_1_0)
  );
  ReduceS_3 n229 ( // @[Top.scala 56:22]
    .clock(n229_clock),
    .reset(n229_reset),
    .valid_up(n229_valid_up),
    .valid_down(n229_valid_down),
    .I_0_0(n229_I_0_0),
    .I_1_0(n229_I_1_0),
    .O_0_0(n229_O_0_0)
  );
  InitialDelayCounter_3 InitialDelayCounter_1 ( // @[Const.scala 11:33]
    .clock(InitialDelayCounter_1_clock),
    .reset(InitialDelayCounter_1_reset),
    .valid_down(InitialDelayCounter_1_valid_down)
  );
  Map2S_11 n232 ( // @[Top.scala 60:22]
    .valid_up(n232_valid_up),
    .valid_down(n232_valid_down),
    .I0_0_0(n232_I0_0_0),
    .I1_0_0(n232_I1_0_0),
    .O_0_0_t0b(n232_O_0_0_t0b),
    .O_0_0_t1b(n232_O_0_0_t1b)
  );
  MapS_8 n243 ( // @[Top.scala 64:22]
    .valid_up(n243_valid_up),
    .valid_down(n243_valid_down),
    .I_0_0_t0b(n243_I_0_0_t0b),
    .I_0_0_t1b(n243_I_0_0_t1b),
    .O_0_0(n243_O_0_0)
  );
  assign valid_down = n243_valid_down; // @[Top.scala 68:16]
  assign O_0_0 = n243_O_0_0; // @[Top.scala 67:7]
  assign InitialDelayCounter_clock = clock;
  assign InitialDelayCounter_reset = reset;
  assign n208_valid_up = valid_up & InitialDelayCounter_valid_down; // @[Top.scala 49:19]
  assign n208_I0_0_0 = I_0_0; // @[Top.scala 47:13]
  assign n208_I0_0_1 = I_0_1; // @[Top.scala 47:13]
  assign n208_I0_1_0 = I_1_0; // @[Top.scala 47:13]
  assign n208_I0_1_1 = I_1_1; // @[Top.scala 47:13]
  assign n219_valid_up = n208_valid_down; // @[Top.scala 52:19]
  assign n219_I_0_0_t0b = n208_O_0_0_t0b; // @[Top.scala 51:12]
  assign n219_I_0_0_t1b = n208_O_0_0_t1b; // @[Top.scala 51:12]
  assign n219_I_0_1_t0b = n208_O_0_1_t0b; // @[Top.scala 51:12]
  assign n219_I_0_1_t1b = n208_O_0_1_t1b; // @[Top.scala 51:12]
  assign n219_I_1_0_t0b = n208_O_1_0_t0b; // @[Top.scala 51:12]
  assign n219_I_1_0_t1b = n208_O_1_0_t1b; // @[Top.scala 51:12]
  assign n219_I_1_1_t0b = n208_O_1_1_t0b; // @[Top.scala 51:12]
  assign n219_I_1_1_t1b = n208_O_1_1_t1b; // @[Top.scala 51:12]
  assign n224_clock = clock;
  assign n224_reset = reset;
  assign n224_valid_up = n219_valid_down; // @[Top.scala 55:19]
  assign n224_I_0_0 = n219_O_0_0; // @[Top.scala 54:12]
  assign n224_I_0_1 = n219_O_0_1; // @[Top.scala 54:12]
  assign n224_I_1_0 = n219_O_1_0; // @[Top.scala 54:12]
  assign n224_I_1_1 = n219_O_1_1; // @[Top.scala 54:12]
  assign n229_clock = clock;
  assign n229_reset = reset;
  assign n229_valid_up = n224_valid_down; // @[Top.scala 58:19]
  assign n229_I_0_0 = n224_O_0_0; // @[Top.scala 57:12]
  assign n229_I_1_0 = n224_O_1_0; // @[Top.scala 57:12]
  assign InitialDelayCounter_1_clock = clock;
  assign InitialDelayCounter_1_reset = reset;
  assign n232_valid_up = n229_valid_down & InitialDelayCounter_1_valid_down; // @[Top.scala 63:19]
  assign n232_I0_0_0 = n229_O_0_0; // @[Top.scala 61:13]
  assign n232_I1_0_0 = 8'h3; // @[Top.scala 62:13]
  assign n243_valid_up = n232_valid_down; // @[Top.scala 66:19]
  assign n243_I_0_0_t0b = n232_O_0_0_t0b; // @[Top.scala 65:12]
  assign n243_I_0_0_t1b = n232_O_0_0_t1b; // @[Top.scala 65:12]
endmodule
module MapS_18(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  fst_op_clock; // @[MapS.scala 9:22]
  wire  fst_op_reset; // @[MapS.scala 9:22]
  wire  fst_op_valid_up; // @[MapS.scala 9:22]
  wire  fst_op_valid_down; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_0_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_0; // @[MapS.scala 9:22]
  wire [7:0] fst_op_I_1_1; // @[MapS.scala 9:22]
  wire [7:0] fst_op_O_0_0; // @[MapS.scala 9:22]
  wire  other_ops_0_clock; // @[MapS.scala 10:86]
  wire  other_ops_0_reset; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_0_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_0_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_1_clock; // @[MapS.scala 10:86]
  wire  other_ops_1_reset; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_1_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_1_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_2_clock; // @[MapS.scala 10:86]
  wire  other_ops_2_reset; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_2_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_2_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_3_clock; // @[MapS.scala 10:86]
  wire  other_ops_3_reset; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_3_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_3_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_4_clock; // @[MapS.scala 10:86]
  wire  other_ops_4_reset; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_4_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_4_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_5_clock; // @[MapS.scala 10:86]
  wire  other_ops_5_reset; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_5_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_5_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_6_clock; // @[MapS.scala 10:86]
  wire  other_ops_6_reset; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_6_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_6_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_7_clock; // @[MapS.scala 10:86]
  wire  other_ops_7_reset; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_7_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_7_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_8_clock; // @[MapS.scala 10:86]
  wire  other_ops_8_reset; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_8_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_8_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_9_clock; // @[MapS.scala 10:86]
  wire  other_ops_9_reset; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_9_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_9_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_10_clock; // @[MapS.scala 10:86]
  wire  other_ops_10_reset; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_10_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_10_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_11_clock; // @[MapS.scala 10:86]
  wire  other_ops_11_reset; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_11_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_11_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_12_clock; // @[MapS.scala 10:86]
  wire  other_ops_12_reset; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_12_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_12_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_13_clock; // @[MapS.scala 10:86]
  wire  other_ops_13_reset; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_13_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_13_O_0_0; // @[MapS.scala 10:86]
  wire  other_ops_14_clock; // @[MapS.scala 10:86]
  wire  other_ops_14_reset; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_up; // @[MapS.scala 10:86]
  wire  other_ops_14_valid_down; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_0_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_0; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_I_1_1; // @[MapS.scala 10:86]
  wire [7:0] other_ops_14_O_0_0; // @[MapS.scala 10:86]
  wire  _T; // @[MapS.scala 23:83]
  wire  _T_1; // @[MapS.scala 23:83]
  wire  _T_2; // @[MapS.scala 23:83]
  wire  _T_3; // @[MapS.scala 23:83]
  wire  _T_4; // @[MapS.scala 23:83]
  wire  _T_5; // @[MapS.scala 23:83]
  wire  _T_6; // @[MapS.scala 23:83]
  wire  _T_7; // @[MapS.scala 23:83]
  wire  _T_8; // @[MapS.scala 23:83]
  wire  _T_9; // @[MapS.scala 23:83]
  wire  _T_10; // @[MapS.scala 23:83]
  wire  _T_11; // @[MapS.scala 23:83]
  wire  _T_12; // @[MapS.scala 23:83]
  wire  _T_13; // @[MapS.scala 23:83]
  Module_1 fst_op ( // @[MapS.scala 9:22]
    .clock(fst_op_clock),
    .reset(fst_op_reset),
    .valid_up(fst_op_valid_up),
    .valid_down(fst_op_valid_down),
    .I_0_0(fst_op_I_0_0),
    .I_0_1(fst_op_I_0_1),
    .I_1_0(fst_op_I_1_0),
    .I_1_1(fst_op_I_1_1),
    .O_0_0(fst_op_O_0_0)
  );
  Module_1 other_ops_0 ( // @[MapS.scala 10:86]
    .clock(other_ops_0_clock),
    .reset(other_ops_0_reset),
    .valid_up(other_ops_0_valid_up),
    .valid_down(other_ops_0_valid_down),
    .I_0_0(other_ops_0_I_0_0),
    .I_0_1(other_ops_0_I_0_1),
    .I_1_0(other_ops_0_I_1_0),
    .I_1_1(other_ops_0_I_1_1),
    .O_0_0(other_ops_0_O_0_0)
  );
  Module_1 other_ops_1 ( // @[MapS.scala 10:86]
    .clock(other_ops_1_clock),
    .reset(other_ops_1_reset),
    .valid_up(other_ops_1_valid_up),
    .valid_down(other_ops_1_valid_down),
    .I_0_0(other_ops_1_I_0_0),
    .I_0_1(other_ops_1_I_0_1),
    .I_1_0(other_ops_1_I_1_0),
    .I_1_1(other_ops_1_I_1_1),
    .O_0_0(other_ops_1_O_0_0)
  );
  Module_1 other_ops_2 ( // @[MapS.scala 10:86]
    .clock(other_ops_2_clock),
    .reset(other_ops_2_reset),
    .valid_up(other_ops_2_valid_up),
    .valid_down(other_ops_2_valid_down),
    .I_0_0(other_ops_2_I_0_0),
    .I_0_1(other_ops_2_I_0_1),
    .I_1_0(other_ops_2_I_1_0),
    .I_1_1(other_ops_2_I_1_1),
    .O_0_0(other_ops_2_O_0_0)
  );
  Module_1 other_ops_3 ( // @[MapS.scala 10:86]
    .clock(other_ops_3_clock),
    .reset(other_ops_3_reset),
    .valid_up(other_ops_3_valid_up),
    .valid_down(other_ops_3_valid_down),
    .I_0_0(other_ops_3_I_0_0),
    .I_0_1(other_ops_3_I_0_1),
    .I_1_0(other_ops_3_I_1_0),
    .I_1_1(other_ops_3_I_1_1),
    .O_0_0(other_ops_3_O_0_0)
  );
  Module_1 other_ops_4 ( // @[MapS.scala 10:86]
    .clock(other_ops_4_clock),
    .reset(other_ops_4_reset),
    .valid_up(other_ops_4_valid_up),
    .valid_down(other_ops_4_valid_down),
    .I_0_0(other_ops_4_I_0_0),
    .I_0_1(other_ops_4_I_0_1),
    .I_1_0(other_ops_4_I_1_0),
    .I_1_1(other_ops_4_I_1_1),
    .O_0_0(other_ops_4_O_0_0)
  );
  Module_1 other_ops_5 ( // @[MapS.scala 10:86]
    .clock(other_ops_5_clock),
    .reset(other_ops_5_reset),
    .valid_up(other_ops_5_valid_up),
    .valid_down(other_ops_5_valid_down),
    .I_0_0(other_ops_5_I_0_0),
    .I_0_1(other_ops_5_I_0_1),
    .I_1_0(other_ops_5_I_1_0),
    .I_1_1(other_ops_5_I_1_1),
    .O_0_0(other_ops_5_O_0_0)
  );
  Module_1 other_ops_6 ( // @[MapS.scala 10:86]
    .clock(other_ops_6_clock),
    .reset(other_ops_6_reset),
    .valid_up(other_ops_6_valid_up),
    .valid_down(other_ops_6_valid_down),
    .I_0_0(other_ops_6_I_0_0),
    .I_0_1(other_ops_6_I_0_1),
    .I_1_0(other_ops_6_I_1_0),
    .I_1_1(other_ops_6_I_1_1),
    .O_0_0(other_ops_6_O_0_0)
  );
  Module_1 other_ops_7 ( // @[MapS.scala 10:86]
    .clock(other_ops_7_clock),
    .reset(other_ops_7_reset),
    .valid_up(other_ops_7_valid_up),
    .valid_down(other_ops_7_valid_down),
    .I_0_0(other_ops_7_I_0_0),
    .I_0_1(other_ops_7_I_0_1),
    .I_1_0(other_ops_7_I_1_0),
    .I_1_1(other_ops_7_I_1_1),
    .O_0_0(other_ops_7_O_0_0)
  );
  Module_1 other_ops_8 ( // @[MapS.scala 10:86]
    .clock(other_ops_8_clock),
    .reset(other_ops_8_reset),
    .valid_up(other_ops_8_valid_up),
    .valid_down(other_ops_8_valid_down),
    .I_0_0(other_ops_8_I_0_0),
    .I_0_1(other_ops_8_I_0_1),
    .I_1_0(other_ops_8_I_1_0),
    .I_1_1(other_ops_8_I_1_1),
    .O_0_0(other_ops_8_O_0_0)
  );
  Module_1 other_ops_9 ( // @[MapS.scala 10:86]
    .clock(other_ops_9_clock),
    .reset(other_ops_9_reset),
    .valid_up(other_ops_9_valid_up),
    .valid_down(other_ops_9_valid_down),
    .I_0_0(other_ops_9_I_0_0),
    .I_0_1(other_ops_9_I_0_1),
    .I_1_0(other_ops_9_I_1_0),
    .I_1_1(other_ops_9_I_1_1),
    .O_0_0(other_ops_9_O_0_0)
  );
  Module_1 other_ops_10 ( // @[MapS.scala 10:86]
    .clock(other_ops_10_clock),
    .reset(other_ops_10_reset),
    .valid_up(other_ops_10_valid_up),
    .valid_down(other_ops_10_valid_down),
    .I_0_0(other_ops_10_I_0_0),
    .I_0_1(other_ops_10_I_0_1),
    .I_1_0(other_ops_10_I_1_0),
    .I_1_1(other_ops_10_I_1_1),
    .O_0_0(other_ops_10_O_0_0)
  );
  Module_1 other_ops_11 ( // @[MapS.scala 10:86]
    .clock(other_ops_11_clock),
    .reset(other_ops_11_reset),
    .valid_up(other_ops_11_valid_up),
    .valid_down(other_ops_11_valid_down),
    .I_0_0(other_ops_11_I_0_0),
    .I_0_1(other_ops_11_I_0_1),
    .I_1_0(other_ops_11_I_1_0),
    .I_1_1(other_ops_11_I_1_1),
    .O_0_0(other_ops_11_O_0_0)
  );
  Module_1 other_ops_12 ( // @[MapS.scala 10:86]
    .clock(other_ops_12_clock),
    .reset(other_ops_12_reset),
    .valid_up(other_ops_12_valid_up),
    .valid_down(other_ops_12_valid_down),
    .I_0_0(other_ops_12_I_0_0),
    .I_0_1(other_ops_12_I_0_1),
    .I_1_0(other_ops_12_I_1_0),
    .I_1_1(other_ops_12_I_1_1),
    .O_0_0(other_ops_12_O_0_0)
  );
  Module_1 other_ops_13 ( // @[MapS.scala 10:86]
    .clock(other_ops_13_clock),
    .reset(other_ops_13_reset),
    .valid_up(other_ops_13_valid_up),
    .valid_down(other_ops_13_valid_down),
    .I_0_0(other_ops_13_I_0_0),
    .I_0_1(other_ops_13_I_0_1),
    .I_1_0(other_ops_13_I_1_0),
    .I_1_1(other_ops_13_I_1_1),
    .O_0_0(other_ops_13_O_0_0)
  );
  Module_1 other_ops_14 ( // @[MapS.scala 10:86]
    .clock(other_ops_14_clock),
    .reset(other_ops_14_reset),
    .valid_up(other_ops_14_valid_up),
    .valid_down(other_ops_14_valid_down),
    .I_0_0(other_ops_14_I_0_0),
    .I_0_1(other_ops_14_I_0_1),
    .I_1_0(other_ops_14_I_1_0),
    .I_1_1(other_ops_14_I_1_1),
    .O_0_0(other_ops_14_O_0_0)
  );
  assign _T = fst_op_valid_down & other_ops_0_valid_down; // @[MapS.scala 23:83]
  assign _T_1 = _T & other_ops_1_valid_down; // @[MapS.scala 23:83]
  assign _T_2 = _T_1 & other_ops_2_valid_down; // @[MapS.scala 23:83]
  assign _T_3 = _T_2 & other_ops_3_valid_down; // @[MapS.scala 23:83]
  assign _T_4 = _T_3 & other_ops_4_valid_down; // @[MapS.scala 23:83]
  assign _T_5 = _T_4 & other_ops_5_valid_down; // @[MapS.scala 23:83]
  assign _T_6 = _T_5 & other_ops_6_valid_down; // @[MapS.scala 23:83]
  assign _T_7 = _T_6 & other_ops_7_valid_down; // @[MapS.scala 23:83]
  assign _T_8 = _T_7 & other_ops_8_valid_down; // @[MapS.scala 23:83]
  assign _T_9 = _T_8 & other_ops_9_valid_down; // @[MapS.scala 23:83]
  assign _T_10 = _T_9 & other_ops_10_valid_down; // @[MapS.scala 23:83]
  assign _T_11 = _T_10 & other_ops_11_valid_down; // @[MapS.scala 23:83]
  assign _T_12 = _T_11 & other_ops_12_valid_down; // @[MapS.scala 23:83]
  assign _T_13 = _T_12 & other_ops_13_valid_down; // @[MapS.scala 23:83]
  assign valid_down = _T_13 & other_ops_14_valid_down; // @[MapS.scala 23:14]
  assign O_0_0_0 = fst_op_O_0_0; // @[MapS.scala 17:8]
  assign O_1_0_0 = other_ops_0_O_0_0; // @[MapS.scala 21:12]
  assign O_2_0_0 = other_ops_1_O_0_0; // @[MapS.scala 21:12]
  assign O_3_0_0 = other_ops_2_O_0_0; // @[MapS.scala 21:12]
  assign O_4_0_0 = other_ops_3_O_0_0; // @[MapS.scala 21:12]
  assign O_5_0_0 = other_ops_4_O_0_0; // @[MapS.scala 21:12]
  assign O_6_0_0 = other_ops_5_O_0_0; // @[MapS.scala 21:12]
  assign O_7_0_0 = other_ops_6_O_0_0; // @[MapS.scala 21:12]
  assign O_8_0_0 = other_ops_7_O_0_0; // @[MapS.scala 21:12]
  assign O_9_0_0 = other_ops_8_O_0_0; // @[MapS.scala 21:12]
  assign O_10_0_0 = other_ops_9_O_0_0; // @[MapS.scala 21:12]
  assign O_11_0_0 = other_ops_10_O_0_0; // @[MapS.scala 21:12]
  assign O_12_0_0 = other_ops_11_O_0_0; // @[MapS.scala 21:12]
  assign O_13_0_0 = other_ops_12_O_0_0; // @[MapS.scala 21:12]
  assign O_14_0_0 = other_ops_13_O_0_0; // @[MapS.scala 21:12]
  assign O_15_0_0 = other_ops_14_O_0_0; // @[MapS.scala 21:12]
  assign fst_op_clock = clock;
  assign fst_op_reset = reset;
  assign fst_op_valid_up = valid_up; // @[MapS.scala 15:19]
  assign fst_op_I_0_0 = I_0_0_0; // @[MapS.scala 16:12]
  assign fst_op_I_0_1 = I_0_0_1; // @[MapS.scala 16:12]
  assign fst_op_I_1_0 = I_0_1_0; // @[MapS.scala 16:12]
  assign fst_op_I_1_1 = I_0_1_1; // @[MapS.scala 16:12]
  assign other_ops_0_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_0_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_0_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_0_I_0_0 = I_1_0_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_0_1 = I_1_0_1; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_0 = I_1_1_0; // @[MapS.scala 20:41]
  assign other_ops_0_I_1_1 = I_1_1_1; // @[MapS.scala 20:41]
  assign other_ops_1_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_1_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_1_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_1_I_0_0 = I_2_0_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_0_1 = I_2_0_1; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_0 = I_2_1_0; // @[MapS.scala 20:41]
  assign other_ops_1_I_1_1 = I_2_1_1; // @[MapS.scala 20:41]
  assign other_ops_2_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_2_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_2_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_2_I_0_0 = I_3_0_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_0_1 = I_3_0_1; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_0 = I_3_1_0; // @[MapS.scala 20:41]
  assign other_ops_2_I_1_1 = I_3_1_1; // @[MapS.scala 20:41]
  assign other_ops_3_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_3_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_3_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_3_I_0_0 = I_4_0_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_0_1 = I_4_0_1; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_0 = I_4_1_0; // @[MapS.scala 20:41]
  assign other_ops_3_I_1_1 = I_4_1_1; // @[MapS.scala 20:41]
  assign other_ops_4_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_4_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_4_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_4_I_0_0 = I_5_0_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_0_1 = I_5_0_1; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_0 = I_5_1_0; // @[MapS.scala 20:41]
  assign other_ops_4_I_1_1 = I_5_1_1; // @[MapS.scala 20:41]
  assign other_ops_5_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_5_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_5_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_5_I_0_0 = I_6_0_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_0_1 = I_6_0_1; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_0 = I_6_1_0; // @[MapS.scala 20:41]
  assign other_ops_5_I_1_1 = I_6_1_1; // @[MapS.scala 20:41]
  assign other_ops_6_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_6_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_6_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_6_I_0_0 = I_7_0_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_0_1 = I_7_0_1; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_0 = I_7_1_0; // @[MapS.scala 20:41]
  assign other_ops_6_I_1_1 = I_7_1_1; // @[MapS.scala 20:41]
  assign other_ops_7_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_7_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_7_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_7_I_0_0 = I_8_0_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_0_1 = I_8_0_1; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_0 = I_8_1_0; // @[MapS.scala 20:41]
  assign other_ops_7_I_1_1 = I_8_1_1; // @[MapS.scala 20:41]
  assign other_ops_8_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_8_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_8_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_8_I_0_0 = I_9_0_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_0_1 = I_9_0_1; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_0 = I_9_1_0; // @[MapS.scala 20:41]
  assign other_ops_8_I_1_1 = I_9_1_1; // @[MapS.scala 20:41]
  assign other_ops_9_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_9_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_9_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_9_I_0_0 = I_10_0_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_0_1 = I_10_0_1; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_0 = I_10_1_0; // @[MapS.scala 20:41]
  assign other_ops_9_I_1_1 = I_10_1_1; // @[MapS.scala 20:41]
  assign other_ops_10_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_10_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_10_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_10_I_0_0 = I_11_0_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_0_1 = I_11_0_1; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_0 = I_11_1_0; // @[MapS.scala 20:41]
  assign other_ops_10_I_1_1 = I_11_1_1; // @[MapS.scala 20:41]
  assign other_ops_11_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_11_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_11_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_11_I_0_0 = I_12_0_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_0_1 = I_12_0_1; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_0 = I_12_1_0; // @[MapS.scala 20:41]
  assign other_ops_11_I_1_1 = I_12_1_1; // @[MapS.scala 20:41]
  assign other_ops_12_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_12_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_12_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_12_I_0_0 = I_13_0_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_0_1 = I_13_0_1; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_0 = I_13_1_0; // @[MapS.scala 20:41]
  assign other_ops_12_I_1_1 = I_13_1_1; // @[MapS.scala 20:41]
  assign other_ops_13_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_13_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_13_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_13_I_0_0 = I_14_0_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_0_1 = I_14_0_1; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_0 = I_14_1_0; // @[MapS.scala 20:41]
  assign other_ops_13_I_1_1 = I_14_1_1; // @[MapS.scala 20:41]
  assign other_ops_14_clock = clock; // @[MapS.scala 10:86]
  assign other_ops_14_reset = reset; // @[MapS.scala 10:86]
  assign other_ops_14_valid_up = valid_up; // @[MapS.scala 19:39]
  assign other_ops_14_I_0_0 = I_15_0_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_0_1 = I_15_0_1; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_0 = I_15_1_0; // @[MapS.scala 20:41]
  assign other_ops_14_I_1_1 = I_15_1_1; // @[MapS.scala 20:41]
endmodule
module MapT_15(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0_0_0,
  input  [7:0] I_0_0_1,
  input  [7:0] I_0_1_0,
  input  [7:0] I_0_1_1,
  input  [7:0] I_1_0_0,
  input  [7:0] I_1_0_1,
  input  [7:0] I_1_1_0,
  input  [7:0] I_1_1_1,
  input  [7:0] I_2_0_0,
  input  [7:0] I_2_0_1,
  input  [7:0] I_2_1_0,
  input  [7:0] I_2_1_1,
  input  [7:0] I_3_0_0,
  input  [7:0] I_3_0_1,
  input  [7:0] I_3_1_0,
  input  [7:0] I_3_1_1,
  input  [7:0] I_4_0_0,
  input  [7:0] I_4_0_1,
  input  [7:0] I_4_1_0,
  input  [7:0] I_4_1_1,
  input  [7:0] I_5_0_0,
  input  [7:0] I_5_0_1,
  input  [7:0] I_5_1_0,
  input  [7:0] I_5_1_1,
  input  [7:0] I_6_0_0,
  input  [7:0] I_6_0_1,
  input  [7:0] I_6_1_0,
  input  [7:0] I_6_1_1,
  input  [7:0] I_7_0_0,
  input  [7:0] I_7_0_1,
  input  [7:0] I_7_1_0,
  input  [7:0] I_7_1_1,
  input  [7:0] I_8_0_0,
  input  [7:0] I_8_0_1,
  input  [7:0] I_8_1_0,
  input  [7:0] I_8_1_1,
  input  [7:0] I_9_0_0,
  input  [7:0] I_9_0_1,
  input  [7:0] I_9_1_0,
  input  [7:0] I_9_1_1,
  input  [7:0] I_10_0_0,
  input  [7:0] I_10_0_1,
  input  [7:0] I_10_1_0,
  input  [7:0] I_10_1_1,
  input  [7:0] I_11_0_0,
  input  [7:0] I_11_0_1,
  input  [7:0] I_11_1_0,
  input  [7:0] I_11_1_1,
  input  [7:0] I_12_0_0,
  input  [7:0] I_12_0_1,
  input  [7:0] I_12_1_0,
  input  [7:0] I_12_1_1,
  input  [7:0] I_13_0_0,
  input  [7:0] I_13_0_1,
  input  [7:0] I_13_1_0,
  input  [7:0] I_13_1_1,
  input  [7:0] I_14_0_0,
  input  [7:0] I_14_0_1,
  input  [7:0] I_14_1_0,
  input  [7:0] I_14_1_1,
  input  [7:0] I_15_0_0,
  input  [7:0] I_15_0_1,
  input  [7:0] I_15_1_0,
  input  [7:0] I_15_1_1,
  output [7:0] O_0_0_0,
  output [7:0] O_1_0_0,
  output [7:0] O_2_0_0,
  output [7:0] O_3_0_0,
  output [7:0] O_4_0_0,
  output [7:0] O_5_0_0,
  output [7:0] O_6_0_0,
  output [7:0] O_7_0_0,
  output [7:0] O_8_0_0,
  output [7:0] O_9_0_0,
  output [7:0] O_10_0_0,
  output [7:0] O_11_0_0,
  output [7:0] O_12_0_0,
  output [7:0] O_13_0_0,
  output [7:0] O_14_0_0,
  output [7:0] O_15_0_0
);
  wire  op_clock; // @[MapT.scala 8:20]
  wire  op_reset; // @[MapT.scala 8:20]
  wire  op_valid_up; // @[MapT.scala 8:20]
  wire  op_valid_down; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_0_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_1_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_2_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_3_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_4_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_5_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_6_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_7_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_8_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_9_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_10_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_11_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_12_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_13_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_14_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_0_1; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_0; // @[MapT.scala 8:20]
  wire [7:0] op_I_15_1_1; // @[MapT.scala 8:20]
  wire [7:0] op_O_0_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_1_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_2_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_3_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_4_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_5_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_6_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_7_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_8_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_9_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_10_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_11_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_12_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_13_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_14_0_0; // @[MapT.scala 8:20]
  wire [7:0] op_O_15_0_0; // @[MapT.scala 8:20]
  MapS_18 op ( // @[MapT.scala 8:20]
    .clock(op_clock),
    .reset(op_reset),
    .valid_up(op_valid_up),
    .valid_down(op_valid_down),
    .I_0_0_0(op_I_0_0_0),
    .I_0_0_1(op_I_0_0_1),
    .I_0_1_0(op_I_0_1_0),
    .I_0_1_1(op_I_0_1_1),
    .I_1_0_0(op_I_1_0_0),
    .I_1_0_1(op_I_1_0_1),
    .I_1_1_0(op_I_1_1_0),
    .I_1_1_1(op_I_1_1_1),
    .I_2_0_0(op_I_2_0_0),
    .I_2_0_1(op_I_2_0_1),
    .I_2_1_0(op_I_2_1_0),
    .I_2_1_1(op_I_2_1_1),
    .I_3_0_0(op_I_3_0_0),
    .I_3_0_1(op_I_3_0_1),
    .I_3_1_0(op_I_3_1_0),
    .I_3_1_1(op_I_3_1_1),
    .I_4_0_0(op_I_4_0_0),
    .I_4_0_1(op_I_4_0_1),
    .I_4_1_0(op_I_4_1_0),
    .I_4_1_1(op_I_4_1_1),
    .I_5_0_0(op_I_5_0_0),
    .I_5_0_1(op_I_5_0_1),
    .I_5_1_0(op_I_5_1_0),
    .I_5_1_1(op_I_5_1_1),
    .I_6_0_0(op_I_6_0_0),
    .I_6_0_1(op_I_6_0_1),
    .I_6_1_0(op_I_6_1_0),
    .I_6_1_1(op_I_6_1_1),
    .I_7_0_0(op_I_7_0_0),
    .I_7_0_1(op_I_7_0_1),
    .I_7_1_0(op_I_7_1_0),
    .I_7_1_1(op_I_7_1_1),
    .I_8_0_0(op_I_8_0_0),
    .I_8_0_1(op_I_8_0_1),
    .I_8_1_0(op_I_8_1_0),
    .I_8_1_1(op_I_8_1_1),
    .I_9_0_0(op_I_9_0_0),
    .I_9_0_1(op_I_9_0_1),
    .I_9_1_0(op_I_9_1_0),
    .I_9_1_1(op_I_9_1_1),
    .I_10_0_0(op_I_10_0_0),
    .I_10_0_1(op_I_10_0_1),
    .I_10_1_0(op_I_10_1_0),
    .I_10_1_1(op_I_10_1_1),
    .I_11_0_0(op_I_11_0_0),
    .I_11_0_1(op_I_11_0_1),
    .I_11_1_0(op_I_11_1_0),
    .I_11_1_1(op_I_11_1_1),
    .I_12_0_0(op_I_12_0_0),
    .I_12_0_1(op_I_12_0_1),
    .I_12_1_0(op_I_12_1_0),
    .I_12_1_1(op_I_12_1_1),
    .I_13_0_0(op_I_13_0_0),
    .I_13_0_1(op_I_13_0_1),
    .I_13_1_0(op_I_13_1_0),
    .I_13_1_1(op_I_13_1_1),
    .I_14_0_0(op_I_14_0_0),
    .I_14_0_1(op_I_14_0_1),
    .I_14_1_0(op_I_14_1_0),
    .I_14_1_1(op_I_14_1_1),
    .I_15_0_0(op_I_15_0_0),
    .I_15_0_1(op_I_15_0_1),
    .I_15_1_0(op_I_15_1_0),
    .I_15_1_1(op_I_15_1_1),
    .O_0_0_0(op_O_0_0_0),
    .O_1_0_0(op_O_1_0_0),
    .O_2_0_0(op_O_2_0_0),
    .O_3_0_0(op_O_3_0_0),
    .O_4_0_0(op_O_4_0_0),
    .O_5_0_0(op_O_5_0_0),
    .O_6_0_0(op_O_6_0_0),
    .O_7_0_0(op_O_7_0_0),
    .O_8_0_0(op_O_8_0_0),
    .O_9_0_0(op_O_9_0_0),
    .O_10_0_0(op_O_10_0_0),
    .O_11_0_0(op_O_11_0_0),
    .O_12_0_0(op_O_12_0_0),
    .O_13_0_0(op_O_13_0_0),
    .O_14_0_0(op_O_14_0_0),
    .O_15_0_0(op_O_15_0_0)
  );
  assign valid_down = op_valid_down; // @[MapT.scala 16:16]
  assign O_0_0_0 = op_O_0_0_0; // @[MapT.scala 15:7]
  assign O_1_0_0 = op_O_1_0_0; // @[MapT.scala 15:7]
  assign O_2_0_0 = op_O_2_0_0; // @[MapT.scala 15:7]
  assign O_3_0_0 = op_O_3_0_0; // @[MapT.scala 15:7]
  assign O_4_0_0 = op_O_4_0_0; // @[MapT.scala 15:7]
  assign O_5_0_0 = op_O_5_0_0; // @[MapT.scala 15:7]
  assign O_6_0_0 = op_O_6_0_0; // @[MapT.scala 15:7]
  assign O_7_0_0 = op_O_7_0_0; // @[MapT.scala 15:7]
  assign O_8_0_0 = op_O_8_0_0; // @[MapT.scala 15:7]
  assign O_9_0_0 = op_O_9_0_0; // @[MapT.scala 15:7]
  assign O_10_0_0 = op_O_10_0_0; // @[MapT.scala 15:7]
  assign O_11_0_0 = op_O_11_0_0; // @[MapT.scala 15:7]
  assign O_12_0_0 = op_O_12_0_0; // @[MapT.scala 15:7]
  assign O_13_0_0 = op_O_13_0_0; // @[MapT.scala 15:7]
  assign O_14_0_0 = op_O_14_0_0; // @[MapT.scala 15:7]
  assign O_15_0_0 = op_O_15_0_0; // @[MapT.scala 15:7]
  assign op_clock = clock;
  assign op_reset = reset;
  assign op_valid_up = valid_up; // @[MapT.scala 13:17]
  assign op_I_0_0_0 = I_0_0_0; // @[MapT.scala 14:10]
  assign op_I_0_0_1 = I_0_0_1; // @[MapT.scala 14:10]
  assign op_I_0_1_0 = I_0_1_0; // @[MapT.scala 14:10]
  assign op_I_0_1_1 = I_0_1_1; // @[MapT.scala 14:10]
  assign op_I_1_0_0 = I_1_0_0; // @[MapT.scala 14:10]
  assign op_I_1_0_1 = I_1_0_1; // @[MapT.scala 14:10]
  assign op_I_1_1_0 = I_1_1_0; // @[MapT.scala 14:10]
  assign op_I_1_1_1 = I_1_1_1; // @[MapT.scala 14:10]
  assign op_I_2_0_0 = I_2_0_0; // @[MapT.scala 14:10]
  assign op_I_2_0_1 = I_2_0_1; // @[MapT.scala 14:10]
  assign op_I_2_1_0 = I_2_1_0; // @[MapT.scala 14:10]
  assign op_I_2_1_1 = I_2_1_1; // @[MapT.scala 14:10]
  assign op_I_3_0_0 = I_3_0_0; // @[MapT.scala 14:10]
  assign op_I_3_0_1 = I_3_0_1; // @[MapT.scala 14:10]
  assign op_I_3_1_0 = I_3_1_0; // @[MapT.scala 14:10]
  assign op_I_3_1_1 = I_3_1_1; // @[MapT.scala 14:10]
  assign op_I_4_0_0 = I_4_0_0; // @[MapT.scala 14:10]
  assign op_I_4_0_1 = I_4_0_1; // @[MapT.scala 14:10]
  assign op_I_4_1_0 = I_4_1_0; // @[MapT.scala 14:10]
  assign op_I_4_1_1 = I_4_1_1; // @[MapT.scala 14:10]
  assign op_I_5_0_0 = I_5_0_0; // @[MapT.scala 14:10]
  assign op_I_5_0_1 = I_5_0_1; // @[MapT.scala 14:10]
  assign op_I_5_1_0 = I_5_1_0; // @[MapT.scala 14:10]
  assign op_I_5_1_1 = I_5_1_1; // @[MapT.scala 14:10]
  assign op_I_6_0_0 = I_6_0_0; // @[MapT.scala 14:10]
  assign op_I_6_0_1 = I_6_0_1; // @[MapT.scala 14:10]
  assign op_I_6_1_0 = I_6_1_0; // @[MapT.scala 14:10]
  assign op_I_6_1_1 = I_6_1_1; // @[MapT.scala 14:10]
  assign op_I_7_0_0 = I_7_0_0; // @[MapT.scala 14:10]
  assign op_I_7_0_1 = I_7_0_1; // @[MapT.scala 14:10]
  assign op_I_7_1_0 = I_7_1_0; // @[MapT.scala 14:10]
  assign op_I_7_1_1 = I_7_1_1; // @[MapT.scala 14:10]
  assign op_I_8_0_0 = I_8_0_0; // @[MapT.scala 14:10]
  assign op_I_8_0_1 = I_8_0_1; // @[MapT.scala 14:10]
  assign op_I_8_1_0 = I_8_1_0; // @[MapT.scala 14:10]
  assign op_I_8_1_1 = I_8_1_1; // @[MapT.scala 14:10]
  assign op_I_9_0_0 = I_9_0_0; // @[MapT.scala 14:10]
  assign op_I_9_0_1 = I_9_0_1; // @[MapT.scala 14:10]
  assign op_I_9_1_0 = I_9_1_0; // @[MapT.scala 14:10]
  assign op_I_9_1_1 = I_9_1_1; // @[MapT.scala 14:10]
  assign op_I_10_0_0 = I_10_0_0; // @[MapT.scala 14:10]
  assign op_I_10_0_1 = I_10_0_1; // @[MapT.scala 14:10]
  assign op_I_10_1_0 = I_10_1_0; // @[MapT.scala 14:10]
  assign op_I_10_1_1 = I_10_1_1; // @[MapT.scala 14:10]
  assign op_I_11_0_0 = I_11_0_0; // @[MapT.scala 14:10]
  assign op_I_11_0_1 = I_11_0_1; // @[MapT.scala 14:10]
  assign op_I_11_1_0 = I_11_1_0; // @[MapT.scala 14:10]
  assign op_I_11_1_1 = I_11_1_1; // @[MapT.scala 14:10]
  assign op_I_12_0_0 = I_12_0_0; // @[MapT.scala 14:10]
  assign op_I_12_0_1 = I_12_0_1; // @[MapT.scala 14:10]
  assign op_I_12_1_0 = I_12_1_0; // @[MapT.scala 14:10]
  assign op_I_12_1_1 = I_12_1_1; // @[MapT.scala 14:10]
  assign op_I_13_0_0 = I_13_0_0; // @[MapT.scala 14:10]
  assign op_I_13_0_1 = I_13_0_1; // @[MapT.scala 14:10]
  assign op_I_13_1_0 = I_13_1_0; // @[MapT.scala 14:10]
  assign op_I_13_1_1 = I_13_1_1; // @[MapT.scala 14:10]
  assign op_I_14_0_0 = I_14_0_0; // @[MapT.scala 14:10]
  assign op_I_14_0_1 = I_14_0_1; // @[MapT.scala 14:10]
  assign op_I_14_1_0 = I_14_1_0; // @[MapT.scala 14:10]
  assign op_I_14_1_1 = I_14_1_1; // @[MapT.scala 14:10]
  assign op_I_15_0_0 = I_15_0_0; // @[MapT.scala 14:10]
  assign op_I_15_0_1 = I_15_0_1; // @[MapT.scala 14:10]
  assign op_I_15_1_0 = I_15_1_0; // @[MapT.scala 14:10]
  assign op_I_15_1_1 = I_15_1_1; // @[MapT.scala 14:10]
endmodule
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [7:0] I_0,
  input  [7:0] I_1,
  input  [7:0] I_2,
  input  [7:0] I_3,
  input  [7:0] I_4,
  input  [7:0] I_5,
  input  [7:0] I_6,
  input  [7:0] I_7,
  input  [7:0] I_8,
  input  [7:0] I_9,
  input  [7:0] I_10,
  input  [7:0] I_11,
  input  [7:0] I_12,
  input  [7:0] I_13,
  input  [7:0] I_14,
  input  [7:0] I_15,
  output [7:0] O_0,
  output [7:0] O_1,
  output [7:0] O_2,
  output [7:0] O_3,
  output [7:0] O_4,
  output [7:0] O_5,
  output [7:0] O_6,
  output [7:0] O_7,
  output [7:0] O_8,
  output [7:0] O_9,
  output [7:0] O_10,
  output [7:0] O_11,
  output [7:0] O_12,
  output [7:0] O_13,
  output [7:0] O_14,
  output [7:0] O_15
);
  wire  n1_clock; // @[Top.scala 74:20]
  wire  n1_reset; // @[Top.scala 74:20]
  wire  n1_valid_up; // @[Top.scala 74:20]
  wire  n1_valid_down; // @[Top.scala 74:20]
  wire [7:0] n1_I_0; // @[Top.scala 74:20]
  wire [7:0] n1_I_1; // @[Top.scala 74:20]
  wire [7:0] n1_I_2; // @[Top.scala 74:20]
  wire [7:0] n1_I_3; // @[Top.scala 74:20]
  wire [7:0] n1_I_4; // @[Top.scala 74:20]
  wire [7:0] n1_I_5; // @[Top.scala 74:20]
  wire [7:0] n1_I_6; // @[Top.scala 74:20]
  wire [7:0] n1_I_7; // @[Top.scala 74:20]
  wire [7:0] n1_I_8; // @[Top.scala 74:20]
  wire [7:0] n1_I_9; // @[Top.scala 74:20]
  wire [7:0] n1_I_10; // @[Top.scala 74:20]
  wire [7:0] n1_I_11; // @[Top.scala 74:20]
  wire [7:0] n1_I_12; // @[Top.scala 74:20]
  wire [7:0] n1_I_13; // @[Top.scala 74:20]
  wire [7:0] n1_I_14; // @[Top.scala 74:20]
  wire [7:0] n1_I_15; // @[Top.scala 74:20]
  wire [7:0] n1_O_0; // @[Top.scala 74:20]
  wire [7:0] n1_O_1; // @[Top.scala 74:20]
  wire [7:0] n1_O_2; // @[Top.scala 74:20]
  wire [7:0] n1_O_3; // @[Top.scala 74:20]
  wire [7:0] n1_O_4; // @[Top.scala 74:20]
  wire [7:0] n1_O_5; // @[Top.scala 74:20]
  wire [7:0] n1_O_6; // @[Top.scala 74:20]
  wire [7:0] n1_O_7; // @[Top.scala 74:20]
  wire [7:0] n1_O_8; // @[Top.scala 74:20]
  wire [7:0] n1_O_9; // @[Top.scala 74:20]
  wire [7:0] n1_O_10; // @[Top.scala 74:20]
  wire [7:0] n1_O_11; // @[Top.scala 74:20]
  wire [7:0] n1_O_12; // @[Top.scala 74:20]
  wire [7:0] n1_O_13; // @[Top.scala 74:20]
  wire [7:0] n1_O_14; // @[Top.scala 74:20]
  wire [7:0] n1_O_15; // @[Top.scala 74:20]
  wire  n2_clock; // @[Top.scala 77:20]
  wire  n2_reset; // @[Top.scala 77:20]
  wire  n2_valid_up; // @[Top.scala 77:20]
  wire  n2_valid_down; // @[Top.scala 77:20]
  wire [7:0] n2_I_0; // @[Top.scala 77:20]
  wire [7:0] n2_I_1; // @[Top.scala 77:20]
  wire [7:0] n2_I_2; // @[Top.scala 77:20]
  wire [7:0] n2_I_3; // @[Top.scala 77:20]
  wire [7:0] n2_I_4; // @[Top.scala 77:20]
  wire [7:0] n2_I_5; // @[Top.scala 77:20]
  wire [7:0] n2_I_6; // @[Top.scala 77:20]
  wire [7:0] n2_I_7; // @[Top.scala 77:20]
  wire [7:0] n2_I_8; // @[Top.scala 77:20]
  wire [7:0] n2_I_9; // @[Top.scala 77:20]
  wire [7:0] n2_I_10; // @[Top.scala 77:20]
  wire [7:0] n2_I_11; // @[Top.scala 77:20]
  wire [7:0] n2_I_12; // @[Top.scala 77:20]
  wire [7:0] n2_I_13; // @[Top.scala 77:20]
  wire [7:0] n2_I_14; // @[Top.scala 77:20]
  wire [7:0] n2_I_15; // @[Top.scala 77:20]
  wire [7:0] n2_O_0; // @[Top.scala 77:20]
  wire [7:0] n2_O_1; // @[Top.scala 77:20]
  wire [7:0] n2_O_2; // @[Top.scala 77:20]
  wire [7:0] n2_O_3; // @[Top.scala 77:20]
  wire [7:0] n2_O_4; // @[Top.scala 77:20]
  wire [7:0] n2_O_5; // @[Top.scala 77:20]
  wire [7:0] n2_O_6; // @[Top.scala 77:20]
  wire [7:0] n2_O_7; // @[Top.scala 77:20]
  wire [7:0] n2_O_8; // @[Top.scala 77:20]
  wire [7:0] n2_O_9; // @[Top.scala 77:20]
  wire [7:0] n2_O_10; // @[Top.scala 77:20]
  wire [7:0] n2_O_11; // @[Top.scala 77:20]
  wire [7:0] n2_O_12; // @[Top.scala 77:20]
  wire [7:0] n2_O_13; // @[Top.scala 77:20]
  wire [7:0] n2_O_14; // @[Top.scala 77:20]
  wire [7:0] n2_O_15; // @[Top.scala 77:20]
  wire  n3_clock; // @[Top.scala 80:20]
  wire  n3_reset; // @[Top.scala 80:20]
  wire  n3_valid_up; // @[Top.scala 80:20]
  wire  n3_valid_down; // @[Top.scala 80:20]
  wire [7:0] n3_I_0; // @[Top.scala 80:20]
  wire [7:0] n3_I_1; // @[Top.scala 80:20]
  wire [7:0] n3_I_2; // @[Top.scala 80:20]
  wire [7:0] n3_I_3; // @[Top.scala 80:20]
  wire [7:0] n3_I_4; // @[Top.scala 80:20]
  wire [7:0] n3_I_5; // @[Top.scala 80:20]
  wire [7:0] n3_I_6; // @[Top.scala 80:20]
  wire [7:0] n3_I_7; // @[Top.scala 80:20]
  wire [7:0] n3_I_8; // @[Top.scala 80:20]
  wire [7:0] n3_I_9; // @[Top.scala 80:20]
  wire [7:0] n3_I_10; // @[Top.scala 80:20]
  wire [7:0] n3_I_11; // @[Top.scala 80:20]
  wire [7:0] n3_I_12; // @[Top.scala 80:20]
  wire [7:0] n3_I_13; // @[Top.scala 80:20]
  wire [7:0] n3_I_14; // @[Top.scala 80:20]
  wire [7:0] n3_I_15; // @[Top.scala 80:20]
  wire [7:0] n3_O_0; // @[Top.scala 80:20]
  wire [7:0] n3_O_1; // @[Top.scala 80:20]
  wire [7:0] n3_O_2; // @[Top.scala 80:20]
  wire [7:0] n3_O_3; // @[Top.scala 80:20]
  wire [7:0] n3_O_4; // @[Top.scala 80:20]
  wire [7:0] n3_O_5; // @[Top.scala 80:20]
  wire [7:0] n3_O_6; // @[Top.scala 80:20]
  wire [7:0] n3_O_7; // @[Top.scala 80:20]
  wire [7:0] n3_O_8; // @[Top.scala 80:20]
  wire [7:0] n3_O_9; // @[Top.scala 80:20]
  wire [7:0] n3_O_10; // @[Top.scala 80:20]
  wire [7:0] n3_O_11; // @[Top.scala 80:20]
  wire [7:0] n3_O_12; // @[Top.scala 80:20]
  wire [7:0] n3_O_13; // @[Top.scala 80:20]
  wire [7:0] n3_O_14; // @[Top.scala 80:20]
  wire [7:0] n3_O_15; // @[Top.scala 80:20]
  wire  n4_clock; // @[Top.scala 83:20]
  wire  n4_valid_up; // @[Top.scala 83:20]
  wire  n4_valid_down; // @[Top.scala 83:20]
  wire [7:0] n4_I_0; // @[Top.scala 83:20]
  wire [7:0] n4_I_1; // @[Top.scala 83:20]
  wire [7:0] n4_I_2; // @[Top.scala 83:20]
  wire [7:0] n4_I_3; // @[Top.scala 83:20]
  wire [7:0] n4_I_4; // @[Top.scala 83:20]
  wire [7:0] n4_I_5; // @[Top.scala 83:20]
  wire [7:0] n4_I_6; // @[Top.scala 83:20]
  wire [7:0] n4_I_7; // @[Top.scala 83:20]
  wire [7:0] n4_I_8; // @[Top.scala 83:20]
  wire [7:0] n4_I_9; // @[Top.scala 83:20]
  wire [7:0] n4_I_10; // @[Top.scala 83:20]
  wire [7:0] n4_I_11; // @[Top.scala 83:20]
  wire [7:0] n4_I_12; // @[Top.scala 83:20]
  wire [7:0] n4_I_13; // @[Top.scala 83:20]
  wire [7:0] n4_I_14; // @[Top.scala 83:20]
  wire [7:0] n4_I_15; // @[Top.scala 83:20]
  wire [7:0] n4_O_0; // @[Top.scala 83:20]
  wire [7:0] n4_O_1; // @[Top.scala 83:20]
  wire [7:0] n4_O_2; // @[Top.scala 83:20]
  wire [7:0] n4_O_3; // @[Top.scala 83:20]
  wire [7:0] n4_O_4; // @[Top.scala 83:20]
  wire [7:0] n4_O_5; // @[Top.scala 83:20]
  wire [7:0] n4_O_6; // @[Top.scala 83:20]
  wire [7:0] n4_O_7; // @[Top.scala 83:20]
  wire [7:0] n4_O_8; // @[Top.scala 83:20]
  wire [7:0] n4_O_9; // @[Top.scala 83:20]
  wire [7:0] n4_O_10; // @[Top.scala 83:20]
  wire [7:0] n4_O_11; // @[Top.scala 83:20]
  wire [7:0] n4_O_12; // @[Top.scala 83:20]
  wire [7:0] n4_O_13; // @[Top.scala 83:20]
  wire [7:0] n4_O_14; // @[Top.scala 83:20]
  wire [7:0] n4_O_15; // @[Top.scala 83:20]
  wire  n5_clock; // @[Top.scala 86:20]
  wire  n5_valid_up; // @[Top.scala 86:20]
  wire  n5_valid_down; // @[Top.scala 86:20]
  wire [7:0] n5_I_0; // @[Top.scala 86:20]
  wire [7:0] n5_I_1; // @[Top.scala 86:20]
  wire [7:0] n5_I_2; // @[Top.scala 86:20]
  wire [7:0] n5_I_3; // @[Top.scala 86:20]
  wire [7:0] n5_I_4; // @[Top.scala 86:20]
  wire [7:0] n5_I_5; // @[Top.scala 86:20]
  wire [7:0] n5_I_6; // @[Top.scala 86:20]
  wire [7:0] n5_I_7; // @[Top.scala 86:20]
  wire [7:0] n5_I_8; // @[Top.scala 86:20]
  wire [7:0] n5_I_9; // @[Top.scala 86:20]
  wire [7:0] n5_I_10; // @[Top.scala 86:20]
  wire [7:0] n5_I_11; // @[Top.scala 86:20]
  wire [7:0] n5_I_12; // @[Top.scala 86:20]
  wire [7:0] n5_I_13; // @[Top.scala 86:20]
  wire [7:0] n5_I_14; // @[Top.scala 86:20]
  wire [7:0] n5_I_15; // @[Top.scala 86:20]
  wire [7:0] n5_O_0; // @[Top.scala 86:20]
  wire [7:0] n5_O_1; // @[Top.scala 86:20]
  wire [7:0] n5_O_2; // @[Top.scala 86:20]
  wire [7:0] n5_O_3; // @[Top.scala 86:20]
  wire [7:0] n5_O_4; // @[Top.scala 86:20]
  wire [7:0] n5_O_5; // @[Top.scala 86:20]
  wire [7:0] n5_O_6; // @[Top.scala 86:20]
  wire [7:0] n5_O_7; // @[Top.scala 86:20]
  wire [7:0] n5_O_8; // @[Top.scala 86:20]
  wire [7:0] n5_O_9; // @[Top.scala 86:20]
  wire [7:0] n5_O_10; // @[Top.scala 86:20]
  wire [7:0] n5_O_11; // @[Top.scala 86:20]
  wire [7:0] n5_O_12; // @[Top.scala 86:20]
  wire [7:0] n5_O_13; // @[Top.scala 86:20]
  wire [7:0] n5_O_14; // @[Top.scala 86:20]
  wire [7:0] n5_O_15; // @[Top.scala 86:20]
  wire  n6_valid_up; // @[Top.scala 89:20]
  wire  n6_valid_down; // @[Top.scala 89:20]
  wire [7:0] n6_I0_0; // @[Top.scala 89:20]
  wire [7:0] n6_I0_1; // @[Top.scala 89:20]
  wire [7:0] n6_I0_2; // @[Top.scala 89:20]
  wire [7:0] n6_I0_3; // @[Top.scala 89:20]
  wire [7:0] n6_I0_4; // @[Top.scala 89:20]
  wire [7:0] n6_I0_5; // @[Top.scala 89:20]
  wire [7:0] n6_I0_6; // @[Top.scala 89:20]
  wire [7:0] n6_I0_7; // @[Top.scala 89:20]
  wire [7:0] n6_I0_8; // @[Top.scala 89:20]
  wire [7:0] n6_I0_9; // @[Top.scala 89:20]
  wire [7:0] n6_I0_10; // @[Top.scala 89:20]
  wire [7:0] n6_I0_11; // @[Top.scala 89:20]
  wire [7:0] n6_I0_12; // @[Top.scala 89:20]
  wire [7:0] n6_I0_13; // @[Top.scala 89:20]
  wire [7:0] n6_I0_14; // @[Top.scala 89:20]
  wire [7:0] n6_I0_15; // @[Top.scala 89:20]
  wire [7:0] n6_I1_0; // @[Top.scala 89:20]
  wire [7:0] n6_I1_1; // @[Top.scala 89:20]
  wire [7:0] n6_I1_2; // @[Top.scala 89:20]
  wire [7:0] n6_I1_3; // @[Top.scala 89:20]
  wire [7:0] n6_I1_4; // @[Top.scala 89:20]
  wire [7:0] n6_I1_5; // @[Top.scala 89:20]
  wire [7:0] n6_I1_6; // @[Top.scala 89:20]
  wire [7:0] n6_I1_7; // @[Top.scala 89:20]
  wire [7:0] n6_I1_8; // @[Top.scala 89:20]
  wire [7:0] n6_I1_9; // @[Top.scala 89:20]
  wire [7:0] n6_I1_10; // @[Top.scala 89:20]
  wire [7:0] n6_I1_11; // @[Top.scala 89:20]
  wire [7:0] n6_I1_12; // @[Top.scala 89:20]
  wire [7:0] n6_I1_13; // @[Top.scala 89:20]
  wire [7:0] n6_I1_14; // @[Top.scala 89:20]
  wire [7:0] n6_I1_15; // @[Top.scala 89:20]
  wire [7:0] n6_O_0_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_0_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_1_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_1_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_2_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_2_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_3_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_3_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_4_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_4_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_5_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_5_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_6_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_6_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_7_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_7_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_8_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_8_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_9_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_9_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_10_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_10_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_11_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_11_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_12_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_12_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_13_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_13_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_14_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_14_1; // @[Top.scala 89:20]
  wire [7:0] n6_O_15_0; // @[Top.scala 89:20]
  wire [7:0] n6_O_15_1; // @[Top.scala 89:20]
  wire  n13_valid_up; // @[Top.scala 93:21]
  wire  n13_valid_down; // @[Top.scala 93:21]
  wire [7:0] n13_I0_0_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_0_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_1_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_1_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_2_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_2_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_3_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_3_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_4_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_4_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_5_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_5_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_6_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_6_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_7_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_7_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_8_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_8_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_9_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_9_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_10_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_10_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_11_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_11_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_12_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_12_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_13_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_13_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_14_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_14_1; // @[Top.scala 93:21]
  wire [7:0] n13_I0_15_0; // @[Top.scala 93:21]
  wire [7:0] n13_I0_15_1; // @[Top.scala 93:21]
  wire [7:0] n13_I1_0; // @[Top.scala 93:21]
  wire [7:0] n13_I1_1; // @[Top.scala 93:21]
  wire [7:0] n13_I1_2; // @[Top.scala 93:21]
  wire [7:0] n13_I1_3; // @[Top.scala 93:21]
  wire [7:0] n13_I1_4; // @[Top.scala 93:21]
  wire [7:0] n13_I1_5; // @[Top.scala 93:21]
  wire [7:0] n13_I1_6; // @[Top.scala 93:21]
  wire [7:0] n13_I1_7; // @[Top.scala 93:21]
  wire [7:0] n13_I1_8; // @[Top.scala 93:21]
  wire [7:0] n13_I1_9; // @[Top.scala 93:21]
  wire [7:0] n13_I1_10; // @[Top.scala 93:21]
  wire [7:0] n13_I1_11; // @[Top.scala 93:21]
  wire [7:0] n13_I1_12; // @[Top.scala 93:21]
  wire [7:0] n13_I1_13; // @[Top.scala 93:21]
  wire [7:0] n13_I1_14; // @[Top.scala 93:21]
  wire [7:0] n13_I1_15; // @[Top.scala 93:21]
  wire [7:0] n13_O_0_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_0_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_0_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_1_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_1_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_1_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_2_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_2_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_2_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_3_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_3_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_3_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_4_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_4_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_4_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_5_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_5_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_5_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_6_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_6_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_6_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_7_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_7_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_7_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_8_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_8_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_8_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_9_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_9_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_9_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_10_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_10_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_10_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_11_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_11_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_11_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_12_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_12_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_12_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_13_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_13_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_13_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_14_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_14_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_14_2; // @[Top.scala 93:21]
  wire [7:0] n13_O_15_0; // @[Top.scala 93:21]
  wire [7:0] n13_O_15_1; // @[Top.scala 93:21]
  wire [7:0] n13_O_15_2; // @[Top.scala 93:21]
  wire  n22_valid_up; // @[Top.scala 97:21]
  wire  n22_valid_down; // @[Top.scala 97:21]
  wire [7:0] n22_I_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_1_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_1_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_1_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_2_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_2_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_2_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_3_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_3_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_3_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_4_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_4_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_4_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_5_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_5_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_5_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_6_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_6_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_6_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_7_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_7_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_7_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_8_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_8_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_8_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_9_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_9_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_9_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_10_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_10_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_10_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_11_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_11_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_11_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_12_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_12_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_12_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_13_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_13_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_13_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_14_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_14_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_14_2; // @[Top.scala 97:21]
  wire [7:0] n22_I_15_0; // @[Top.scala 97:21]
  wire [7:0] n22_I_15_1; // @[Top.scala 97:21]
  wire [7:0] n22_I_15_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_0_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_0_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_0_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_1_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_1_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_1_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_2_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_2_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_2_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_3_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_3_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_3_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_4_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_4_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_4_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_5_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_5_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_5_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_6_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_6_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_6_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_7_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_7_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_7_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_8_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_8_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_8_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_9_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_9_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_9_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_10_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_10_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_10_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_11_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_11_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_11_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_12_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_12_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_12_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_13_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_13_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_13_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_14_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_14_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_14_0_2; // @[Top.scala 97:21]
  wire [7:0] n22_O_15_0_0; // @[Top.scala 97:21]
  wire [7:0] n22_O_15_0_1; // @[Top.scala 97:21]
  wire [7:0] n22_O_15_0_2; // @[Top.scala 97:21]
  wire  n29_valid_up; // @[Top.scala 100:21]
  wire  n29_valid_down; // @[Top.scala 100:21]
  wire [7:0] n29_I_0_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_0_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_0_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_1_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_1_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_1_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_2_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_2_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_2_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_3_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_3_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_3_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_4_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_4_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_4_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_5_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_5_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_5_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_6_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_6_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_6_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_7_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_7_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_7_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_8_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_8_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_8_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_9_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_9_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_9_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_10_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_10_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_10_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_11_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_11_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_11_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_12_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_12_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_12_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_13_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_13_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_13_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_14_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_14_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_14_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_I_15_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_I_15_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_I_15_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_0_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_0_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_0_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_1_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_1_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_1_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_2_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_2_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_2_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_3_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_3_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_3_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_4_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_4_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_4_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_5_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_5_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_5_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_6_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_6_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_6_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_7_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_7_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_7_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_8_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_8_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_8_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_9_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_9_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_9_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_10_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_10_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_10_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_11_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_11_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_11_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_12_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_12_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_12_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_13_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_13_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_13_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_14_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_14_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_14_2; // @[Top.scala 100:21]
  wire [7:0] n29_O_15_0; // @[Top.scala 100:21]
  wire [7:0] n29_O_15_1; // @[Top.scala 100:21]
  wire [7:0] n29_O_15_2; // @[Top.scala 100:21]
  wire  n30_clock; // @[Top.scala 103:21]
  wire  n30_valid_up; // @[Top.scala 103:21]
  wire  n30_valid_down; // @[Top.scala 103:21]
  wire [7:0] n30_I_0; // @[Top.scala 103:21]
  wire [7:0] n30_I_1; // @[Top.scala 103:21]
  wire [7:0] n30_I_2; // @[Top.scala 103:21]
  wire [7:0] n30_I_3; // @[Top.scala 103:21]
  wire [7:0] n30_I_4; // @[Top.scala 103:21]
  wire [7:0] n30_I_5; // @[Top.scala 103:21]
  wire [7:0] n30_I_6; // @[Top.scala 103:21]
  wire [7:0] n30_I_7; // @[Top.scala 103:21]
  wire [7:0] n30_I_8; // @[Top.scala 103:21]
  wire [7:0] n30_I_9; // @[Top.scala 103:21]
  wire [7:0] n30_I_10; // @[Top.scala 103:21]
  wire [7:0] n30_I_11; // @[Top.scala 103:21]
  wire [7:0] n30_I_12; // @[Top.scala 103:21]
  wire [7:0] n30_I_13; // @[Top.scala 103:21]
  wire [7:0] n30_I_14; // @[Top.scala 103:21]
  wire [7:0] n30_I_15; // @[Top.scala 103:21]
  wire [7:0] n30_O_0; // @[Top.scala 103:21]
  wire [7:0] n30_O_1; // @[Top.scala 103:21]
  wire [7:0] n30_O_2; // @[Top.scala 103:21]
  wire [7:0] n30_O_3; // @[Top.scala 103:21]
  wire [7:0] n30_O_4; // @[Top.scala 103:21]
  wire [7:0] n30_O_5; // @[Top.scala 103:21]
  wire [7:0] n30_O_6; // @[Top.scala 103:21]
  wire [7:0] n30_O_7; // @[Top.scala 103:21]
  wire [7:0] n30_O_8; // @[Top.scala 103:21]
  wire [7:0] n30_O_9; // @[Top.scala 103:21]
  wire [7:0] n30_O_10; // @[Top.scala 103:21]
  wire [7:0] n30_O_11; // @[Top.scala 103:21]
  wire [7:0] n30_O_12; // @[Top.scala 103:21]
  wire [7:0] n30_O_13; // @[Top.scala 103:21]
  wire [7:0] n30_O_14; // @[Top.scala 103:21]
  wire [7:0] n30_O_15; // @[Top.scala 103:21]
  wire  n31_clock; // @[Top.scala 106:21]
  wire  n31_valid_up; // @[Top.scala 106:21]
  wire  n31_valid_down; // @[Top.scala 106:21]
  wire [7:0] n31_I_0; // @[Top.scala 106:21]
  wire [7:0] n31_I_1; // @[Top.scala 106:21]
  wire [7:0] n31_I_2; // @[Top.scala 106:21]
  wire [7:0] n31_I_3; // @[Top.scala 106:21]
  wire [7:0] n31_I_4; // @[Top.scala 106:21]
  wire [7:0] n31_I_5; // @[Top.scala 106:21]
  wire [7:0] n31_I_6; // @[Top.scala 106:21]
  wire [7:0] n31_I_7; // @[Top.scala 106:21]
  wire [7:0] n31_I_8; // @[Top.scala 106:21]
  wire [7:0] n31_I_9; // @[Top.scala 106:21]
  wire [7:0] n31_I_10; // @[Top.scala 106:21]
  wire [7:0] n31_I_11; // @[Top.scala 106:21]
  wire [7:0] n31_I_12; // @[Top.scala 106:21]
  wire [7:0] n31_I_13; // @[Top.scala 106:21]
  wire [7:0] n31_I_14; // @[Top.scala 106:21]
  wire [7:0] n31_I_15; // @[Top.scala 106:21]
  wire [7:0] n31_O_0; // @[Top.scala 106:21]
  wire [7:0] n31_O_1; // @[Top.scala 106:21]
  wire [7:0] n31_O_2; // @[Top.scala 106:21]
  wire [7:0] n31_O_3; // @[Top.scala 106:21]
  wire [7:0] n31_O_4; // @[Top.scala 106:21]
  wire [7:0] n31_O_5; // @[Top.scala 106:21]
  wire [7:0] n31_O_6; // @[Top.scala 106:21]
  wire [7:0] n31_O_7; // @[Top.scala 106:21]
  wire [7:0] n31_O_8; // @[Top.scala 106:21]
  wire [7:0] n31_O_9; // @[Top.scala 106:21]
  wire [7:0] n31_O_10; // @[Top.scala 106:21]
  wire [7:0] n31_O_11; // @[Top.scala 106:21]
  wire [7:0] n31_O_12; // @[Top.scala 106:21]
  wire [7:0] n31_O_13; // @[Top.scala 106:21]
  wire [7:0] n31_O_14; // @[Top.scala 106:21]
  wire [7:0] n31_O_15; // @[Top.scala 106:21]
  wire  n32_valid_up; // @[Top.scala 109:21]
  wire  n32_valid_down; // @[Top.scala 109:21]
  wire [7:0] n32_I0_0; // @[Top.scala 109:21]
  wire [7:0] n32_I0_1; // @[Top.scala 109:21]
  wire [7:0] n32_I0_2; // @[Top.scala 109:21]
  wire [7:0] n32_I0_3; // @[Top.scala 109:21]
  wire [7:0] n32_I0_4; // @[Top.scala 109:21]
  wire [7:0] n32_I0_5; // @[Top.scala 109:21]
  wire [7:0] n32_I0_6; // @[Top.scala 109:21]
  wire [7:0] n32_I0_7; // @[Top.scala 109:21]
  wire [7:0] n32_I0_8; // @[Top.scala 109:21]
  wire [7:0] n32_I0_9; // @[Top.scala 109:21]
  wire [7:0] n32_I0_10; // @[Top.scala 109:21]
  wire [7:0] n32_I0_11; // @[Top.scala 109:21]
  wire [7:0] n32_I0_12; // @[Top.scala 109:21]
  wire [7:0] n32_I0_13; // @[Top.scala 109:21]
  wire [7:0] n32_I0_14; // @[Top.scala 109:21]
  wire [7:0] n32_I0_15; // @[Top.scala 109:21]
  wire [7:0] n32_I1_0; // @[Top.scala 109:21]
  wire [7:0] n32_I1_1; // @[Top.scala 109:21]
  wire [7:0] n32_I1_2; // @[Top.scala 109:21]
  wire [7:0] n32_I1_3; // @[Top.scala 109:21]
  wire [7:0] n32_I1_4; // @[Top.scala 109:21]
  wire [7:0] n32_I1_5; // @[Top.scala 109:21]
  wire [7:0] n32_I1_6; // @[Top.scala 109:21]
  wire [7:0] n32_I1_7; // @[Top.scala 109:21]
  wire [7:0] n32_I1_8; // @[Top.scala 109:21]
  wire [7:0] n32_I1_9; // @[Top.scala 109:21]
  wire [7:0] n32_I1_10; // @[Top.scala 109:21]
  wire [7:0] n32_I1_11; // @[Top.scala 109:21]
  wire [7:0] n32_I1_12; // @[Top.scala 109:21]
  wire [7:0] n32_I1_13; // @[Top.scala 109:21]
  wire [7:0] n32_I1_14; // @[Top.scala 109:21]
  wire [7:0] n32_I1_15; // @[Top.scala 109:21]
  wire [7:0] n32_O_0_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_0_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_1_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_1_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_2_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_2_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_3_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_3_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_4_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_4_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_5_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_5_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_6_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_6_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_7_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_7_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_8_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_8_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_9_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_9_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_10_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_10_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_11_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_11_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_12_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_12_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_13_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_13_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_14_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_14_1; // @[Top.scala 109:21]
  wire [7:0] n32_O_15_0; // @[Top.scala 109:21]
  wire [7:0] n32_O_15_1; // @[Top.scala 109:21]
  wire  n39_valid_up; // @[Top.scala 113:21]
  wire  n39_valid_down; // @[Top.scala 113:21]
  wire [7:0] n39_I0_0_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_0_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_1_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_1_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_2_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_2_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_3_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_3_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_4_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_4_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_5_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_5_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_6_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_6_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_7_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_7_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_8_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_8_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_9_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_9_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_10_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_10_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_11_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_11_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_12_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_12_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_13_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_13_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_14_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_14_1; // @[Top.scala 113:21]
  wire [7:0] n39_I0_15_0; // @[Top.scala 113:21]
  wire [7:0] n39_I0_15_1; // @[Top.scala 113:21]
  wire [7:0] n39_I1_0; // @[Top.scala 113:21]
  wire [7:0] n39_I1_1; // @[Top.scala 113:21]
  wire [7:0] n39_I1_2; // @[Top.scala 113:21]
  wire [7:0] n39_I1_3; // @[Top.scala 113:21]
  wire [7:0] n39_I1_4; // @[Top.scala 113:21]
  wire [7:0] n39_I1_5; // @[Top.scala 113:21]
  wire [7:0] n39_I1_6; // @[Top.scala 113:21]
  wire [7:0] n39_I1_7; // @[Top.scala 113:21]
  wire [7:0] n39_I1_8; // @[Top.scala 113:21]
  wire [7:0] n39_I1_9; // @[Top.scala 113:21]
  wire [7:0] n39_I1_10; // @[Top.scala 113:21]
  wire [7:0] n39_I1_11; // @[Top.scala 113:21]
  wire [7:0] n39_I1_12; // @[Top.scala 113:21]
  wire [7:0] n39_I1_13; // @[Top.scala 113:21]
  wire [7:0] n39_I1_14; // @[Top.scala 113:21]
  wire [7:0] n39_I1_15; // @[Top.scala 113:21]
  wire [7:0] n39_O_0_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_0_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_0_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_1_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_1_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_1_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_2_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_2_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_2_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_3_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_3_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_3_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_4_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_4_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_4_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_5_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_5_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_5_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_6_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_6_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_6_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_7_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_7_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_7_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_8_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_8_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_8_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_9_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_9_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_9_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_10_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_10_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_10_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_11_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_11_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_11_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_12_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_12_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_12_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_13_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_13_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_13_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_14_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_14_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_14_2; // @[Top.scala 113:21]
  wire [7:0] n39_O_15_0; // @[Top.scala 113:21]
  wire [7:0] n39_O_15_1; // @[Top.scala 113:21]
  wire [7:0] n39_O_15_2; // @[Top.scala 113:21]
  wire  n48_valid_up; // @[Top.scala 117:21]
  wire  n48_valid_down; // @[Top.scala 117:21]
  wire [7:0] n48_I_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_1_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_1_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_1_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_2_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_2_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_2_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_3_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_3_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_3_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_4_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_4_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_4_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_5_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_5_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_5_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_6_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_6_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_6_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_7_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_7_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_7_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_8_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_8_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_8_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_9_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_9_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_9_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_10_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_10_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_10_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_11_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_11_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_11_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_12_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_12_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_12_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_13_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_13_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_13_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_14_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_14_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_14_2; // @[Top.scala 117:21]
  wire [7:0] n48_I_15_0; // @[Top.scala 117:21]
  wire [7:0] n48_I_15_1; // @[Top.scala 117:21]
  wire [7:0] n48_I_15_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_0_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_0_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_0_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_1_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_1_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_1_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_2_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_2_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_2_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_3_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_3_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_3_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_4_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_4_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_4_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_5_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_5_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_5_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_6_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_6_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_6_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_7_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_7_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_7_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_8_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_8_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_8_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_9_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_9_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_9_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_10_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_10_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_10_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_11_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_11_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_11_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_12_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_12_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_12_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_13_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_13_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_13_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_14_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_14_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_14_0_2; // @[Top.scala 117:21]
  wire [7:0] n48_O_15_0_0; // @[Top.scala 117:21]
  wire [7:0] n48_O_15_0_1; // @[Top.scala 117:21]
  wire [7:0] n48_O_15_0_2; // @[Top.scala 117:21]
  wire  n55_valid_up; // @[Top.scala 120:21]
  wire  n55_valid_down; // @[Top.scala 120:21]
  wire [7:0] n55_I_0_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_0_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_0_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_1_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_1_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_1_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_2_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_2_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_2_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_3_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_3_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_3_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_4_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_4_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_4_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_5_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_5_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_5_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_6_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_6_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_6_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_7_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_7_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_7_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_8_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_8_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_8_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_9_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_9_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_9_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_10_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_10_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_10_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_11_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_11_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_11_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_12_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_12_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_12_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_13_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_13_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_13_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_14_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_14_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_14_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_I_15_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_I_15_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_I_15_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_0_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_0_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_0_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_1_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_1_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_1_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_2_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_2_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_2_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_3_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_3_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_3_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_4_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_4_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_4_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_5_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_5_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_5_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_6_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_6_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_6_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_7_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_7_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_7_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_8_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_8_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_8_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_9_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_9_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_9_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_10_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_10_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_10_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_11_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_11_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_11_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_12_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_12_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_12_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_13_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_13_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_13_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_14_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_14_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_14_2; // @[Top.scala 120:21]
  wire [7:0] n55_O_15_0; // @[Top.scala 120:21]
  wire [7:0] n55_O_15_1; // @[Top.scala 120:21]
  wire [7:0] n55_O_15_2; // @[Top.scala 120:21]
  wire  n56_valid_up; // @[Top.scala 123:21]
  wire  n56_valid_down; // @[Top.scala 123:21]
  wire [7:0] n56_I0_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_2_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_2_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_2_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_3_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_3_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_3_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_4_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_4_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_4_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_5_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_5_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_5_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_6_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_6_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_6_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_7_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_7_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_7_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_8_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_8_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_8_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_9_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_9_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_9_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_10_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_10_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_10_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_11_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_11_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_11_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_12_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_12_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_12_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_13_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_13_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_13_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_14_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_14_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_14_2; // @[Top.scala 123:21]
  wire [7:0] n56_I0_15_0; // @[Top.scala 123:21]
  wire [7:0] n56_I0_15_1; // @[Top.scala 123:21]
  wire [7:0] n56_I0_15_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_2_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_2_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_2_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_3_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_3_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_3_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_4_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_4_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_4_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_5_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_5_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_5_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_6_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_6_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_6_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_7_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_7_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_7_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_8_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_8_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_8_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_9_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_9_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_9_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_10_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_10_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_10_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_11_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_11_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_11_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_12_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_12_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_12_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_13_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_13_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_13_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_14_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_14_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_14_2; // @[Top.scala 123:21]
  wire [7:0] n56_I1_15_0; // @[Top.scala 123:21]
  wire [7:0] n56_I1_15_1; // @[Top.scala 123:21]
  wire [7:0] n56_I1_15_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_0_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_0_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_0_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_0_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_0_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_0_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_1_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_1_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_1_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_1_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_1_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_1_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_2_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_2_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_2_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_2_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_2_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_2_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_3_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_3_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_3_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_3_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_3_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_3_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_4_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_4_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_4_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_4_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_4_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_4_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_5_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_5_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_5_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_5_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_5_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_5_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_6_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_6_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_6_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_6_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_6_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_6_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_7_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_7_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_7_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_7_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_7_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_7_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_8_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_8_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_8_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_8_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_8_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_8_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_9_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_9_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_9_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_9_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_9_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_9_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_10_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_10_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_10_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_10_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_10_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_10_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_11_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_11_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_11_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_11_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_11_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_11_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_12_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_12_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_12_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_12_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_12_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_12_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_13_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_13_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_13_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_13_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_13_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_13_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_14_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_14_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_14_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_14_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_14_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_14_1_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_15_0_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_15_0_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_15_0_2; // @[Top.scala 123:21]
  wire [7:0] n56_O_15_1_0; // @[Top.scala 123:21]
  wire [7:0] n56_O_15_1_1; // @[Top.scala 123:21]
  wire [7:0] n56_O_15_1_2; // @[Top.scala 123:21]
  wire  n63_clock; // @[Top.scala 127:21]
  wire  n63_valid_up; // @[Top.scala 127:21]
  wire  n63_valid_down; // @[Top.scala 127:21]
  wire [7:0] n63_I_0; // @[Top.scala 127:21]
  wire [7:0] n63_I_1; // @[Top.scala 127:21]
  wire [7:0] n63_I_2; // @[Top.scala 127:21]
  wire [7:0] n63_I_3; // @[Top.scala 127:21]
  wire [7:0] n63_I_4; // @[Top.scala 127:21]
  wire [7:0] n63_I_5; // @[Top.scala 127:21]
  wire [7:0] n63_I_6; // @[Top.scala 127:21]
  wire [7:0] n63_I_7; // @[Top.scala 127:21]
  wire [7:0] n63_I_8; // @[Top.scala 127:21]
  wire [7:0] n63_I_9; // @[Top.scala 127:21]
  wire [7:0] n63_I_10; // @[Top.scala 127:21]
  wire [7:0] n63_I_11; // @[Top.scala 127:21]
  wire [7:0] n63_I_12; // @[Top.scala 127:21]
  wire [7:0] n63_I_13; // @[Top.scala 127:21]
  wire [7:0] n63_I_14; // @[Top.scala 127:21]
  wire [7:0] n63_I_15; // @[Top.scala 127:21]
  wire [7:0] n63_O_0; // @[Top.scala 127:21]
  wire [7:0] n63_O_1; // @[Top.scala 127:21]
  wire [7:0] n63_O_2; // @[Top.scala 127:21]
  wire [7:0] n63_O_3; // @[Top.scala 127:21]
  wire [7:0] n63_O_4; // @[Top.scala 127:21]
  wire [7:0] n63_O_5; // @[Top.scala 127:21]
  wire [7:0] n63_O_6; // @[Top.scala 127:21]
  wire [7:0] n63_O_7; // @[Top.scala 127:21]
  wire [7:0] n63_O_8; // @[Top.scala 127:21]
  wire [7:0] n63_O_9; // @[Top.scala 127:21]
  wire [7:0] n63_O_10; // @[Top.scala 127:21]
  wire [7:0] n63_O_11; // @[Top.scala 127:21]
  wire [7:0] n63_O_12; // @[Top.scala 127:21]
  wire [7:0] n63_O_13; // @[Top.scala 127:21]
  wire [7:0] n63_O_14; // @[Top.scala 127:21]
  wire [7:0] n63_O_15; // @[Top.scala 127:21]
  wire  n64_clock; // @[Top.scala 130:21]
  wire  n64_valid_up; // @[Top.scala 130:21]
  wire  n64_valid_down; // @[Top.scala 130:21]
  wire [7:0] n64_I_0; // @[Top.scala 130:21]
  wire [7:0] n64_I_1; // @[Top.scala 130:21]
  wire [7:0] n64_I_2; // @[Top.scala 130:21]
  wire [7:0] n64_I_3; // @[Top.scala 130:21]
  wire [7:0] n64_I_4; // @[Top.scala 130:21]
  wire [7:0] n64_I_5; // @[Top.scala 130:21]
  wire [7:0] n64_I_6; // @[Top.scala 130:21]
  wire [7:0] n64_I_7; // @[Top.scala 130:21]
  wire [7:0] n64_I_8; // @[Top.scala 130:21]
  wire [7:0] n64_I_9; // @[Top.scala 130:21]
  wire [7:0] n64_I_10; // @[Top.scala 130:21]
  wire [7:0] n64_I_11; // @[Top.scala 130:21]
  wire [7:0] n64_I_12; // @[Top.scala 130:21]
  wire [7:0] n64_I_13; // @[Top.scala 130:21]
  wire [7:0] n64_I_14; // @[Top.scala 130:21]
  wire [7:0] n64_I_15; // @[Top.scala 130:21]
  wire [7:0] n64_O_0; // @[Top.scala 130:21]
  wire [7:0] n64_O_1; // @[Top.scala 130:21]
  wire [7:0] n64_O_2; // @[Top.scala 130:21]
  wire [7:0] n64_O_3; // @[Top.scala 130:21]
  wire [7:0] n64_O_4; // @[Top.scala 130:21]
  wire [7:0] n64_O_5; // @[Top.scala 130:21]
  wire [7:0] n64_O_6; // @[Top.scala 130:21]
  wire [7:0] n64_O_7; // @[Top.scala 130:21]
  wire [7:0] n64_O_8; // @[Top.scala 130:21]
  wire [7:0] n64_O_9; // @[Top.scala 130:21]
  wire [7:0] n64_O_10; // @[Top.scala 130:21]
  wire [7:0] n64_O_11; // @[Top.scala 130:21]
  wire [7:0] n64_O_12; // @[Top.scala 130:21]
  wire [7:0] n64_O_13; // @[Top.scala 130:21]
  wire [7:0] n64_O_14; // @[Top.scala 130:21]
  wire [7:0] n64_O_15; // @[Top.scala 130:21]
  wire  n65_valid_up; // @[Top.scala 133:21]
  wire  n65_valid_down; // @[Top.scala 133:21]
  wire [7:0] n65_I0_0; // @[Top.scala 133:21]
  wire [7:0] n65_I0_1; // @[Top.scala 133:21]
  wire [7:0] n65_I0_2; // @[Top.scala 133:21]
  wire [7:0] n65_I0_3; // @[Top.scala 133:21]
  wire [7:0] n65_I0_4; // @[Top.scala 133:21]
  wire [7:0] n65_I0_5; // @[Top.scala 133:21]
  wire [7:0] n65_I0_6; // @[Top.scala 133:21]
  wire [7:0] n65_I0_7; // @[Top.scala 133:21]
  wire [7:0] n65_I0_8; // @[Top.scala 133:21]
  wire [7:0] n65_I0_9; // @[Top.scala 133:21]
  wire [7:0] n65_I0_10; // @[Top.scala 133:21]
  wire [7:0] n65_I0_11; // @[Top.scala 133:21]
  wire [7:0] n65_I0_12; // @[Top.scala 133:21]
  wire [7:0] n65_I0_13; // @[Top.scala 133:21]
  wire [7:0] n65_I0_14; // @[Top.scala 133:21]
  wire [7:0] n65_I0_15; // @[Top.scala 133:21]
  wire [7:0] n65_I1_0; // @[Top.scala 133:21]
  wire [7:0] n65_I1_1; // @[Top.scala 133:21]
  wire [7:0] n65_I1_2; // @[Top.scala 133:21]
  wire [7:0] n65_I1_3; // @[Top.scala 133:21]
  wire [7:0] n65_I1_4; // @[Top.scala 133:21]
  wire [7:0] n65_I1_5; // @[Top.scala 133:21]
  wire [7:0] n65_I1_6; // @[Top.scala 133:21]
  wire [7:0] n65_I1_7; // @[Top.scala 133:21]
  wire [7:0] n65_I1_8; // @[Top.scala 133:21]
  wire [7:0] n65_I1_9; // @[Top.scala 133:21]
  wire [7:0] n65_I1_10; // @[Top.scala 133:21]
  wire [7:0] n65_I1_11; // @[Top.scala 133:21]
  wire [7:0] n65_I1_12; // @[Top.scala 133:21]
  wire [7:0] n65_I1_13; // @[Top.scala 133:21]
  wire [7:0] n65_I1_14; // @[Top.scala 133:21]
  wire [7:0] n65_I1_15; // @[Top.scala 133:21]
  wire [7:0] n65_O_0_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_0_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_1_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_1_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_2_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_2_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_3_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_3_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_4_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_4_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_5_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_5_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_6_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_6_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_7_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_7_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_8_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_8_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_9_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_9_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_10_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_10_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_11_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_11_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_12_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_12_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_13_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_13_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_14_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_14_1; // @[Top.scala 133:21]
  wire [7:0] n65_O_15_0; // @[Top.scala 133:21]
  wire [7:0] n65_O_15_1; // @[Top.scala 133:21]
  wire  n72_valid_up; // @[Top.scala 137:21]
  wire  n72_valid_down; // @[Top.scala 137:21]
  wire [7:0] n72_I0_0_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_0_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_1_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_1_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_2_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_2_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_3_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_3_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_4_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_4_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_5_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_5_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_6_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_6_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_7_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_7_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_8_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_8_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_9_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_9_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_10_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_10_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_11_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_11_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_12_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_12_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_13_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_13_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_14_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_14_1; // @[Top.scala 137:21]
  wire [7:0] n72_I0_15_0; // @[Top.scala 137:21]
  wire [7:0] n72_I0_15_1; // @[Top.scala 137:21]
  wire [7:0] n72_I1_0; // @[Top.scala 137:21]
  wire [7:0] n72_I1_1; // @[Top.scala 137:21]
  wire [7:0] n72_I1_2; // @[Top.scala 137:21]
  wire [7:0] n72_I1_3; // @[Top.scala 137:21]
  wire [7:0] n72_I1_4; // @[Top.scala 137:21]
  wire [7:0] n72_I1_5; // @[Top.scala 137:21]
  wire [7:0] n72_I1_6; // @[Top.scala 137:21]
  wire [7:0] n72_I1_7; // @[Top.scala 137:21]
  wire [7:0] n72_I1_8; // @[Top.scala 137:21]
  wire [7:0] n72_I1_9; // @[Top.scala 137:21]
  wire [7:0] n72_I1_10; // @[Top.scala 137:21]
  wire [7:0] n72_I1_11; // @[Top.scala 137:21]
  wire [7:0] n72_I1_12; // @[Top.scala 137:21]
  wire [7:0] n72_I1_13; // @[Top.scala 137:21]
  wire [7:0] n72_I1_14; // @[Top.scala 137:21]
  wire [7:0] n72_I1_15; // @[Top.scala 137:21]
  wire [7:0] n72_O_0_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_0_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_0_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_1_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_1_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_1_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_2_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_2_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_2_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_3_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_3_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_3_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_4_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_4_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_4_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_5_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_5_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_5_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_6_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_6_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_6_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_7_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_7_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_7_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_8_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_8_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_8_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_9_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_9_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_9_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_10_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_10_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_10_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_11_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_11_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_11_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_12_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_12_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_12_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_13_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_13_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_13_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_14_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_14_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_14_2; // @[Top.scala 137:21]
  wire [7:0] n72_O_15_0; // @[Top.scala 137:21]
  wire [7:0] n72_O_15_1; // @[Top.scala 137:21]
  wire [7:0] n72_O_15_2; // @[Top.scala 137:21]
  wire  n81_valid_up; // @[Top.scala 141:21]
  wire  n81_valid_down; // @[Top.scala 141:21]
  wire [7:0] n81_I_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_1_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_1_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_1_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_2_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_2_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_2_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_3_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_3_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_3_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_4_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_4_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_4_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_5_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_5_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_5_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_6_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_6_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_6_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_7_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_7_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_7_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_8_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_8_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_8_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_9_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_9_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_9_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_10_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_10_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_10_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_11_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_11_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_11_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_12_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_12_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_12_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_13_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_13_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_13_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_14_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_14_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_14_2; // @[Top.scala 141:21]
  wire [7:0] n81_I_15_0; // @[Top.scala 141:21]
  wire [7:0] n81_I_15_1; // @[Top.scala 141:21]
  wire [7:0] n81_I_15_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_0_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_0_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_0_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_1_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_1_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_1_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_2_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_2_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_2_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_3_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_3_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_3_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_4_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_4_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_4_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_5_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_5_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_5_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_6_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_6_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_6_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_7_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_7_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_7_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_8_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_8_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_8_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_9_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_9_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_9_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_10_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_10_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_10_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_11_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_11_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_11_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_12_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_12_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_12_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_13_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_13_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_13_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_14_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_14_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_14_0_2; // @[Top.scala 141:21]
  wire [7:0] n81_O_15_0_0; // @[Top.scala 141:21]
  wire [7:0] n81_O_15_0_1; // @[Top.scala 141:21]
  wire [7:0] n81_O_15_0_2; // @[Top.scala 141:21]
  wire  n88_valid_up; // @[Top.scala 144:21]
  wire  n88_valid_down; // @[Top.scala 144:21]
  wire [7:0] n88_I_0_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_0_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_0_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_1_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_1_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_1_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_2_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_2_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_2_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_3_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_3_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_3_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_4_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_4_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_4_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_5_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_5_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_5_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_6_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_6_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_6_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_7_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_7_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_7_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_8_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_8_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_8_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_9_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_9_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_9_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_10_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_10_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_10_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_11_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_11_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_11_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_12_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_12_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_12_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_13_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_13_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_13_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_14_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_14_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_14_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_I_15_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_I_15_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_I_15_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_0_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_0_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_0_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_1_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_1_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_1_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_2_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_2_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_2_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_3_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_3_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_3_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_4_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_4_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_4_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_5_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_5_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_5_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_6_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_6_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_6_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_7_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_7_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_7_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_8_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_8_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_8_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_9_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_9_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_9_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_10_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_10_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_10_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_11_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_11_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_11_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_12_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_12_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_12_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_13_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_13_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_13_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_14_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_14_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_14_2; // @[Top.scala 144:21]
  wire [7:0] n88_O_15_0; // @[Top.scala 144:21]
  wire [7:0] n88_O_15_1; // @[Top.scala 144:21]
  wire [7:0] n88_O_15_2; // @[Top.scala 144:21]
  wire  n89_valid_up; // @[Top.scala 147:21]
  wire  n89_valid_down; // @[Top.scala 147:21]
  wire [7:0] n89_I0_0_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_0_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_0_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_0_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_0_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_0_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_1_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_1_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_1_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_1_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_1_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_1_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_2_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_2_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_2_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_2_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_2_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_2_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_3_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_3_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_3_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_3_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_3_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_3_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_4_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_4_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_4_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_4_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_4_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_4_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_5_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_5_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_5_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_5_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_5_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_5_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_6_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_6_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_6_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_6_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_6_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_6_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_7_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_7_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_7_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_7_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_7_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_7_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_8_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_8_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_8_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_8_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_8_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_8_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_9_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_9_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_9_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_9_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_9_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_9_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_10_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_10_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_10_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_10_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_10_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_10_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_11_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_11_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_11_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_11_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_11_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_11_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_12_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_12_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_12_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_12_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_12_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_12_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_13_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_13_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_13_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_13_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_13_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_13_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_14_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_14_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_14_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_14_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_14_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_14_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_15_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_15_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_15_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I0_15_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I0_15_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I0_15_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_3_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_3_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_3_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_4_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_4_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_4_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_5_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_5_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_5_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_6_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_6_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_6_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_7_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_7_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_7_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_8_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_8_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_8_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_9_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_9_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_9_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_10_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_10_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_10_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_11_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_11_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_11_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_12_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_12_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_12_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_13_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_13_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_13_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_14_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_14_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_14_2; // @[Top.scala 147:21]
  wire [7:0] n89_I1_15_0; // @[Top.scala 147:21]
  wire [7:0] n89_I1_15_1; // @[Top.scala 147:21]
  wire [7:0] n89_I1_15_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_0_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_1_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_2_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_3_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_4_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_5_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_6_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_7_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_8_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_9_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_10_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_11_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_12_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_13_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_14_2_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_0_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_0_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_0_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_1_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_1_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_1_2; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_2_0; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_2_1; // @[Top.scala 147:21]
  wire [7:0] n89_O_15_2_2; // @[Top.scala 147:21]
  wire  n98_valid_up; // @[Top.scala 151:21]
  wire  n98_valid_down; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_1_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_2_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_3_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_4_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_5_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_6_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_7_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_8_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_9_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_10_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_11_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_12_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_13_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_14_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_I_15_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_0_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_1_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_2_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_3_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_4_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_5_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_6_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_7_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_8_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_9_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_10_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_11_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_12_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_13_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_14_0_2_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_0_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_0_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_0_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_1_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_1_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_1_2; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_2_0; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_2_1; // @[Top.scala 151:21]
  wire [7:0] n98_O_15_0_2_2; // @[Top.scala 151:21]
  wire  n105_valid_up; // @[Top.scala 154:22]
  wire  n105_valid_down; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_0_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_1_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_2_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_3_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_4_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_5_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_6_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_7_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_8_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_9_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_10_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_11_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_12_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_13_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_14_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_I_15_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_0_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_1_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_2_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_3_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_4_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_5_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_6_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_7_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_8_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_9_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_10_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_11_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_12_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_13_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_14_2_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_0_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_0_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_0_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_1_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_1_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_1_2; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_2_0; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_2_1; // @[Top.scala 154:22]
  wire [7:0] n105_O_15_2_2; // @[Top.scala 154:22]
  wire  n147_clock; // @[Top.scala 157:22]
  wire  n147_reset; // @[Top.scala 157:22]
  wire  n147_valid_up; // @[Top.scala 157:22]
  wire  n147_valid_down; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_0_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_1_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_2_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_3_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_4_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_5_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_6_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_7_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_8_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_9_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_10_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_11_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_12_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_13_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_14_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_0_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_0_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_1_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_1_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_1_2; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_2_0; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_2_1; // @[Top.scala 157:22]
  wire [7:0] n147_I_15_2_2; // @[Top.scala 157:22]
  wire [7:0] n147_O_0_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_1_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_2_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_3_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_4_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_5_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_6_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_7_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_8_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_9_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_10_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_11_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_12_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_13_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_14_0_0; // @[Top.scala 157:22]
  wire [7:0] n147_O_15_0_0; // @[Top.scala 157:22]
  wire  n148_valid_up; // @[Top.scala 160:22]
  wire  n148_valid_down; // @[Top.scala 160:22]
  wire [7:0] n148_I_0_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_1_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_2_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_3_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_4_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_5_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_6_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_7_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_8_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_9_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_10_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_11_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_12_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_13_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_14_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_I_15_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_0_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_1_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_2_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_3_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_4_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_5_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_6_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_7_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_8_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_9_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_10_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_11_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_12_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_13_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_14_0; // @[Top.scala 160:22]
  wire [7:0] n148_O_15_0; // @[Top.scala 160:22]
  wire  n149_valid_up; // @[Top.scala 163:22]
  wire  n149_valid_down; // @[Top.scala 163:22]
  wire [7:0] n149_I_0_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_1_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_2_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_3_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_4_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_5_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_6_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_7_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_8_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_9_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_10_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_11_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_12_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_13_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_14_0; // @[Top.scala 163:22]
  wire [7:0] n149_I_15_0; // @[Top.scala 163:22]
  wire [7:0] n149_O_0; // @[Top.scala 163:22]
  wire [7:0] n149_O_1; // @[Top.scala 163:22]
  wire [7:0] n149_O_2; // @[Top.scala 163:22]
  wire [7:0] n149_O_3; // @[Top.scala 163:22]
  wire [7:0] n149_O_4; // @[Top.scala 163:22]
  wire [7:0] n149_O_5; // @[Top.scala 163:22]
  wire [7:0] n149_O_6; // @[Top.scala 163:22]
  wire [7:0] n149_O_7; // @[Top.scala 163:22]
  wire [7:0] n149_O_8; // @[Top.scala 163:22]
  wire [7:0] n149_O_9; // @[Top.scala 163:22]
  wire [7:0] n149_O_10; // @[Top.scala 163:22]
  wire [7:0] n149_O_11; // @[Top.scala 163:22]
  wire [7:0] n149_O_12; // @[Top.scala 163:22]
  wire [7:0] n149_O_13; // @[Top.scala 163:22]
  wire [7:0] n149_O_14; // @[Top.scala 163:22]
  wire [7:0] n149_O_15; // @[Top.scala 163:22]
  wire  n150_clock; // @[Top.scala 166:22]
  wire  n150_reset; // @[Top.scala 166:22]
  wire  n150_valid_up; // @[Top.scala 166:22]
  wire  n150_valid_down; // @[Top.scala 166:22]
  wire [7:0] n150_I_0; // @[Top.scala 166:22]
  wire [7:0] n150_I_1; // @[Top.scala 166:22]
  wire [7:0] n150_I_2; // @[Top.scala 166:22]
  wire [7:0] n150_I_3; // @[Top.scala 166:22]
  wire [7:0] n150_I_4; // @[Top.scala 166:22]
  wire [7:0] n150_I_5; // @[Top.scala 166:22]
  wire [7:0] n150_I_6; // @[Top.scala 166:22]
  wire [7:0] n150_I_7; // @[Top.scala 166:22]
  wire [7:0] n150_I_8; // @[Top.scala 166:22]
  wire [7:0] n150_I_9; // @[Top.scala 166:22]
  wire [7:0] n150_I_10; // @[Top.scala 166:22]
  wire [7:0] n150_I_11; // @[Top.scala 166:22]
  wire [7:0] n150_I_12; // @[Top.scala 166:22]
  wire [7:0] n150_I_13; // @[Top.scala 166:22]
  wire [7:0] n150_I_14; // @[Top.scala 166:22]
  wire [7:0] n150_I_15; // @[Top.scala 166:22]
  wire [7:0] n150_O_0; // @[Top.scala 166:22]
  wire [7:0] n150_O_1; // @[Top.scala 166:22]
  wire [7:0] n150_O_2; // @[Top.scala 166:22]
  wire [7:0] n150_O_3; // @[Top.scala 166:22]
  wire [7:0] n150_O_4; // @[Top.scala 166:22]
  wire [7:0] n150_O_5; // @[Top.scala 166:22]
  wire [7:0] n150_O_6; // @[Top.scala 166:22]
  wire [7:0] n150_O_7; // @[Top.scala 166:22]
  wire [7:0] n150_O_8; // @[Top.scala 166:22]
  wire [7:0] n150_O_9; // @[Top.scala 166:22]
  wire [7:0] n150_O_10; // @[Top.scala 166:22]
  wire [7:0] n150_O_11; // @[Top.scala 166:22]
  wire [7:0] n150_O_12; // @[Top.scala 166:22]
  wire [7:0] n150_O_13; // @[Top.scala 166:22]
  wire [7:0] n150_O_14; // @[Top.scala 166:22]
  wire [7:0] n150_O_15; // @[Top.scala 166:22]
  wire  n151_clock; // @[Top.scala 169:22]
  wire  n151_valid_up; // @[Top.scala 169:22]
  wire  n151_valid_down; // @[Top.scala 169:22]
  wire [7:0] n151_I_0; // @[Top.scala 169:22]
  wire [7:0] n151_I_1; // @[Top.scala 169:22]
  wire [7:0] n151_I_2; // @[Top.scala 169:22]
  wire [7:0] n151_I_3; // @[Top.scala 169:22]
  wire [7:0] n151_I_4; // @[Top.scala 169:22]
  wire [7:0] n151_I_5; // @[Top.scala 169:22]
  wire [7:0] n151_I_6; // @[Top.scala 169:22]
  wire [7:0] n151_I_7; // @[Top.scala 169:22]
  wire [7:0] n151_I_8; // @[Top.scala 169:22]
  wire [7:0] n151_I_9; // @[Top.scala 169:22]
  wire [7:0] n151_I_10; // @[Top.scala 169:22]
  wire [7:0] n151_I_11; // @[Top.scala 169:22]
  wire [7:0] n151_I_12; // @[Top.scala 169:22]
  wire [7:0] n151_I_13; // @[Top.scala 169:22]
  wire [7:0] n151_I_14; // @[Top.scala 169:22]
  wire [7:0] n151_I_15; // @[Top.scala 169:22]
  wire [7:0] n151_O_0; // @[Top.scala 169:22]
  wire [7:0] n151_O_1; // @[Top.scala 169:22]
  wire [7:0] n151_O_2; // @[Top.scala 169:22]
  wire [7:0] n151_O_3; // @[Top.scala 169:22]
  wire [7:0] n151_O_4; // @[Top.scala 169:22]
  wire [7:0] n151_O_5; // @[Top.scala 169:22]
  wire [7:0] n151_O_6; // @[Top.scala 169:22]
  wire [7:0] n151_O_7; // @[Top.scala 169:22]
  wire [7:0] n151_O_8; // @[Top.scala 169:22]
  wire [7:0] n151_O_9; // @[Top.scala 169:22]
  wire [7:0] n151_O_10; // @[Top.scala 169:22]
  wire [7:0] n151_O_11; // @[Top.scala 169:22]
  wire [7:0] n151_O_12; // @[Top.scala 169:22]
  wire [7:0] n151_O_13; // @[Top.scala 169:22]
  wire [7:0] n151_O_14; // @[Top.scala 169:22]
  wire [7:0] n151_O_15; // @[Top.scala 169:22]
  wire  n152_valid_up; // @[Top.scala 172:22]
  wire  n152_valid_down; // @[Top.scala 172:22]
  wire [7:0] n152_I0_0; // @[Top.scala 172:22]
  wire [7:0] n152_I0_1; // @[Top.scala 172:22]
  wire [7:0] n152_I0_2; // @[Top.scala 172:22]
  wire [7:0] n152_I0_3; // @[Top.scala 172:22]
  wire [7:0] n152_I0_4; // @[Top.scala 172:22]
  wire [7:0] n152_I0_5; // @[Top.scala 172:22]
  wire [7:0] n152_I0_6; // @[Top.scala 172:22]
  wire [7:0] n152_I0_7; // @[Top.scala 172:22]
  wire [7:0] n152_I0_8; // @[Top.scala 172:22]
  wire [7:0] n152_I0_9; // @[Top.scala 172:22]
  wire [7:0] n152_I0_10; // @[Top.scala 172:22]
  wire [7:0] n152_I0_11; // @[Top.scala 172:22]
  wire [7:0] n152_I0_12; // @[Top.scala 172:22]
  wire [7:0] n152_I0_13; // @[Top.scala 172:22]
  wire [7:0] n152_I0_14; // @[Top.scala 172:22]
  wire [7:0] n152_I0_15; // @[Top.scala 172:22]
  wire [7:0] n152_I1_0; // @[Top.scala 172:22]
  wire [7:0] n152_I1_1; // @[Top.scala 172:22]
  wire [7:0] n152_I1_2; // @[Top.scala 172:22]
  wire [7:0] n152_I1_3; // @[Top.scala 172:22]
  wire [7:0] n152_I1_4; // @[Top.scala 172:22]
  wire [7:0] n152_I1_5; // @[Top.scala 172:22]
  wire [7:0] n152_I1_6; // @[Top.scala 172:22]
  wire [7:0] n152_I1_7; // @[Top.scala 172:22]
  wire [7:0] n152_I1_8; // @[Top.scala 172:22]
  wire [7:0] n152_I1_9; // @[Top.scala 172:22]
  wire [7:0] n152_I1_10; // @[Top.scala 172:22]
  wire [7:0] n152_I1_11; // @[Top.scala 172:22]
  wire [7:0] n152_I1_12; // @[Top.scala 172:22]
  wire [7:0] n152_I1_13; // @[Top.scala 172:22]
  wire [7:0] n152_I1_14; // @[Top.scala 172:22]
  wire [7:0] n152_I1_15; // @[Top.scala 172:22]
  wire [7:0] n152_O_0_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_0_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_1_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_1_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_2_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_2_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_3_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_3_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_4_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_4_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_5_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_5_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_6_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_6_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_7_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_7_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_8_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_8_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_9_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_9_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_10_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_10_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_11_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_11_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_12_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_12_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_13_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_13_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_14_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_14_1; // @[Top.scala 172:22]
  wire [7:0] n152_O_15_0; // @[Top.scala 172:22]
  wire [7:0] n152_O_15_1; // @[Top.scala 172:22]
  wire  n161_valid_up; // @[Top.scala 176:22]
  wire  n161_valid_down; // @[Top.scala 176:22]
  wire [7:0] n161_I_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_1_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_1_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_2_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_2_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_3_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_3_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_4_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_4_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_5_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_5_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_6_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_6_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_7_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_7_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_8_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_8_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_9_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_9_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_10_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_10_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_11_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_11_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_12_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_12_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_13_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_13_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_14_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_14_1; // @[Top.scala 176:22]
  wire [7:0] n161_I_15_0; // @[Top.scala 176:22]
  wire [7:0] n161_I_15_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_0_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_0_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_1_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_1_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_2_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_2_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_3_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_3_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_4_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_4_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_5_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_5_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_6_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_6_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_7_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_7_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_8_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_8_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_9_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_9_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_10_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_10_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_11_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_11_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_12_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_12_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_13_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_13_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_14_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_14_0_1; // @[Top.scala 176:22]
  wire [7:0] n161_O_15_0_0; // @[Top.scala 176:22]
  wire [7:0] n161_O_15_0_1; // @[Top.scala 176:22]
  wire  n168_valid_up; // @[Top.scala 179:22]
  wire  n168_valid_down; // @[Top.scala 179:22]
  wire [7:0] n168_I_0_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_0_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_1_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_1_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_2_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_2_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_3_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_3_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_4_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_4_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_5_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_5_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_6_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_6_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_7_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_7_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_8_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_8_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_9_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_9_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_10_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_10_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_11_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_11_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_12_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_12_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_13_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_13_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_14_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_14_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_I_15_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_I_15_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_0_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_0_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_1_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_1_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_2_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_2_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_3_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_3_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_4_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_4_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_5_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_5_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_6_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_6_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_7_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_7_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_8_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_8_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_9_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_9_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_10_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_10_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_11_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_11_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_12_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_12_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_13_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_13_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_14_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_14_1; // @[Top.scala 179:22]
  wire [7:0] n168_O_15_0; // @[Top.scala 179:22]
  wire [7:0] n168_O_15_1; // @[Top.scala 179:22]
  wire  n169_clock; // @[Top.scala 182:22]
  wire  n169_valid_up; // @[Top.scala 182:22]
  wire  n169_valid_down; // @[Top.scala 182:22]
  wire [7:0] n169_I_0; // @[Top.scala 182:22]
  wire [7:0] n169_I_1; // @[Top.scala 182:22]
  wire [7:0] n169_I_2; // @[Top.scala 182:22]
  wire [7:0] n169_I_3; // @[Top.scala 182:22]
  wire [7:0] n169_I_4; // @[Top.scala 182:22]
  wire [7:0] n169_I_5; // @[Top.scala 182:22]
  wire [7:0] n169_I_6; // @[Top.scala 182:22]
  wire [7:0] n169_I_7; // @[Top.scala 182:22]
  wire [7:0] n169_I_8; // @[Top.scala 182:22]
  wire [7:0] n169_I_9; // @[Top.scala 182:22]
  wire [7:0] n169_I_10; // @[Top.scala 182:22]
  wire [7:0] n169_I_11; // @[Top.scala 182:22]
  wire [7:0] n169_I_12; // @[Top.scala 182:22]
  wire [7:0] n169_I_13; // @[Top.scala 182:22]
  wire [7:0] n169_I_14; // @[Top.scala 182:22]
  wire [7:0] n169_I_15; // @[Top.scala 182:22]
  wire [7:0] n169_O_0; // @[Top.scala 182:22]
  wire [7:0] n169_O_1; // @[Top.scala 182:22]
  wire [7:0] n169_O_2; // @[Top.scala 182:22]
  wire [7:0] n169_O_3; // @[Top.scala 182:22]
  wire [7:0] n169_O_4; // @[Top.scala 182:22]
  wire [7:0] n169_O_5; // @[Top.scala 182:22]
  wire [7:0] n169_O_6; // @[Top.scala 182:22]
  wire [7:0] n169_O_7; // @[Top.scala 182:22]
  wire [7:0] n169_O_8; // @[Top.scala 182:22]
  wire [7:0] n169_O_9; // @[Top.scala 182:22]
  wire [7:0] n169_O_10; // @[Top.scala 182:22]
  wire [7:0] n169_O_11; // @[Top.scala 182:22]
  wire [7:0] n169_O_12; // @[Top.scala 182:22]
  wire [7:0] n169_O_13; // @[Top.scala 182:22]
  wire [7:0] n169_O_14; // @[Top.scala 182:22]
  wire [7:0] n169_O_15; // @[Top.scala 182:22]
  wire  n170_valid_up; // @[Top.scala 185:22]
  wire  n170_valid_down; // @[Top.scala 185:22]
  wire [7:0] n170_I0_0; // @[Top.scala 185:22]
  wire [7:0] n170_I0_1; // @[Top.scala 185:22]
  wire [7:0] n170_I0_2; // @[Top.scala 185:22]
  wire [7:0] n170_I0_3; // @[Top.scala 185:22]
  wire [7:0] n170_I0_4; // @[Top.scala 185:22]
  wire [7:0] n170_I0_5; // @[Top.scala 185:22]
  wire [7:0] n170_I0_6; // @[Top.scala 185:22]
  wire [7:0] n170_I0_7; // @[Top.scala 185:22]
  wire [7:0] n170_I0_8; // @[Top.scala 185:22]
  wire [7:0] n170_I0_9; // @[Top.scala 185:22]
  wire [7:0] n170_I0_10; // @[Top.scala 185:22]
  wire [7:0] n170_I0_11; // @[Top.scala 185:22]
  wire [7:0] n170_I0_12; // @[Top.scala 185:22]
  wire [7:0] n170_I0_13; // @[Top.scala 185:22]
  wire [7:0] n170_I0_14; // @[Top.scala 185:22]
  wire [7:0] n170_I0_15; // @[Top.scala 185:22]
  wire [7:0] n170_I1_0; // @[Top.scala 185:22]
  wire [7:0] n170_I1_1; // @[Top.scala 185:22]
  wire [7:0] n170_I1_2; // @[Top.scala 185:22]
  wire [7:0] n170_I1_3; // @[Top.scala 185:22]
  wire [7:0] n170_I1_4; // @[Top.scala 185:22]
  wire [7:0] n170_I1_5; // @[Top.scala 185:22]
  wire [7:0] n170_I1_6; // @[Top.scala 185:22]
  wire [7:0] n170_I1_7; // @[Top.scala 185:22]
  wire [7:0] n170_I1_8; // @[Top.scala 185:22]
  wire [7:0] n170_I1_9; // @[Top.scala 185:22]
  wire [7:0] n170_I1_10; // @[Top.scala 185:22]
  wire [7:0] n170_I1_11; // @[Top.scala 185:22]
  wire [7:0] n170_I1_12; // @[Top.scala 185:22]
  wire [7:0] n170_I1_13; // @[Top.scala 185:22]
  wire [7:0] n170_I1_14; // @[Top.scala 185:22]
  wire [7:0] n170_I1_15; // @[Top.scala 185:22]
  wire [7:0] n170_O_0_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_0_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_1_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_1_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_2_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_2_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_3_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_3_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_4_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_4_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_5_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_5_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_6_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_6_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_7_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_7_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_8_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_8_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_9_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_9_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_10_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_10_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_11_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_11_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_12_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_12_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_13_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_13_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_14_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_14_1; // @[Top.scala 185:22]
  wire [7:0] n170_O_15_0; // @[Top.scala 185:22]
  wire [7:0] n170_O_15_1; // @[Top.scala 185:22]
  wire  n179_valid_up; // @[Top.scala 189:22]
  wire  n179_valid_down; // @[Top.scala 189:22]
  wire [7:0] n179_I_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_1_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_1_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_2_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_2_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_3_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_3_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_4_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_4_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_5_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_5_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_6_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_6_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_7_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_7_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_8_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_8_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_9_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_9_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_10_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_10_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_11_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_11_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_12_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_12_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_13_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_13_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_14_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_14_1; // @[Top.scala 189:22]
  wire [7:0] n179_I_15_0; // @[Top.scala 189:22]
  wire [7:0] n179_I_15_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_0_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_0_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_1_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_1_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_2_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_2_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_3_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_3_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_4_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_4_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_5_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_5_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_6_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_6_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_7_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_7_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_8_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_8_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_9_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_9_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_10_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_10_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_11_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_11_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_12_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_12_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_13_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_13_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_14_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_14_0_1; // @[Top.scala 189:22]
  wire [7:0] n179_O_15_0_0; // @[Top.scala 189:22]
  wire [7:0] n179_O_15_0_1; // @[Top.scala 189:22]
  wire  n186_valid_up; // @[Top.scala 192:22]
  wire  n186_valid_down; // @[Top.scala 192:22]
  wire [7:0] n186_I_0_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_0_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_1_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_1_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_2_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_2_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_3_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_3_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_4_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_4_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_5_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_5_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_6_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_6_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_7_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_7_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_8_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_8_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_9_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_9_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_10_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_10_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_11_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_11_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_12_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_12_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_13_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_13_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_14_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_14_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_I_15_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_I_15_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_0_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_0_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_1_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_1_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_2_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_2_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_3_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_3_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_4_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_4_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_5_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_5_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_6_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_6_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_7_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_7_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_8_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_8_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_9_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_9_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_10_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_10_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_11_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_11_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_12_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_12_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_13_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_13_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_14_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_14_1; // @[Top.scala 192:22]
  wire [7:0] n186_O_15_0; // @[Top.scala 192:22]
  wire [7:0] n186_O_15_1; // @[Top.scala 192:22]
  wire  n187_valid_up; // @[Top.scala 195:22]
  wire  n187_valid_down; // @[Top.scala 195:22]
  wire [7:0] n187_I0_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_2_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_2_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_3_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_3_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_4_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_4_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_5_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_5_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_6_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_6_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_7_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_7_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_8_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_8_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_9_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_9_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_10_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_10_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_11_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_11_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_12_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_12_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_13_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_13_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_14_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_14_1; // @[Top.scala 195:22]
  wire [7:0] n187_I0_15_0; // @[Top.scala 195:22]
  wire [7:0] n187_I0_15_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_2_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_2_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_3_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_3_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_4_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_4_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_5_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_5_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_6_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_6_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_7_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_7_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_8_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_8_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_9_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_9_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_10_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_10_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_11_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_11_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_12_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_12_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_13_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_13_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_14_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_14_1; // @[Top.scala 195:22]
  wire [7:0] n187_I1_15_0; // @[Top.scala 195:22]
  wire [7:0] n187_I1_15_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_0_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_0_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_0_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_0_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_1_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_1_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_1_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_1_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_2_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_2_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_2_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_2_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_3_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_3_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_3_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_3_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_4_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_4_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_4_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_4_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_5_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_5_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_5_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_5_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_6_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_6_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_6_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_6_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_7_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_7_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_7_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_7_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_8_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_8_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_8_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_8_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_9_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_9_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_9_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_9_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_10_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_10_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_10_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_10_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_11_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_11_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_11_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_11_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_12_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_12_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_12_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_12_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_13_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_13_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_13_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_13_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_14_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_14_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_14_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_14_1_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_15_0_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_15_0_1; // @[Top.scala 195:22]
  wire [7:0] n187_O_15_1_0; // @[Top.scala 195:22]
  wire [7:0] n187_O_15_1_1; // @[Top.scala 195:22]
  wire  n196_valid_up; // @[Top.scala 199:22]
  wire  n196_valid_down; // @[Top.scala 199:22]
  wire [7:0] n196_I_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_1_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_1_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_1_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_1_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_2_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_2_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_2_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_2_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_3_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_3_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_3_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_3_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_4_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_4_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_4_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_4_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_5_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_5_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_5_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_5_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_6_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_6_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_6_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_6_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_7_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_7_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_7_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_7_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_8_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_8_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_8_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_8_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_9_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_9_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_9_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_9_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_10_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_10_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_10_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_10_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_11_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_11_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_11_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_11_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_12_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_12_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_12_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_12_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_13_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_13_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_13_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_13_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_14_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_14_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_14_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_14_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_15_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_15_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_I_15_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_I_15_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_0_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_0_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_0_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_0_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_1_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_1_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_1_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_1_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_2_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_2_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_2_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_2_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_3_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_3_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_3_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_3_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_4_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_4_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_4_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_4_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_5_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_5_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_5_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_5_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_6_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_6_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_6_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_6_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_7_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_7_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_7_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_7_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_8_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_8_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_8_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_8_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_9_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_9_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_9_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_9_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_10_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_10_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_10_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_10_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_11_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_11_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_11_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_11_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_12_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_12_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_12_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_12_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_13_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_13_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_13_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_13_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_14_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_14_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_14_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_14_0_1_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_15_0_0_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_15_0_0_1; // @[Top.scala 199:22]
  wire [7:0] n196_O_15_0_1_0; // @[Top.scala 199:22]
  wire [7:0] n196_O_15_0_1_1; // @[Top.scala 199:22]
  wire  n203_valid_up; // @[Top.scala 202:22]
  wire  n203_valid_down; // @[Top.scala 202:22]
  wire [7:0] n203_I_0_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_0_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_0_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_0_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_1_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_1_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_1_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_1_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_2_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_2_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_2_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_2_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_3_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_3_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_3_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_3_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_4_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_4_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_4_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_4_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_5_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_5_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_5_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_5_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_6_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_6_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_6_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_6_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_7_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_7_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_7_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_7_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_8_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_8_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_8_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_8_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_9_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_9_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_9_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_9_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_10_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_10_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_10_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_10_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_11_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_11_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_11_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_11_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_12_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_12_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_12_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_12_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_13_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_13_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_13_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_13_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_14_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_14_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_14_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_14_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_15_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_15_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_I_15_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_I_15_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_0_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_0_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_0_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_0_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_1_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_1_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_1_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_1_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_2_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_2_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_2_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_2_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_3_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_3_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_3_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_3_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_4_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_4_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_4_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_4_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_5_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_5_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_5_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_5_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_6_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_6_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_6_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_6_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_7_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_7_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_7_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_7_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_8_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_8_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_8_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_8_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_9_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_9_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_9_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_9_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_10_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_10_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_10_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_10_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_11_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_11_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_11_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_11_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_12_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_12_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_12_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_12_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_13_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_13_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_13_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_13_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_14_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_14_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_14_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_14_1_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_15_0_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_15_0_1; // @[Top.scala 202:22]
  wire [7:0] n203_O_15_1_0; // @[Top.scala 202:22]
  wire [7:0] n203_O_15_1_1; // @[Top.scala 202:22]
  wire  n245_clock; // @[Top.scala 205:22]
  wire  n245_reset; // @[Top.scala 205:22]
  wire  n245_valid_up; // @[Top.scala 205:22]
  wire  n245_valid_down; // @[Top.scala 205:22]
  wire [7:0] n245_I_0_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_0_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_0_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_0_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_1_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_1_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_1_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_1_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_2_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_2_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_2_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_2_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_3_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_3_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_3_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_3_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_4_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_4_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_4_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_4_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_5_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_5_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_5_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_5_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_6_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_6_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_6_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_6_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_7_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_7_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_7_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_7_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_8_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_8_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_8_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_8_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_9_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_9_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_9_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_9_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_10_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_10_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_10_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_10_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_11_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_11_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_11_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_11_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_12_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_12_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_12_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_12_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_13_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_13_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_13_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_13_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_14_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_14_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_14_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_14_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_15_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_15_0_1; // @[Top.scala 205:22]
  wire [7:0] n245_I_15_1_0; // @[Top.scala 205:22]
  wire [7:0] n245_I_15_1_1; // @[Top.scala 205:22]
  wire [7:0] n245_O_0_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_1_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_2_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_3_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_4_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_5_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_6_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_7_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_8_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_9_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_10_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_11_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_12_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_13_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_14_0_0; // @[Top.scala 205:22]
  wire [7:0] n245_O_15_0_0; // @[Top.scala 205:22]
  wire  n246_valid_up; // @[Top.scala 208:22]
  wire  n246_valid_down; // @[Top.scala 208:22]
  wire [7:0] n246_I_0_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_1_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_2_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_3_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_4_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_5_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_6_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_7_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_8_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_9_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_10_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_11_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_12_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_13_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_14_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_I_15_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_0_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_1_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_2_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_3_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_4_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_5_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_6_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_7_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_8_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_9_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_10_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_11_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_12_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_13_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_14_0; // @[Top.scala 208:22]
  wire [7:0] n246_O_15_0; // @[Top.scala 208:22]
  wire  n247_valid_up; // @[Top.scala 211:22]
  wire  n247_valid_down; // @[Top.scala 211:22]
  wire [7:0] n247_I_0_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_1_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_2_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_3_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_4_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_5_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_6_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_7_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_8_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_9_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_10_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_11_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_12_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_13_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_14_0; // @[Top.scala 211:22]
  wire [7:0] n247_I_15_0; // @[Top.scala 211:22]
  wire [7:0] n247_O_0; // @[Top.scala 211:22]
  wire [7:0] n247_O_1; // @[Top.scala 211:22]
  wire [7:0] n247_O_2; // @[Top.scala 211:22]
  wire [7:0] n247_O_3; // @[Top.scala 211:22]
  wire [7:0] n247_O_4; // @[Top.scala 211:22]
  wire [7:0] n247_O_5; // @[Top.scala 211:22]
  wire [7:0] n247_O_6; // @[Top.scala 211:22]
  wire [7:0] n247_O_7; // @[Top.scala 211:22]
  wire [7:0] n247_O_8; // @[Top.scala 211:22]
  wire [7:0] n247_O_9; // @[Top.scala 211:22]
  wire [7:0] n247_O_10; // @[Top.scala 211:22]
  wire [7:0] n247_O_11; // @[Top.scala 211:22]
  wire [7:0] n247_O_12; // @[Top.scala 211:22]
  wire [7:0] n247_O_13; // @[Top.scala 211:22]
  wire [7:0] n247_O_14; // @[Top.scala 211:22]
  wire [7:0] n247_O_15; // @[Top.scala 211:22]
  wire  n248_clock; // @[Top.scala 214:22]
  wire  n248_reset; // @[Top.scala 214:22]
  wire  n248_valid_up; // @[Top.scala 214:22]
  wire  n248_valid_down; // @[Top.scala 214:22]
  wire [7:0] n248_I_0; // @[Top.scala 214:22]
  wire [7:0] n248_I_1; // @[Top.scala 214:22]
  wire [7:0] n248_I_2; // @[Top.scala 214:22]
  wire [7:0] n248_I_3; // @[Top.scala 214:22]
  wire [7:0] n248_I_4; // @[Top.scala 214:22]
  wire [7:0] n248_I_5; // @[Top.scala 214:22]
  wire [7:0] n248_I_6; // @[Top.scala 214:22]
  wire [7:0] n248_I_7; // @[Top.scala 214:22]
  wire [7:0] n248_I_8; // @[Top.scala 214:22]
  wire [7:0] n248_I_9; // @[Top.scala 214:22]
  wire [7:0] n248_I_10; // @[Top.scala 214:22]
  wire [7:0] n248_I_11; // @[Top.scala 214:22]
  wire [7:0] n248_I_12; // @[Top.scala 214:22]
  wire [7:0] n248_I_13; // @[Top.scala 214:22]
  wire [7:0] n248_I_14; // @[Top.scala 214:22]
  wire [7:0] n248_I_15; // @[Top.scala 214:22]
  wire [7:0] n248_O_0; // @[Top.scala 214:22]
  wire [7:0] n248_O_1; // @[Top.scala 214:22]
  wire [7:0] n248_O_2; // @[Top.scala 214:22]
  wire [7:0] n248_O_3; // @[Top.scala 214:22]
  wire [7:0] n248_O_4; // @[Top.scala 214:22]
  wire [7:0] n248_O_5; // @[Top.scala 214:22]
  wire [7:0] n248_O_6; // @[Top.scala 214:22]
  wire [7:0] n248_O_7; // @[Top.scala 214:22]
  wire [7:0] n248_O_8; // @[Top.scala 214:22]
  wire [7:0] n248_O_9; // @[Top.scala 214:22]
  wire [7:0] n248_O_10; // @[Top.scala 214:22]
  wire [7:0] n248_O_11; // @[Top.scala 214:22]
  wire [7:0] n248_O_12; // @[Top.scala 214:22]
  wire [7:0] n248_O_13; // @[Top.scala 214:22]
  wire [7:0] n248_O_14; // @[Top.scala 214:22]
  wire [7:0] n248_O_15; // @[Top.scala 214:22]
  wire  n249_clock; // @[Top.scala 217:22]
  wire  n249_reset; // @[Top.scala 217:22]
  wire  n249_valid_up; // @[Top.scala 217:22]
  wire  n249_valid_down; // @[Top.scala 217:22]
  wire [7:0] n249_I_0; // @[Top.scala 217:22]
  wire [7:0] n249_I_1; // @[Top.scala 217:22]
  wire [7:0] n249_I_2; // @[Top.scala 217:22]
  wire [7:0] n249_I_3; // @[Top.scala 217:22]
  wire [7:0] n249_I_4; // @[Top.scala 217:22]
  wire [7:0] n249_I_5; // @[Top.scala 217:22]
  wire [7:0] n249_I_6; // @[Top.scala 217:22]
  wire [7:0] n249_I_7; // @[Top.scala 217:22]
  wire [7:0] n249_I_8; // @[Top.scala 217:22]
  wire [7:0] n249_I_9; // @[Top.scala 217:22]
  wire [7:0] n249_I_10; // @[Top.scala 217:22]
  wire [7:0] n249_I_11; // @[Top.scala 217:22]
  wire [7:0] n249_I_12; // @[Top.scala 217:22]
  wire [7:0] n249_I_13; // @[Top.scala 217:22]
  wire [7:0] n249_I_14; // @[Top.scala 217:22]
  wire [7:0] n249_I_15; // @[Top.scala 217:22]
  wire [7:0] n249_O_0; // @[Top.scala 217:22]
  wire [7:0] n249_O_1; // @[Top.scala 217:22]
  wire [7:0] n249_O_2; // @[Top.scala 217:22]
  wire [7:0] n249_O_3; // @[Top.scala 217:22]
  wire [7:0] n249_O_4; // @[Top.scala 217:22]
  wire [7:0] n249_O_5; // @[Top.scala 217:22]
  wire [7:0] n249_O_6; // @[Top.scala 217:22]
  wire [7:0] n249_O_7; // @[Top.scala 217:22]
  wire [7:0] n249_O_8; // @[Top.scala 217:22]
  wire [7:0] n249_O_9; // @[Top.scala 217:22]
  wire [7:0] n249_O_10; // @[Top.scala 217:22]
  wire [7:0] n249_O_11; // @[Top.scala 217:22]
  wire [7:0] n249_O_12; // @[Top.scala 217:22]
  wire [7:0] n249_O_13; // @[Top.scala 217:22]
  wire [7:0] n249_O_14; // @[Top.scala 217:22]
  wire [7:0] n249_O_15; // @[Top.scala 217:22]
  wire  n250_clock; // @[Top.scala 220:22]
  wire  n250_reset; // @[Top.scala 220:22]
  wire  n250_valid_up; // @[Top.scala 220:22]
  wire  n250_valid_down; // @[Top.scala 220:22]
  wire [7:0] n250_I_0; // @[Top.scala 220:22]
  wire [7:0] n250_I_1; // @[Top.scala 220:22]
  wire [7:0] n250_I_2; // @[Top.scala 220:22]
  wire [7:0] n250_I_3; // @[Top.scala 220:22]
  wire [7:0] n250_I_4; // @[Top.scala 220:22]
  wire [7:0] n250_I_5; // @[Top.scala 220:22]
  wire [7:0] n250_I_6; // @[Top.scala 220:22]
  wire [7:0] n250_I_7; // @[Top.scala 220:22]
  wire [7:0] n250_I_8; // @[Top.scala 220:22]
  wire [7:0] n250_I_9; // @[Top.scala 220:22]
  wire [7:0] n250_I_10; // @[Top.scala 220:22]
  wire [7:0] n250_I_11; // @[Top.scala 220:22]
  wire [7:0] n250_I_12; // @[Top.scala 220:22]
  wire [7:0] n250_I_13; // @[Top.scala 220:22]
  wire [7:0] n250_I_14; // @[Top.scala 220:22]
  wire [7:0] n250_I_15; // @[Top.scala 220:22]
  wire [7:0] n250_O_0; // @[Top.scala 220:22]
  wire [7:0] n250_O_1; // @[Top.scala 220:22]
  wire [7:0] n250_O_2; // @[Top.scala 220:22]
  wire [7:0] n250_O_3; // @[Top.scala 220:22]
  wire [7:0] n250_O_4; // @[Top.scala 220:22]
  wire [7:0] n250_O_5; // @[Top.scala 220:22]
  wire [7:0] n250_O_6; // @[Top.scala 220:22]
  wire [7:0] n250_O_7; // @[Top.scala 220:22]
  wire [7:0] n250_O_8; // @[Top.scala 220:22]
  wire [7:0] n250_O_9; // @[Top.scala 220:22]
  wire [7:0] n250_O_10; // @[Top.scala 220:22]
  wire [7:0] n250_O_11; // @[Top.scala 220:22]
  wire [7:0] n250_O_12; // @[Top.scala 220:22]
  wire [7:0] n250_O_13; // @[Top.scala 220:22]
  wire [7:0] n250_O_14; // @[Top.scala 220:22]
  wire [7:0] n250_O_15; // @[Top.scala 220:22]
  FIFO n1 ( // @[Top.scala 74:20]
    .clock(n1_clock),
    .reset(n1_reset),
    .valid_up(n1_valid_up),
    .valid_down(n1_valid_down),
    .I_0(n1_I_0),
    .I_1(n1_I_1),
    .I_2(n1_I_2),
    .I_3(n1_I_3),
    .I_4(n1_I_4),
    .I_5(n1_I_5),
    .I_6(n1_I_6),
    .I_7(n1_I_7),
    .I_8(n1_I_8),
    .I_9(n1_I_9),
    .I_10(n1_I_10),
    .I_11(n1_I_11),
    .I_12(n1_I_12),
    .I_13(n1_I_13),
    .I_14(n1_I_14),
    .I_15(n1_I_15),
    .O_0(n1_O_0),
    .O_1(n1_O_1),
    .O_2(n1_O_2),
    .O_3(n1_O_3),
    .O_4(n1_O_4),
    .O_5(n1_O_5),
    .O_6(n1_O_6),
    .O_7(n1_O_7),
    .O_8(n1_O_8),
    .O_9(n1_O_9),
    .O_10(n1_O_10),
    .O_11(n1_O_11),
    .O_12(n1_O_12),
    .O_13(n1_O_13),
    .O_14(n1_O_14),
    .O_15(n1_O_15)
  );
  ShiftTS n2 ( // @[Top.scala 77:20]
    .clock(n2_clock),
    .reset(n2_reset),
    .valid_up(n2_valid_up),
    .valid_down(n2_valid_down),
    .I_0(n2_I_0),
    .I_1(n2_I_1),
    .I_2(n2_I_2),
    .I_3(n2_I_3),
    .I_4(n2_I_4),
    .I_5(n2_I_5),
    .I_6(n2_I_6),
    .I_7(n2_I_7),
    .I_8(n2_I_8),
    .I_9(n2_I_9),
    .I_10(n2_I_10),
    .I_11(n2_I_11),
    .I_12(n2_I_12),
    .I_13(n2_I_13),
    .I_14(n2_I_14),
    .I_15(n2_I_15),
    .O_0(n2_O_0),
    .O_1(n2_O_1),
    .O_2(n2_O_2),
    .O_3(n2_O_3),
    .O_4(n2_O_4),
    .O_5(n2_O_5),
    .O_6(n2_O_6),
    .O_7(n2_O_7),
    .O_8(n2_O_8),
    .O_9(n2_O_9),
    .O_10(n2_O_10),
    .O_11(n2_O_11),
    .O_12(n2_O_12),
    .O_13(n2_O_13),
    .O_14(n2_O_14),
    .O_15(n2_O_15)
  );
  ShiftTS n3 ( // @[Top.scala 80:20]
    .clock(n3_clock),
    .reset(n3_reset),
    .valid_up(n3_valid_up),
    .valid_down(n3_valid_down),
    .I_0(n3_I_0),
    .I_1(n3_I_1),
    .I_2(n3_I_2),
    .I_3(n3_I_3),
    .I_4(n3_I_4),
    .I_5(n3_I_5),
    .I_6(n3_I_6),
    .I_7(n3_I_7),
    .I_8(n3_I_8),
    .I_9(n3_I_9),
    .I_10(n3_I_10),
    .I_11(n3_I_11),
    .I_12(n3_I_12),
    .I_13(n3_I_13),
    .I_14(n3_I_14),
    .I_15(n3_I_15),
    .O_0(n3_O_0),
    .O_1(n3_O_1),
    .O_2(n3_O_2),
    .O_3(n3_O_3),
    .O_4(n3_O_4),
    .O_5(n3_O_5),
    .O_6(n3_O_6),
    .O_7(n3_O_7),
    .O_8(n3_O_8),
    .O_9(n3_O_9),
    .O_10(n3_O_10),
    .O_11(n3_O_11),
    .O_12(n3_O_12),
    .O_13(n3_O_13),
    .O_14(n3_O_14),
    .O_15(n3_O_15)
  );
  ShiftTS_2 n4 ( // @[Top.scala 83:20]
    .clock(n4_clock),
    .valid_up(n4_valid_up),
    .valid_down(n4_valid_down),
    .I_0(n4_I_0),
    .I_1(n4_I_1),
    .I_2(n4_I_2),
    .I_3(n4_I_3),
    .I_4(n4_I_4),
    .I_5(n4_I_5),
    .I_6(n4_I_6),
    .I_7(n4_I_7),
    .I_8(n4_I_8),
    .I_9(n4_I_9),
    .I_10(n4_I_10),
    .I_11(n4_I_11),
    .I_12(n4_I_12),
    .I_13(n4_I_13),
    .I_14(n4_I_14),
    .I_15(n4_I_15),
    .O_0(n4_O_0),
    .O_1(n4_O_1),
    .O_2(n4_O_2),
    .O_3(n4_O_3),
    .O_4(n4_O_4),
    .O_5(n4_O_5),
    .O_6(n4_O_6),
    .O_7(n4_O_7),
    .O_8(n4_O_8),
    .O_9(n4_O_9),
    .O_10(n4_O_10),
    .O_11(n4_O_11),
    .O_12(n4_O_12),
    .O_13(n4_O_13),
    .O_14(n4_O_14),
    .O_15(n4_O_15)
  );
  ShiftTS_2 n5 ( // @[Top.scala 86:20]
    .clock(n5_clock),
    .valid_up(n5_valid_up),
    .valid_down(n5_valid_down),
    .I_0(n5_I_0),
    .I_1(n5_I_1),
    .I_2(n5_I_2),
    .I_3(n5_I_3),
    .I_4(n5_I_4),
    .I_5(n5_I_5),
    .I_6(n5_I_6),
    .I_7(n5_I_7),
    .I_8(n5_I_8),
    .I_9(n5_I_9),
    .I_10(n5_I_10),
    .I_11(n5_I_11),
    .I_12(n5_I_12),
    .I_13(n5_I_13),
    .I_14(n5_I_14),
    .I_15(n5_I_15),
    .O_0(n5_O_0),
    .O_1(n5_O_1),
    .O_2(n5_O_2),
    .O_3(n5_O_3),
    .O_4(n5_O_4),
    .O_5(n5_O_5),
    .O_6(n5_O_6),
    .O_7(n5_O_7),
    .O_8(n5_O_8),
    .O_9(n5_O_9),
    .O_10(n5_O_10),
    .O_11(n5_O_11),
    .O_12(n5_O_12),
    .O_13(n5_O_13),
    .O_14(n5_O_14),
    .O_15(n5_O_15)
  );
  Map2T n6 ( // @[Top.scala 89:20]
    .valid_up(n6_valid_up),
    .valid_down(n6_valid_down),
    .I0_0(n6_I0_0),
    .I0_1(n6_I0_1),
    .I0_2(n6_I0_2),
    .I0_3(n6_I0_3),
    .I0_4(n6_I0_4),
    .I0_5(n6_I0_5),
    .I0_6(n6_I0_6),
    .I0_7(n6_I0_7),
    .I0_8(n6_I0_8),
    .I0_9(n6_I0_9),
    .I0_10(n6_I0_10),
    .I0_11(n6_I0_11),
    .I0_12(n6_I0_12),
    .I0_13(n6_I0_13),
    .I0_14(n6_I0_14),
    .I0_15(n6_I0_15),
    .I1_0(n6_I1_0),
    .I1_1(n6_I1_1),
    .I1_2(n6_I1_2),
    .I1_3(n6_I1_3),
    .I1_4(n6_I1_4),
    .I1_5(n6_I1_5),
    .I1_6(n6_I1_6),
    .I1_7(n6_I1_7),
    .I1_8(n6_I1_8),
    .I1_9(n6_I1_9),
    .I1_10(n6_I1_10),
    .I1_11(n6_I1_11),
    .I1_12(n6_I1_12),
    .I1_13(n6_I1_13),
    .I1_14(n6_I1_14),
    .I1_15(n6_I1_15),
    .O_0_0(n6_O_0_0),
    .O_0_1(n6_O_0_1),
    .O_1_0(n6_O_1_0),
    .O_1_1(n6_O_1_1),
    .O_2_0(n6_O_2_0),
    .O_2_1(n6_O_2_1),
    .O_3_0(n6_O_3_0),
    .O_3_1(n6_O_3_1),
    .O_4_0(n6_O_4_0),
    .O_4_1(n6_O_4_1),
    .O_5_0(n6_O_5_0),
    .O_5_1(n6_O_5_1),
    .O_6_0(n6_O_6_0),
    .O_6_1(n6_O_6_1),
    .O_7_0(n6_O_7_0),
    .O_7_1(n6_O_7_1),
    .O_8_0(n6_O_8_0),
    .O_8_1(n6_O_8_1),
    .O_9_0(n6_O_9_0),
    .O_9_1(n6_O_9_1),
    .O_10_0(n6_O_10_0),
    .O_10_1(n6_O_10_1),
    .O_11_0(n6_O_11_0),
    .O_11_1(n6_O_11_1),
    .O_12_0(n6_O_12_0),
    .O_12_1(n6_O_12_1),
    .O_13_0(n6_O_13_0),
    .O_13_1(n6_O_13_1),
    .O_14_0(n6_O_14_0),
    .O_14_1(n6_O_14_1),
    .O_15_0(n6_O_15_0),
    .O_15_1(n6_O_15_1)
  );
  Map2T_1 n13 ( // @[Top.scala 93:21]
    .valid_up(n13_valid_up),
    .valid_down(n13_valid_down),
    .I0_0_0(n13_I0_0_0),
    .I0_0_1(n13_I0_0_1),
    .I0_1_0(n13_I0_1_0),
    .I0_1_1(n13_I0_1_1),
    .I0_2_0(n13_I0_2_0),
    .I0_2_1(n13_I0_2_1),
    .I0_3_0(n13_I0_3_0),
    .I0_3_1(n13_I0_3_1),
    .I0_4_0(n13_I0_4_0),
    .I0_4_1(n13_I0_4_1),
    .I0_5_0(n13_I0_5_0),
    .I0_5_1(n13_I0_5_1),
    .I0_6_0(n13_I0_6_0),
    .I0_6_1(n13_I0_6_1),
    .I0_7_0(n13_I0_7_0),
    .I0_7_1(n13_I0_7_1),
    .I0_8_0(n13_I0_8_0),
    .I0_8_1(n13_I0_8_1),
    .I0_9_0(n13_I0_9_0),
    .I0_9_1(n13_I0_9_1),
    .I0_10_0(n13_I0_10_0),
    .I0_10_1(n13_I0_10_1),
    .I0_11_0(n13_I0_11_0),
    .I0_11_1(n13_I0_11_1),
    .I0_12_0(n13_I0_12_0),
    .I0_12_1(n13_I0_12_1),
    .I0_13_0(n13_I0_13_0),
    .I0_13_1(n13_I0_13_1),
    .I0_14_0(n13_I0_14_0),
    .I0_14_1(n13_I0_14_1),
    .I0_15_0(n13_I0_15_0),
    .I0_15_1(n13_I0_15_1),
    .I1_0(n13_I1_0),
    .I1_1(n13_I1_1),
    .I1_2(n13_I1_2),
    .I1_3(n13_I1_3),
    .I1_4(n13_I1_4),
    .I1_5(n13_I1_5),
    .I1_6(n13_I1_6),
    .I1_7(n13_I1_7),
    .I1_8(n13_I1_8),
    .I1_9(n13_I1_9),
    .I1_10(n13_I1_10),
    .I1_11(n13_I1_11),
    .I1_12(n13_I1_12),
    .I1_13(n13_I1_13),
    .I1_14(n13_I1_14),
    .I1_15(n13_I1_15),
    .O_0_0(n13_O_0_0),
    .O_0_1(n13_O_0_1),
    .O_0_2(n13_O_0_2),
    .O_1_0(n13_O_1_0),
    .O_1_1(n13_O_1_1),
    .O_1_2(n13_O_1_2),
    .O_2_0(n13_O_2_0),
    .O_2_1(n13_O_2_1),
    .O_2_2(n13_O_2_2),
    .O_3_0(n13_O_3_0),
    .O_3_1(n13_O_3_1),
    .O_3_2(n13_O_3_2),
    .O_4_0(n13_O_4_0),
    .O_4_1(n13_O_4_1),
    .O_4_2(n13_O_4_2),
    .O_5_0(n13_O_5_0),
    .O_5_1(n13_O_5_1),
    .O_5_2(n13_O_5_2),
    .O_6_0(n13_O_6_0),
    .O_6_1(n13_O_6_1),
    .O_6_2(n13_O_6_2),
    .O_7_0(n13_O_7_0),
    .O_7_1(n13_O_7_1),
    .O_7_2(n13_O_7_2),
    .O_8_0(n13_O_8_0),
    .O_8_1(n13_O_8_1),
    .O_8_2(n13_O_8_2),
    .O_9_0(n13_O_9_0),
    .O_9_1(n13_O_9_1),
    .O_9_2(n13_O_9_2),
    .O_10_0(n13_O_10_0),
    .O_10_1(n13_O_10_1),
    .O_10_2(n13_O_10_2),
    .O_11_0(n13_O_11_0),
    .O_11_1(n13_O_11_1),
    .O_11_2(n13_O_11_2),
    .O_12_0(n13_O_12_0),
    .O_12_1(n13_O_12_1),
    .O_12_2(n13_O_12_2),
    .O_13_0(n13_O_13_0),
    .O_13_1(n13_O_13_1),
    .O_13_2(n13_O_13_2),
    .O_14_0(n13_O_14_0),
    .O_14_1(n13_O_14_1),
    .O_14_2(n13_O_14_2),
    .O_15_0(n13_O_15_0),
    .O_15_1(n13_O_15_1),
    .O_15_2(n13_O_15_2)
  );
  MapT n22 ( // @[Top.scala 97:21]
    .valid_up(n22_valid_up),
    .valid_down(n22_valid_down),
    .I_0_0(n22_I_0_0),
    .I_0_1(n22_I_0_1),
    .I_0_2(n22_I_0_2),
    .I_1_0(n22_I_1_0),
    .I_1_1(n22_I_1_1),
    .I_1_2(n22_I_1_2),
    .I_2_0(n22_I_2_0),
    .I_2_1(n22_I_2_1),
    .I_2_2(n22_I_2_2),
    .I_3_0(n22_I_3_0),
    .I_3_1(n22_I_3_1),
    .I_3_2(n22_I_3_2),
    .I_4_0(n22_I_4_0),
    .I_4_1(n22_I_4_1),
    .I_4_2(n22_I_4_2),
    .I_5_0(n22_I_5_0),
    .I_5_1(n22_I_5_1),
    .I_5_2(n22_I_5_2),
    .I_6_0(n22_I_6_0),
    .I_6_1(n22_I_6_1),
    .I_6_2(n22_I_6_2),
    .I_7_0(n22_I_7_0),
    .I_7_1(n22_I_7_1),
    .I_7_2(n22_I_7_2),
    .I_8_0(n22_I_8_0),
    .I_8_1(n22_I_8_1),
    .I_8_2(n22_I_8_2),
    .I_9_0(n22_I_9_0),
    .I_9_1(n22_I_9_1),
    .I_9_2(n22_I_9_2),
    .I_10_0(n22_I_10_0),
    .I_10_1(n22_I_10_1),
    .I_10_2(n22_I_10_2),
    .I_11_0(n22_I_11_0),
    .I_11_1(n22_I_11_1),
    .I_11_2(n22_I_11_2),
    .I_12_0(n22_I_12_0),
    .I_12_1(n22_I_12_1),
    .I_12_2(n22_I_12_2),
    .I_13_0(n22_I_13_0),
    .I_13_1(n22_I_13_1),
    .I_13_2(n22_I_13_2),
    .I_14_0(n22_I_14_0),
    .I_14_1(n22_I_14_1),
    .I_14_2(n22_I_14_2),
    .I_15_0(n22_I_15_0),
    .I_15_1(n22_I_15_1),
    .I_15_2(n22_I_15_2),
    .O_0_0_0(n22_O_0_0_0),
    .O_0_0_1(n22_O_0_0_1),
    .O_0_0_2(n22_O_0_0_2),
    .O_1_0_0(n22_O_1_0_0),
    .O_1_0_1(n22_O_1_0_1),
    .O_1_0_2(n22_O_1_0_2),
    .O_2_0_0(n22_O_2_0_0),
    .O_2_0_1(n22_O_2_0_1),
    .O_2_0_2(n22_O_2_0_2),
    .O_3_0_0(n22_O_3_0_0),
    .O_3_0_1(n22_O_3_0_1),
    .O_3_0_2(n22_O_3_0_2),
    .O_4_0_0(n22_O_4_0_0),
    .O_4_0_1(n22_O_4_0_1),
    .O_4_0_2(n22_O_4_0_2),
    .O_5_0_0(n22_O_5_0_0),
    .O_5_0_1(n22_O_5_0_1),
    .O_5_0_2(n22_O_5_0_2),
    .O_6_0_0(n22_O_6_0_0),
    .O_6_0_1(n22_O_6_0_1),
    .O_6_0_2(n22_O_6_0_2),
    .O_7_0_0(n22_O_7_0_0),
    .O_7_0_1(n22_O_7_0_1),
    .O_7_0_2(n22_O_7_0_2),
    .O_8_0_0(n22_O_8_0_0),
    .O_8_0_1(n22_O_8_0_1),
    .O_8_0_2(n22_O_8_0_2),
    .O_9_0_0(n22_O_9_0_0),
    .O_9_0_1(n22_O_9_0_1),
    .O_9_0_2(n22_O_9_0_2),
    .O_10_0_0(n22_O_10_0_0),
    .O_10_0_1(n22_O_10_0_1),
    .O_10_0_2(n22_O_10_0_2),
    .O_11_0_0(n22_O_11_0_0),
    .O_11_0_1(n22_O_11_0_1),
    .O_11_0_2(n22_O_11_0_2),
    .O_12_0_0(n22_O_12_0_0),
    .O_12_0_1(n22_O_12_0_1),
    .O_12_0_2(n22_O_12_0_2),
    .O_13_0_0(n22_O_13_0_0),
    .O_13_0_1(n22_O_13_0_1),
    .O_13_0_2(n22_O_13_0_2),
    .O_14_0_0(n22_O_14_0_0),
    .O_14_0_1(n22_O_14_0_1),
    .O_14_0_2(n22_O_14_0_2),
    .O_15_0_0(n22_O_15_0_0),
    .O_15_0_1(n22_O_15_0_1),
    .O_15_0_2(n22_O_15_0_2)
  );
  MapT_1 n29 ( // @[Top.scala 100:21]
    .valid_up(n29_valid_up),
    .valid_down(n29_valid_down),
    .I_0_0_0(n29_I_0_0_0),
    .I_0_0_1(n29_I_0_0_1),
    .I_0_0_2(n29_I_0_0_2),
    .I_1_0_0(n29_I_1_0_0),
    .I_1_0_1(n29_I_1_0_1),
    .I_1_0_2(n29_I_1_0_2),
    .I_2_0_0(n29_I_2_0_0),
    .I_2_0_1(n29_I_2_0_1),
    .I_2_0_2(n29_I_2_0_2),
    .I_3_0_0(n29_I_3_0_0),
    .I_3_0_1(n29_I_3_0_1),
    .I_3_0_2(n29_I_3_0_2),
    .I_4_0_0(n29_I_4_0_0),
    .I_4_0_1(n29_I_4_0_1),
    .I_4_0_2(n29_I_4_0_2),
    .I_5_0_0(n29_I_5_0_0),
    .I_5_0_1(n29_I_5_0_1),
    .I_5_0_2(n29_I_5_0_2),
    .I_6_0_0(n29_I_6_0_0),
    .I_6_0_1(n29_I_6_0_1),
    .I_6_0_2(n29_I_6_0_2),
    .I_7_0_0(n29_I_7_0_0),
    .I_7_0_1(n29_I_7_0_1),
    .I_7_0_2(n29_I_7_0_2),
    .I_8_0_0(n29_I_8_0_0),
    .I_8_0_1(n29_I_8_0_1),
    .I_8_0_2(n29_I_8_0_2),
    .I_9_0_0(n29_I_9_0_0),
    .I_9_0_1(n29_I_9_0_1),
    .I_9_0_2(n29_I_9_0_2),
    .I_10_0_0(n29_I_10_0_0),
    .I_10_0_1(n29_I_10_0_1),
    .I_10_0_2(n29_I_10_0_2),
    .I_11_0_0(n29_I_11_0_0),
    .I_11_0_1(n29_I_11_0_1),
    .I_11_0_2(n29_I_11_0_2),
    .I_12_0_0(n29_I_12_0_0),
    .I_12_0_1(n29_I_12_0_1),
    .I_12_0_2(n29_I_12_0_2),
    .I_13_0_0(n29_I_13_0_0),
    .I_13_0_1(n29_I_13_0_1),
    .I_13_0_2(n29_I_13_0_2),
    .I_14_0_0(n29_I_14_0_0),
    .I_14_0_1(n29_I_14_0_1),
    .I_14_0_2(n29_I_14_0_2),
    .I_15_0_0(n29_I_15_0_0),
    .I_15_0_1(n29_I_15_0_1),
    .I_15_0_2(n29_I_15_0_2),
    .O_0_0(n29_O_0_0),
    .O_0_1(n29_O_0_1),
    .O_0_2(n29_O_0_2),
    .O_1_0(n29_O_1_0),
    .O_1_1(n29_O_1_1),
    .O_1_2(n29_O_1_2),
    .O_2_0(n29_O_2_0),
    .O_2_1(n29_O_2_1),
    .O_2_2(n29_O_2_2),
    .O_3_0(n29_O_3_0),
    .O_3_1(n29_O_3_1),
    .O_3_2(n29_O_3_2),
    .O_4_0(n29_O_4_0),
    .O_4_1(n29_O_4_1),
    .O_4_2(n29_O_4_2),
    .O_5_0(n29_O_5_0),
    .O_5_1(n29_O_5_1),
    .O_5_2(n29_O_5_2),
    .O_6_0(n29_O_6_0),
    .O_6_1(n29_O_6_1),
    .O_6_2(n29_O_6_2),
    .O_7_0(n29_O_7_0),
    .O_7_1(n29_O_7_1),
    .O_7_2(n29_O_7_2),
    .O_8_0(n29_O_8_0),
    .O_8_1(n29_O_8_1),
    .O_8_2(n29_O_8_2),
    .O_9_0(n29_O_9_0),
    .O_9_1(n29_O_9_1),
    .O_9_2(n29_O_9_2),
    .O_10_0(n29_O_10_0),
    .O_10_1(n29_O_10_1),
    .O_10_2(n29_O_10_2),
    .O_11_0(n29_O_11_0),
    .O_11_1(n29_O_11_1),
    .O_11_2(n29_O_11_2),
    .O_12_0(n29_O_12_0),
    .O_12_1(n29_O_12_1),
    .O_12_2(n29_O_12_2),
    .O_13_0(n29_O_13_0),
    .O_13_1(n29_O_13_1),
    .O_13_2(n29_O_13_2),
    .O_14_0(n29_O_14_0),
    .O_14_1(n29_O_14_1),
    .O_14_2(n29_O_14_2),
    .O_15_0(n29_O_15_0),
    .O_15_1(n29_O_15_1),
    .O_15_2(n29_O_15_2)
  );
  ShiftTS_2 n30 ( // @[Top.scala 103:21]
    .clock(n30_clock),
    .valid_up(n30_valid_up),
    .valid_down(n30_valid_down),
    .I_0(n30_I_0),
    .I_1(n30_I_1),
    .I_2(n30_I_2),
    .I_3(n30_I_3),
    .I_4(n30_I_4),
    .I_5(n30_I_5),
    .I_6(n30_I_6),
    .I_7(n30_I_7),
    .I_8(n30_I_8),
    .I_9(n30_I_9),
    .I_10(n30_I_10),
    .I_11(n30_I_11),
    .I_12(n30_I_12),
    .I_13(n30_I_13),
    .I_14(n30_I_14),
    .I_15(n30_I_15),
    .O_0(n30_O_0),
    .O_1(n30_O_1),
    .O_2(n30_O_2),
    .O_3(n30_O_3),
    .O_4(n30_O_4),
    .O_5(n30_O_5),
    .O_6(n30_O_6),
    .O_7(n30_O_7),
    .O_8(n30_O_8),
    .O_9(n30_O_9),
    .O_10(n30_O_10),
    .O_11(n30_O_11),
    .O_12(n30_O_12),
    .O_13(n30_O_13),
    .O_14(n30_O_14),
    .O_15(n30_O_15)
  );
  ShiftTS_2 n31 ( // @[Top.scala 106:21]
    .clock(n31_clock),
    .valid_up(n31_valid_up),
    .valid_down(n31_valid_down),
    .I_0(n31_I_0),
    .I_1(n31_I_1),
    .I_2(n31_I_2),
    .I_3(n31_I_3),
    .I_4(n31_I_4),
    .I_5(n31_I_5),
    .I_6(n31_I_6),
    .I_7(n31_I_7),
    .I_8(n31_I_8),
    .I_9(n31_I_9),
    .I_10(n31_I_10),
    .I_11(n31_I_11),
    .I_12(n31_I_12),
    .I_13(n31_I_13),
    .I_14(n31_I_14),
    .I_15(n31_I_15),
    .O_0(n31_O_0),
    .O_1(n31_O_1),
    .O_2(n31_O_2),
    .O_3(n31_O_3),
    .O_4(n31_O_4),
    .O_5(n31_O_5),
    .O_6(n31_O_6),
    .O_7(n31_O_7),
    .O_8(n31_O_8),
    .O_9(n31_O_9),
    .O_10(n31_O_10),
    .O_11(n31_O_11),
    .O_12(n31_O_12),
    .O_13(n31_O_13),
    .O_14(n31_O_14),
    .O_15(n31_O_15)
  );
  Map2T n32 ( // @[Top.scala 109:21]
    .valid_up(n32_valid_up),
    .valid_down(n32_valid_down),
    .I0_0(n32_I0_0),
    .I0_1(n32_I0_1),
    .I0_2(n32_I0_2),
    .I0_3(n32_I0_3),
    .I0_4(n32_I0_4),
    .I0_5(n32_I0_5),
    .I0_6(n32_I0_6),
    .I0_7(n32_I0_7),
    .I0_8(n32_I0_8),
    .I0_9(n32_I0_9),
    .I0_10(n32_I0_10),
    .I0_11(n32_I0_11),
    .I0_12(n32_I0_12),
    .I0_13(n32_I0_13),
    .I0_14(n32_I0_14),
    .I0_15(n32_I0_15),
    .I1_0(n32_I1_0),
    .I1_1(n32_I1_1),
    .I1_2(n32_I1_2),
    .I1_3(n32_I1_3),
    .I1_4(n32_I1_4),
    .I1_5(n32_I1_5),
    .I1_6(n32_I1_6),
    .I1_7(n32_I1_7),
    .I1_8(n32_I1_8),
    .I1_9(n32_I1_9),
    .I1_10(n32_I1_10),
    .I1_11(n32_I1_11),
    .I1_12(n32_I1_12),
    .I1_13(n32_I1_13),
    .I1_14(n32_I1_14),
    .I1_15(n32_I1_15),
    .O_0_0(n32_O_0_0),
    .O_0_1(n32_O_0_1),
    .O_1_0(n32_O_1_0),
    .O_1_1(n32_O_1_1),
    .O_2_0(n32_O_2_0),
    .O_2_1(n32_O_2_1),
    .O_3_0(n32_O_3_0),
    .O_3_1(n32_O_3_1),
    .O_4_0(n32_O_4_0),
    .O_4_1(n32_O_4_1),
    .O_5_0(n32_O_5_0),
    .O_5_1(n32_O_5_1),
    .O_6_0(n32_O_6_0),
    .O_6_1(n32_O_6_1),
    .O_7_0(n32_O_7_0),
    .O_7_1(n32_O_7_1),
    .O_8_0(n32_O_8_0),
    .O_8_1(n32_O_8_1),
    .O_9_0(n32_O_9_0),
    .O_9_1(n32_O_9_1),
    .O_10_0(n32_O_10_0),
    .O_10_1(n32_O_10_1),
    .O_11_0(n32_O_11_0),
    .O_11_1(n32_O_11_1),
    .O_12_0(n32_O_12_0),
    .O_12_1(n32_O_12_1),
    .O_13_0(n32_O_13_0),
    .O_13_1(n32_O_13_1),
    .O_14_0(n32_O_14_0),
    .O_14_1(n32_O_14_1),
    .O_15_0(n32_O_15_0),
    .O_15_1(n32_O_15_1)
  );
  Map2T_1 n39 ( // @[Top.scala 113:21]
    .valid_up(n39_valid_up),
    .valid_down(n39_valid_down),
    .I0_0_0(n39_I0_0_0),
    .I0_0_1(n39_I0_0_1),
    .I0_1_0(n39_I0_1_0),
    .I0_1_1(n39_I0_1_1),
    .I0_2_0(n39_I0_2_0),
    .I0_2_1(n39_I0_2_1),
    .I0_3_0(n39_I0_3_0),
    .I0_3_1(n39_I0_3_1),
    .I0_4_0(n39_I0_4_0),
    .I0_4_1(n39_I0_4_1),
    .I0_5_0(n39_I0_5_0),
    .I0_5_1(n39_I0_5_1),
    .I0_6_0(n39_I0_6_0),
    .I0_6_1(n39_I0_6_1),
    .I0_7_0(n39_I0_7_0),
    .I0_7_1(n39_I0_7_1),
    .I0_8_0(n39_I0_8_0),
    .I0_8_1(n39_I0_8_1),
    .I0_9_0(n39_I0_9_0),
    .I0_9_1(n39_I0_9_1),
    .I0_10_0(n39_I0_10_0),
    .I0_10_1(n39_I0_10_1),
    .I0_11_0(n39_I0_11_0),
    .I0_11_1(n39_I0_11_1),
    .I0_12_0(n39_I0_12_0),
    .I0_12_1(n39_I0_12_1),
    .I0_13_0(n39_I0_13_0),
    .I0_13_1(n39_I0_13_1),
    .I0_14_0(n39_I0_14_0),
    .I0_14_1(n39_I0_14_1),
    .I0_15_0(n39_I0_15_0),
    .I0_15_1(n39_I0_15_1),
    .I1_0(n39_I1_0),
    .I1_1(n39_I1_1),
    .I1_2(n39_I1_2),
    .I1_3(n39_I1_3),
    .I1_4(n39_I1_4),
    .I1_5(n39_I1_5),
    .I1_6(n39_I1_6),
    .I1_7(n39_I1_7),
    .I1_8(n39_I1_8),
    .I1_9(n39_I1_9),
    .I1_10(n39_I1_10),
    .I1_11(n39_I1_11),
    .I1_12(n39_I1_12),
    .I1_13(n39_I1_13),
    .I1_14(n39_I1_14),
    .I1_15(n39_I1_15),
    .O_0_0(n39_O_0_0),
    .O_0_1(n39_O_0_1),
    .O_0_2(n39_O_0_2),
    .O_1_0(n39_O_1_0),
    .O_1_1(n39_O_1_1),
    .O_1_2(n39_O_1_2),
    .O_2_0(n39_O_2_0),
    .O_2_1(n39_O_2_1),
    .O_2_2(n39_O_2_2),
    .O_3_0(n39_O_3_0),
    .O_3_1(n39_O_3_1),
    .O_3_2(n39_O_3_2),
    .O_4_0(n39_O_4_0),
    .O_4_1(n39_O_4_1),
    .O_4_2(n39_O_4_2),
    .O_5_0(n39_O_5_0),
    .O_5_1(n39_O_5_1),
    .O_5_2(n39_O_5_2),
    .O_6_0(n39_O_6_0),
    .O_6_1(n39_O_6_1),
    .O_6_2(n39_O_6_2),
    .O_7_0(n39_O_7_0),
    .O_7_1(n39_O_7_1),
    .O_7_2(n39_O_7_2),
    .O_8_0(n39_O_8_0),
    .O_8_1(n39_O_8_1),
    .O_8_2(n39_O_8_2),
    .O_9_0(n39_O_9_0),
    .O_9_1(n39_O_9_1),
    .O_9_2(n39_O_9_2),
    .O_10_0(n39_O_10_0),
    .O_10_1(n39_O_10_1),
    .O_10_2(n39_O_10_2),
    .O_11_0(n39_O_11_0),
    .O_11_1(n39_O_11_1),
    .O_11_2(n39_O_11_2),
    .O_12_0(n39_O_12_0),
    .O_12_1(n39_O_12_1),
    .O_12_2(n39_O_12_2),
    .O_13_0(n39_O_13_0),
    .O_13_1(n39_O_13_1),
    .O_13_2(n39_O_13_2),
    .O_14_0(n39_O_14_0),
    .O_14_1(n39_O_14_1),
    .O_14_2(n39_O_14_2),
    .O_15_0(n39_O_15_0),
    .O_15_1(n39_O_15_1),
    .O_15_2(n39_O_15_2)
  );
  MapT n48 ( // @[Top.scala 117:21]
    .valid_up(n48_valid_up),
    .valid_down(n48_valid_down),
    .I_0_0(n48_I_0_0),
    .I_0_1(n48_I_0_1),
    .I_0_2(n48_I_0_2),
    .I_1_0(n48_I_1_0),
    .I_1_1(n48_I_1_1),
    .I_1_2(n48_I_1_2),
    .I_2_0(n48_I_2_0),
    .I_2_1(n48_I_2_1),
    .I_2_2(n48_I_2_2),
    .I_3_0(n48_I_3_0),
    .I_3_1(n48_I_3_1),
    .I_3_2(n48_I_3_2),
    .I_4_0(n48_I_4_0),
    .I_4_1(n48_I_4_1),
    .I_4_2(n48_I_4_2),
    .I_5_0(n48_I_5_0),
    .I_5_1(n48_I_5_1),
    .I_5_2(n48_I_5_2),
    .I_6_0(n48_I_6_0),
    .I_6_1(n48_I_6_1),
    .I_6_2(n48_I_6_2),
    .I_7_0(n48_I_7_0),
    .I_7_1(n48_I_7_1),
    .I_7_2(n48_I_7_2),
    .I_8_0(n48_I_8_0),
    .I_8_1(n48_I_8_1),
    .I_8_2(n48_I_8_2),
    .I_9_0(n48_I_9_0),
    .I_9_1(n48_I_9_1),
    .I_9_2(n48_I_9_2),
    .I_10_0(n48_I_10_0),
    .I_10_1(n48_I_10_1),
    .I_10_2(n48_I_10_2),
    .I_11_0(n48_I_11_0),
    .I_11_1(n48_I_11_1),
    .I_11_2(n48_I_11_2),
    .I_12_0(n48_I_12_0),
    .I_12_1(n48_I_12_1),
    .I_12_2(n48_I_12_2),
    .I_13_0(n48_I_13_0),
    .I_13_1(n48_I_13_1),
    .I_13_2(n48_I_13_2),
    .I_14_0(n48_I_14_0),
    .I_14_1(n48_I_14_1),
    .I_14_2(n48_I_14_2),
    .I_15_0(n48_I_15_0),
    .I_15_1(n48_I_15_1),
    .I_15_2(n48_I_15_2),
    .O_0_0_0(n48_O_0_0_0),
    .O_0_0_1(n48_O_0_0_1),
    .O_0_0_2(n48_O_0_0_2),
    .O_1_0_0(n48_O_1_0_0),
    .O_1_0_1(n48_O_1_0_1),
    .O_1_0_2(n48_O_1_0_2),
    .O_2_0_0(n48_O_2_0_0),
    .O_2_0_1(n48_O_2_0_1),
    .O_2_0_2(n48_O_2_0_2),
    .O_3_0_0(n48_O_3_0_0),
    .O_3_0_1(n48_O_3_0_1),
    .O_3_0_2(n48_O_3_0_2),
    .O_4_0_0(n48_O_4_0_0),
    .O_4_0_1(n48_O_4_0_1),
    .O_4_0_2(n48_O_4_0_2),
    .O_5_0_0(n48_O_5_0_0),
    .O_5_0_1(n48_O_5_0_1),
    .O_5_0_2(n48_O_5_0_2),
    .O_6_0_0(n48_O_6_0_0),
    .O_6_0_1(n48_O_6_0_1),
    .O_6_0_2(n48_O_6_0_2),
    .O_7_0_0(n48_O_7_0_0),
    .O_7_0_1(n48_O_7_0_1),
    .O_7_0_2(n48_O_7_0_2),
    .O_8_0_0(n48_O_8_0_0),
    .O_8_0_1(n48_O_8_0_1),
    .O_8_0_2(n48_O_8_0_2),
    .O_9_0_0(n48_O_9_0_0),
    .O_9_0_1(n48_O_9_0_1),
    .O_9_0_2(n48_O_9_0_2),
    .O_10_0_0(n48_O_10_0_0),
    .O_10_0_1(n48_O_10_0_1),
    .O_10_0_2(n48_O_10_0_2),
    .O_11_0_0(n48_O_11_0_0),
    .O_11_0_1(n48_O_11_0_1),
    .O_11_0_2(n48_O_11_0_2),
    .O_12_0_0(n48_O_12_0_0),
    .O_12_0_1(n48_O_12_0_1),
    .O_12_0_2(n48_O_12_0_2),
    .O_13_0_0(n48_O_13_0_0),
    .O_13_0_1(n48_O_13_0_1),
    .O_13_0_2(n48_O_13_0_2),
    .O_14_0_0(n48_O_14_0_0),
    .O_14_0_1(n48_O_14_0_1),
    .O_14_0_2(n48_O_14_0_2),
    .O_15_0_0(n48_O_15_0_0),
    .O_15_0_1(n48_O_15_0_1),
    .O_15_0_2(n48_O_15_0_2)
  );
  MapT_1 n55 ( // @[Top.scala 120:21]
    .valid_up(n55_valid_up),
    .valid_down(n55_valid_down),
    .I_0_0_0(n55_I_0_0_0),
    .I_0_0_1(n55_I_0_0_1),
    .I_0_0_2(n55_I_0_0_2),
    .I_1_0_0(n55_I_1_0_0),
    .I_1_0_1(n55_I_1_0_1),
    .I_1_0_2(n55_I_1_0_2),
    .I_2_0_0(n55_I_2_0_0),
    .I_2_0_1(n55_I_2_0_1),
    .I_2_0_2(n55_I_2_0_2),
    .I_3_0_0(n55_I_3_0_0),
    .I_3_0_1(n55_I_3_0_1),
    .I_3_0_2(n55_I_3_0_2),
    .I_4_0_0(n55_I_4_0_0),
    .I_4_0_1(n55_I_4_0_1),
    .I_4_0_2(n55_I_4_0_2),
    .I_5_0_0(n55_I_5_0_0),
    .I_5_0_1(n55_I_5_0_1),
    .I_5_0_2(n55_I_5_0_2),
    .I_6_0_0(n55_I_6_0_0),
    .I_6_0_1(n55_I_6_0_1),
    .I_6_0_2(n55_I_6_0_2),
    .I_7_0_0(n55_I_7_0_0),
    .I_7_0_1(n55_I_7_0_1),
    .I_7_0_2(n55_I_7_0_2),
    .I_8_0_0(n55_I_8_0_0),
    .I_8_0_1(n55_I_8_0_1),
    .I_8_0_2(n55_I_8_0_2),
    .I_9_0_0(n55_I_9_0_0),
    .I_9_0_1(n55_I_9_0_1),
    .I_9_0_2(n55_I_9_0_2),
    .I_10_0_0(n55_I_10_0_0),
    .I_10_0_1(n55_I_10_0_1),
    .I_10_0_2(n55_I_10_0_2),
    .I_11_0_0(n55_I_11_0_0),
    .I_11_0_1(n55_I_11_0_1),
    .I_11_0_2(n55_I_11_0_2),
    .I_12_0_0(n55_I_12_0_0),
    .I_12_0_1(n55_I_12_0_1),
    .I_12_0_2(n55_I_12_0_2),
    .I_13_0_0(n55_I_13_0_0),
    .I_13_0_1(n55_I_13_0_1),
    .I_13_0_2(n55_I_13_0_2),
    .I_14_0_0(n55_I_14_0_0),
    .I_14_0_1(n55_I_14_0_1),
    .I_14_0_2(n55_I_14_0_2),
    .I_15_0_0(n55_I_15_0_0),
    .I_15_0_1(n55_I_15_0_1),
    .I_15_0_2(n55_I_15_0_2),
    .O_0_0(n55_O_0_0),
    .O_0_1(n55_O_0_1),
    .O_0_2(n55_O_0_2),
    .O_1_0(n55_O_1_0),
    .O_1_1(n55_O_1_1),
    .O_1_2(n55_O_1_2),
    .O_2_0(n55_O_2_0),
    .O_2_1(n55_O_2_1),
    .O_2_2(n55_O_2_2),
    .O_3_0(n55_O_3_0),
    .O_3_1(n55_O_3_1),
    .O_3_2(n55_O_3_2),
    .O_4_0(n55_O_4_0),
    .O_4_1(n55_O_4_1),
    .O_4_2(n55_O_4_2),
    .O_5_0(n55_O_5_0),
    .O_5_1(n55_O_5_1),
    .O_5_2(n55_O_5_2),
    .O_6_0(n55_O_6_0),
    .O_6_1(n55_O_6_1),
    .O_6_2(n55_O_6_2),
    .O_7_0(n55_O_7_0),
    .O_7_1(n55_O_7_1),
    .O_7_2(n55_O_7_2),
    .O_8_0(n55_O_8_0),
    .O_8_1(n55_O_8_1),
    .O_8_2(n55_O_8_2),
    .O_9_0(n55_O_9_0),
    .O_9_1(n55_O_9_1),
    .O_9_2(n55_O_9_2),
    .O_10_0(n55_O_10_0),
    .O_10_1(n55_O_10_1),
    .O_10_2(n55_O_10_2),
    .O_11_0(n55_O_11_0),
    .O_11_1(n55_O_11_1),
    .O_11_2(n55_O_11_2),
    .O_12_0(n55_O_12_0),
    .O_12_1(n55_O_12_1),
    .O_12_2(n55_O_12_2),
    .O_13_0(n55_O_13_0),
    .O_13_1(n55_O_13_1),
    .O_13_2(n55_O_13_2),
    .O_14_0(n55_O_14_0),
    .O_14_1(n55_O_14_1),
    .O_14_2(n55_O_14_2),
    .O_15_0(n55_O_15_0),
    .O_15_1(n55_O_15_1),
    .O_15_2(n55_O_15_2)
  );
  Map2T_4 n56 ( // @[Top.scala 123:21]
    .valid_up(n56_valid_up),
    .valid_down(n56_valid_down),
    .I0_0_0(n56_I0_0_0),
    .I0_0_1(n56_I0_0_1),
    .I0_0_2(n56_I0_0_2),
    .I0_1_0(n56_I0_1_0),
    .I0_1_1(n56_I0_1_1),
    .I0_1_2(n56_I0_1_2),
    .I0_2_0(n56_I0_2_0),
    .I0_2_1(n56_I0_2_1),
    .I0_2_2(n56_I0_2_2),
    .I0_3_0(n56_I0_3_0),
    .I0_3_1(n56_I0_3_1),
    .I0_3_2(n56_I0_3_2),
    .I0_4_0(n56_I0_4_0),
    .I0_4_1(n56_I0_4_1),
    .I0_4_2(n56_I0_4_2),
    .I0_5_0(n56_I0_5_0),
    .I0_5_1(n56_I0_5_1),
    .I0_5_2(n56_I0_5_2),
    .I0_6_0(n56_I0_6_0),
    .I0_6_1(n56_I0_6_1),
    .I0_6_2(n56_I0_6_2),
    .I0_7_0(n56_I0_7_0),
    .I0_7_1(n56_I0_7_1),
    .I0_7_2(n56_I0_7_2),
    .I0_8_0(n56_I0_8_0),
    .I0_8_1(n56_I0_8_1),
    .I0_8_2(n56_I0_8_2),
    .I0_9_0(n56_I0_9_0),
    .I0_9_1(n56_I0_9_1),
    .I0_9_2(n56_I0_9_2),
    .I0_10_0(n56_I0_10_0),
    .I0_10_1(n56_I0_10_1),
    .I0_10_2(n56_I0_10_2),
    .I0_11_0(n56_I0_11_0),
    .I0_11_1(n56_I0_11_1),
    .I0_11_2(n56_I0_11_2),
    .I0_12_0(n56_I0_12_0),
    .I0_12_1(n56_I0_12_1),
    .I0_12_2(n56_I0_12_2),
    .I0_13_0(n56_I0_13_0),
    .I0_13_1(n56_I0_13_1),
    .I0_13_2(n56_I0_13_2),
    .I0_14_0(n56_I0_14_0),
    .I0_14_1(n56_I0_14_1),
    .I0_14_2(n56_I0_14_2),
    .I0_15_0(n56_I0_15_0),
    .I0_15_1(n56_I0_15_1),
    .I0_15_2(n56_I0_15_2),
    .I1_0_0(n56_I1_0_0),
    .I1_0_1(n56_I1_0_1),
    .I1_0_2(n56_I1_0_2),
    .I1_1_0(n56_I1_1_0),
    .I1_1_1(n56_I1_1_1),
    .I1_1_2(n56_I1_1_2),
    .I1_2_0(n56_I1_2_0),
    .I1_2_1(n56_I1_2_1),
    .I1_2_2(n56_I1_2_2),
    .I1_3_0(n56_I1_3_0),
    .I1_3_1(n56_I1_3_1),
    .I1_3_2(n56_I1_3_2),
    .I1_4_0(n56_I1_4_0),
    .I1_4_1(n56_I1_4_1),
    .I1_4_2(n56_I1_4_2),
    .I1_5_0(n56_I1_5_0),
    .I1_5_1(n56_I1_5_1),
    .I1_5_2(n56_I1_5_2),
    .I1_6_0(n56_I1_6_0),
    .I1_6_1(n56_I1_6_1),
    .I1_6_2(n56_I1_6_2),
    .I1_7_0(n56_I1_7_0),
    .I1_7_1(n56_I1_7_1),
    .I1_7_2(n56_I1_7_2),
    .I1_8_0(n56_I1_8_0),
    .I1_8_1(n56_I1_8_1),
    .I1_8_2(n56_I1_8_2),
    .I1_9_0(n56_I1_9_0),
    .I1_9_1(n56_I1_9_1),
    .I1_9_2(n56_I1_9_2),
    .I1_10_0(n56_I1_10_0),
    .I1_10_1(n56_I1_10_1),
    .I1_10_2(n56_I1_10_2),
    .I1_11_0(n56_I1_11_0),
    .I1_11_1(n56_I1_11_1),
    .I1_11_2(n56_I1_11_2),
    .I1_12_0(n56_I1_12_0),
    .I1_12_1(n56_I1_12_1),
    .I1_12_2(n56_I1_12_2),
    .I1_13_0(n56_I1_13_0),
    .I1_13_1(n56_I1_13_1),
    .I1_13_2(n56_I1_13_2),
    .I1_14_0(n56_I1_14_0),
    .I1_14_1(n56_I1_14_1),
    .I1_14_2(n56_I1_14_2),
    .I1_15_0(n56_I1_15_0),
    .I1_15_1(n56_I1_15_1),
    .I1_15_2(n56_I1_15_2),
    .O_0_0_0(n56_O_0_0_0),
    .O_0_0_1(n56_O_0_0_1),
    .O_0_0_2(n56_O_0_0_2),
    .O_0_1_0(n56_O_0_1_0),
    .O_0_1_1(n56_O_0_1_1),
    .O_0_1_2(n56_O_0_1_2),
    .O_1_0_0(n56_O_1_0_0),
    .O_1_0_1(n56_O_1_0_1),
    .O_1_0_2(n56_O_1_0_2),
    .O_1_1_0(n56_O_1_1_0),
    .O_1_1_1(n56_O_1_1_1),
    .O_1_1_2(n56_O_1_1_2),
    .O_2_0_0(n56_O_2_0_0),
    .O_2_0_1(n56_O_2_0_1),
    .O_2_0_2(n56_O_2_0_2),
    .O_2_1_0(n56_O_2_1_0),
    .O_2_1_1(n56_O_2_1_1),
    .O_2_1_2(n56_O_2_1_2),
    .O_3_0_0(n56_O_3_0_0),
    .O_3_0_1(n56_O_3_0_1),
    .O_3_0_2(n56_O_3_0_2),
    .O_3_1_0(n56_O_3_1_0),
    .O_3_1_1(n56_O_3_1_1),
    .O_3_1_2(n56_O_3_1_2),
    .O_4_0_0(n56_O_4_0_0),
    .O_4_0_1(n56_O_4_0_1),
    .O_4_0_2(n56_O_4_0_2),
    .O_4_1_0(n56_O_4_1_0),
    .O_4_1_1(n56_O_4_1_1),
    .O_4_1_2(n56_O_4_1_2),
    .O_5_0_0(n56_O_5_0_0),
    .O_5_0_1(n56_O_5_0_1),
    .O_5_0_2(n56_O_5_0_2),
    .O_5_1_0(n56_O_5_1_0),
    .O_5_1_1(n56_O_5_1_1),
    .O_5_1_2(n56_O_5_1_2),
    .O_6_0_0(n56_O_6_0_0),
    .O_6_0_1(n56_O_6_0_1),
    .O_6_0_2(n56_O_6_0_2),
    .O_6_1_0(n56_O_6_1_0),
    .O_6_1_1(n56_O_6_1_1),
    .O_6_1_2(n56_O_6_1_2),
    .O_7_0_0(n56_O_7_0_0),
    .O_7_0_1(n56_O_7_0_1),
    .O_7_0_2(n56_O_7_0_2),
    .O_7_1_0(n56_O_7_1_0),
    .O_7_1_1(n56_O_7_1_1),
    .O_7_1_2(n56_O_7_1_2),
    .O_8_0_0(n56_O_8_0_0),
    .O_8_0_1(n56_O_8_0_1),
    .O_8_0_2(n56_O_8_0_2),
    .O_8_1_0(n56_O_8_1_0),
    .O_8_1_1(n56_O_8_1_1),
    .O_8_1_2(n56_O_8_1_2),
    .O_9_0_0(n56_O_9_0_0),
    .O_9_0_1(n56_O_9_0_1),
    .O_9_0_2(n56_O_9_0_2),
    .O_9_1_0(n56_O_9_1_0),
    .O_9_1_1(n56_O_9_1_1),
    .O_9_1_2(n56_O_9_1_2),
    .O_10_0_0(n56_O_10_0_0),
    .O_10_0_1(n56_O_10_0_1),
    .O_10_0_2(n56_O_10_0_2),
    .O_10_1_0(n56_O_10_1_0),
    .O_10_1_1(n56_O_10_1_1),
    .O_10_1_2(n56_O_10_1_2),
    .O_11_0_0(n56_O_11_0_0),
    .O_11_0_1(n56_O_11_0_1),
    .O_11_0_2(n56_O_11_0_2),
    .O_11_1_0(n56_O_11_1_0),
    .O_11_1_1(n56_O_11_1_1),
    .O_11_1_2(n56_O_11_1_2),
    .O_12_0_0(n56_O_12_0_0),
    .O_12_0_1(n56_O_12_0_1),
    .O_12_0_2(n56_O_12_0_2),
    .O_12_1_0(n56_O_12_1_0),
    .O_12_1_1(n56_O_12_1_1),
    .O_12_1_2(n56_O_12_1_2),
    .O_13_0_0(n56_O_13_0_0),
    .O_13_0_1(n56_O_13_0_1),
    .O_13_0_2(n56_O_13_0_2),
    .O_13_1_0(n56_O_13_1_0),
    .O_13_1_1(n56_O_13_1_1),
    .O_13_1_2(n56_O_13_1_2),
    .O_14_0_0(n56_O_14_0_0),
    .O_14_0_1(n56_O_14_0_1),
    .O_14_0_2(n56_O_14_0_2),
    .O_14_1_0(n56_O_14_1_0),
    .O_14_1_1(n56_O_14_1_1),
    .O_14_1_2(n56_O_14_1_2),
    .O_15_0_0(n56_O_15_0_0),
    .O_15_0_1(n56_O_15_0_1),
    .O_15_0_2(n56_O_15_0_2),
    .O_15_1_0(n56_O_15_1_0),
    .O_15_1_1(n56_O_15_1_1),
    .O_15_1_2(n56_O_15_1_2)
  );
  ShiftTS_2 n63 ( // @[Top.scala 127:21]
    .clock(n63_clock),
    .valid_up(n63_valid_up),
    .valid_down(n63_valid_down),
    .I_0(n63_I_0),
    .I_1(n63_I_1),
    .I_2(n63_I_2),
    .I_3(n63_I_3),
    .I_4(n63_I_4),
    .I_5(n63_I_5),
    .I_6(n63_I_6),
    .I_7(n63_I_7),
    .I_8(n63_I_8),
    .I_9(n63_I_9),
    .I_10(n63_I_10),
    .I_11(n63_I_11),
    .I_12(n63_I_12),
    .I_13(n63_I_13),
    .I_14(n63_I_14),
    .I_15(n63_I_15),
    .O_0(n63_O_0),
    .O_1(n63_O_1),
    .O_2(n63_O_2),
    .O_3(n63_O_3),
    .O_4(n63_O_4),
    .O_5(n63_O_5),
    .O_6(n63_O_6),
    .O_7(n63_O_7),
    .O_8(n63_O_8),
    .O_9(n63_O_9),
    .O_10(n63_O_10),
    .O_11(n63_O_11),
    .O_12(n63_O_12),
    .O_13(n63_O_13),
    .O_14(n63_O_14),
    .O_15(n63_O_15)
  );
  ShiftTS_2 n64 ( // @[Top.scala 130:21]
    .clock(n64_clock),
    .valid_up(n64_valid_up),
    .valid_down(n64_valid_down),
    .I_0(n64_I_0),
    .I_1(n64_I_1),
    .I_2(n64_I_2),
    .I_3(n64_I_3),
    .I_4(n64_I_4),
    .I_5(n64_I_5),
    .I_6(n64_I_6),
    .I_7(n64_I_7),
    .I_8(n64_I_8),
    .I_9(n64_I_9),
    .I_10(n64_I_10),
    .I_11(n64_I_11),
    .I_12(n64_I_12),
    .I_13(n64_I_13),
    .I_14(n64_I_14),
    .I_15(n64_I_15),
    .O_0(n64_O_0),
    .O_1(n64_O_1),
    .O_2(n64_O_2),
    .O_3(n64_O_3),
    .O_4(n64_O_4),
    .O_5(n64_O_5),
    .O_6(n64_O_6),
    .O_7(n64_O_7),
    .O_8(n64_O_8),
    .O_9(n64_O_9),
    .O_10(n64_O_10),
    .O_11(n64_O_11),
    .O_12(n64_O_12),
    .O_13(n64_O_13),
    .O_14(n64_O_14),
    .O_15(n64_O_15)
  );
  Map2T n65 ( // @[Top.scala 133:21]
    .valid_up(n65_valid_up),
    .valid_down(n65_valid_down),
    .I0_0(n65_I0_0),
    .I0_1(n65_I0_1),
    .I0_2(n65_I0_2),
    .I0_3(n65_I0_3),
    .I0_4(n65_I0_4),
    .I0_5(n65_I0_5),
    .I0_6(n65_I0_6),
    .I0_7(n65_I0_7),
    .I0_8(n65_I0_8),
    .I0_9(n65_I0_9),
    .I0_10(n65_I0_10),
    .I0_11(n65_I0_11),
    .I0_12(n65_I0_12),
    .I0_13(n65_I0_13),
    .I0_14(n65_I0_14),
    .I0_15(n65_I0_15),
    .I1_0(n65_I1_0),
    .I1_1(n65_I1_1),
    .I1_2(n65_I1_2),
    .I1_3(n65_I1_3),
    .I1_4(n65_I1_4),
    .I1_5(n65_I1_5),
    .I1_6(n65_I1_6),
    .I1_7(n65_I1_7),
    .I1_8(n65_I1_8),
    .I1_9(n65_I1_9),
    .I1_10(n65_I1_10),
    .I1_11(n65_I1_11),
    .I1_12(n65_I1_12),
    .I1_13(n65_I1_13),
    .I1_14(n65_I1_14),
    .I1_15(n65_I1_15),
    .O_0_0(n65_O_0_0),
    .O_0_1(n65_O_0_1),
    .O_1_0(n65_O_1_0),
    .O_1_1(n65_O_1_1),
    .O_2_0(n65_O_2_0),
    .O_2_1(n65_O_2_1),
    .O_3_0(n65_O_3_0),
    .O_3_1(n65_O_3_1),
    .O_4_0(n65_O_4_0),
    .O_4_1(n65_O_4_1),
    .O_5_0(n65_O_5_0),
    .O_5_1(n65_O_5_1),
    .O_6_0(n65_O_6_0),
    .O_6_1(n65_O_6_1),
    .O_7_0(n65_O_7_0),
    .O_7_1(n65_O_7_1),
    .O_8_0(n65_O_8_0),
    .O_8_1(n65_O_8_1),
    .O_9_0(n65_O_9_0),
    .O_9_1(n65_O_9_1),
    .O_10_0(n65_O_10_0),
    .O_10_1(n65_O_10_1),
    .O_11_0(n65_O_11_0),
    .O_11_1(n65_O_11_1),
    .O_12_0(n65_O_12_0),
    .O_12_1(n65_O_12_1),
    .O_13_0(n65_O_13_0),
    .O_13_1(n65_O_13_1),
    .O_14_0(n65_O_14_0),
    .O_14_1(n65_O_14_1),
    .O_15_0(n65_O_15_0),
    .O_15_1(n65_O_15_1)
  );
  Map2T_1 n72 ( // @[Top.scala 137:21]
    .valid_up(n72_valid_up),
    .valid_down(n72_valid_down),
    .I0_0_0(n72_I0_0_0),
    .I0_0_1(n72_I0_0_1),
    .I0_1_0(n72_I0_1_0),
    .I0_1_1(n72_I0_1_1),
    .I0_2_0(n72_I0_2_0),
    .I0_2_1(n72_I0_2_1),
    .I0_3_0(n72_I0_3_0),
    .I0_3_1(n72_I0_3_1),
    .I0_4_0(n72_I0_4_0),
    .I0_4_1(n72_I0_4_1),
    .I0_5_0(n72_I0_5_0),
    .I0_5_1(n72_I0_5_1),
    .I0_6_0(n72_I0_6_0),
    .I0_6_1(n72_I0_6_1),
    .I0_7_0(n72_I0_7_0),
    .I0_7_1(n72_I0_7_1),
    .I0_8_0(n72_I0_8_0),
    .I0_8_1(n72_I0_8_1),
    .I0_9_0(n72_I0_9_0),
    .I0_9_1(n72_I0_9_1),
    .I0_10_0(n72_I0_10_0),
    .I0_10_1(n72_I0_10_1),
    .I0_11_0(n72_I0_11_0),
    .I0_11_1(n72_I0_11_1),
    .I0_12_0(n72_I0_12_0),
    .I0_12_1(n72_I0_12_1),
    .I0_13_0(n72_I0_13_0),
    .I0_13_1(n72_I0_13_1),
    .I0_14_0(n72_I0_14_0),
    .I0_14_1(n72_I0_14_1),
    .I0_15_0(n72_I0_15_0),
    .I0_15_1(n72_I0_15_1),
    .I1_0(n72_I1_0),
    .I1_1(n72_I1_1),
    .I1_2(n72_I1_2),
    .I1_3(n72_I1_3),
    .I1_4(n72_I1_4),
    .I1_5(n72_I1_5),
    .I1_6(n72_I1_6),
    .I1_7(n72_I1_7),
    .I1_8(n72_I1_8),
    .I1_9(n72_I1_9),
    .I1_10(n72_I1_10),
    .I1_11(n72_I1_11),
    .I1_12(n72_I1_12),
    .I1_13(n72_I1_13),
    .I1_14(n72_I1_14),
    .I1_15(n72_I1_15),
    .O_0_0(n72_O_0_0),
    .O_0_1(n72_O_0_1),
    .O_0_2(n72_O_0_2),
    .O_1_0(n72_O_1_0),
    .O_1_1(n72_O_1_1),
    .O_1_2(n72_O_1_2),
    .O_2_0(n72_O_2_0),
    .O_2_1(n72_O_2_1),
    .O_2_2(n72_O_2_2),
    .O_3_0(n72_O_3_0),
    .O_3_1(n72_O_3_1),
    .O_3_2(n72_O_3_2),
    .O_4_0(n72_O_4_0),
    .O_4_1(n72_O_4_1),
    .O_4_2(n72_O_4_2),
    .O_5_0(n72_O_5_0),
    .O_5_1(n72_O_5_1),
    .O_5_2(n72_O_5_2),
    .O_6_0(n72_O_6_0),
    .O_6_1(n72_O_6_1),
    .O_6_2(n72_O_6_2),
    .O_7_0(n72_O_7_0),
    .O_7_1(n72_O_7_1),
    .O_7_2(n72_O_7_2),
    .O_8_0(n72_O_8_0),
    .O_8_1(n72_O_8_1),
    .O_8_2(n72_O_8_2),
    .O_9_0(n72_O_9_0),
    .O_9_1(n72_O_9_1),
    .O_9_2(n72_O_9_2),
    .O_10_0(n72_O_10_0),
    .O_10_1(n72_O_10_1),
    .O_10_2(n72_O_10_2),
    .O_11_0(n72_O_11_0),
    .O_11_1(n72_O_11_1),
    .O_11_2(n72_O_11_2),
    .O_12_0(n72_O_12_0),
    .O_12_1(n72_O_12_1),
    .O_12_2(n72_O_12_2),
    .O_13_0(n72_O_13_0),
    .O_13_1(n72_O_13_1),
    .O_13_2(n72_O_13_2),
    .O_14_0(n72_O_14_0),
    .O_14_1(n72_O_14_1),
    .O_14_2(n72_O_14_2),
    .O_15_0(n72_O_15_0),
    .O_15_1(n72_O_15_1),
    .O_15_2(n72_O_15_2)
  );
  MapT n81 ( // @[Top.scala 141:21]
    .valid_up(n81_valid_up),
    .valid_down(n81_valid_down),
    .I_0_0(n81_I_0_0),
    .I_0_1(n81_I_0_1),
    .I_0_2(n81_I_0_2),
    .I_1_0(n81_I_1_0),
    .I_1_1(n81_I_1_1),
    .I_1_2(n81_I_1_2),
    .I_2_0(n81_I_2_0),
    .I_2_1(n81_I_2_1),
    .I_2_2(n81_I_2_2),
    .I_3_0(n81_I_3_0),
    .I_3_1(n81_I_3_1),
    .I_3_2(n81_I_3_2),
    .I_4_0(n81_I_4_0),
    .I_4_1(n81_I_4_1),
    .I_4_2(n81_I_4_2),
    .I_5_0(n81_I_5_0),
    .I_5_1(n81_I_5_1),
    .I_5_2(n81_I_5_2),
    .I_6_0(n81_I_6_0),
    .I_6_1(n81_I_6_1),
    .I_6_2(n81_I_6_2),
    .I_7_0(n81_I_7_0),
    .I_7_1(n81_I_7_1),
    .I_7_2(n81_I_7_2),
    .I_8_0(n81_I_8_0),
    .I_8_1(n81_I_8_1),
    .I_8_2(n81_I_8_2),
    .I_9_0(n81_I_9_0),
    .I_9_1(n81_I_9_1),
    .I_9_2(n81_I_9_2),
    .I_10_0(n81_I_10_0),
    .I_10_1(n81_I_10_1),
    .I_10_2(n81_I_10_2),
    .I_11_0(n81_I_11_0),
    .I_11_1(n81_I_11_1),
    .I_11_2(n81_I_11_2),
    .I_12_0(n81_I_12_0),
    .I_12_1(n81_I_12_1),
    .I_12_2(n81_I_12_2),
    .I_13_0(n81_I_13_0),
    .I_13_1(n81_I_13_1),
    .I_13_2(n81_I_13_2),
    .I_14_0(n81_I_14_0),
    .I_14_1(n81_I_14_1),
    .I_14_2(n81_I_14_2),
    .I_15_0(n81_I_15_0),
    .I_15_1(n81_I_15_1),
    .I_15_2(n81_I_15_2),
    .O_0_0_0(n81_O_0_0_0),
    .O_0_0_1(n81_O_0_0_1),
    .O_0_0_2(n81_O_0_0_2),
    .O_1_0_0(n81_O_1_0_0),
    .O_1_0_1(n81_O_1_0_1),
    .O_1_0_2(n81_O_1_0_2),
    .O_2_0_0(n81_O_2_0_0),
    .O_2_0_1(n81_O_2_0_1),
    .O_2_0_2(n81_O_2_0_2),
    .O_3_0_0(n81_O_3_0_0),
    .O_3_0_1(n81_O_3_0_1),
    .O_3_0_2(n81_O_3_0_2),
    .O_4_0_0(n81_O_4_0_0),
    .O_4_0_1(n81_O_4_0_1),
    .O_4_0_2(n81_O_4_0_2),
    .O_5_0_0(n81_O_5_0_0),
    .O_5_0_1(n81_O_5_0_1),
    .O_5_0_2(n81_O_5_0_2),
    .O_6_0_0(n81_O_6_0_0),
    .O_6_0_1(n81_O_6_0_1),
    .O_6_0_2(n81_O_6_0_2),
    .O_7_0_0(n81_O_7_0_0),
    .O_7_0_1(n81_O_7_0_1),
    .O_7_0_2(n81_O_7_0_2),
    .O_8_0_0(n81_O_8_0_0),
    .O_8_0_1(n81_O_8_0_1),
    .O_8_0_2(n81_O_8_0_2),
    .O_9_0_0(n81_O_9_0_0),
    .O_9_0_1(n81_O_9_0_1),
    .O_9_0_2(n81_O_9_0_2),
    .O_10_0_0(n81_O_10_0_0),
    .O_10_0_1(n81_O_10_0_1),
    .O_10_0_2(n81_O_10_0_2),
    .O_11_0_0(n81_O_11_0_0),
    .O_11_0_1(n81_O_11_0_1),
    .O_11_0_2(n81_O_11_0_2),
    .O_12_0_0(n81_O_12_0_0),
    .O_12_0_1(n81_O_12_0_1),
    .O_12_0_2(n81_O_12_0_2),
    .O_13_0_0(n81_O_13_0_0),
    .O_13_0_1(n81_O_13_0_1),
    .O_13_0_2(n81_O_13_0_2),
    .O_14_0_0(n81_O_14_0_0),
    .O_14_0_1(n81_O_14_0_1),
    .O_14_0_2(n81_O_14_0_2),
    .O_15_0_0(n81_O_15_0_0),
    .O_15_0_1(n81_O_15_0_1),
    .O_15_0_2(n81_O_15_0_2)
  );
  MapT_1 n88 ( // @[Top.scala 144:21]
    .valid_up(n88_valid_up),
    .valid_down(n88_valid_down),
    .I_0_0_0(n88_I_0_0_0),
    .I_0_0_1(n88_I_0_0_1),
    .I_0_0_2(n88_I_0_0_2),
    .I_1_0_0(n88_I_1_0_0),
    .I_1_0_1(n88_I_1_0_1),
    .I_1_0_2(n88_I_1_0_2),
    .I_2_0_0(n88_I_2_0_0),
    .I_2_0_1(n88_I_2_0_1),
    .I_2_0_2(n88_I_2_0_2),
    .I_3_0_0(n88_I_3_0_0),
    .I_3_0_1(n88_I_3_0_1),
    .I_3_0_2(n88_I_3_0_2),
    .I_4_0_0(n88_I_4_0_0),
    .I_4_0_1(n88_I_4_0_1),
    .I_4_0_2(n88_I_4_0_2),
    .I_5_0_0(n88_I_5_0_0),
    .I_5_0_1(n88_I_5_0_1),
    .I_5_0_2(n88_I_5_0_2),
    .I_6_0_0(n88_I_6_0_0),
    .I_6_0_1(n88_I_6_0_1),
    .I_6_0_2(n88_I_6_0_2),
    .I_7_0_0(n88_I_7_0_0),
    .I_7_0_1(n88_I_7_0_1),
    .I_7_0_2(n88_I_7_0_2),
    .I_8_0_0(n88_I_8_0_0),
    .I_8_0_1(n88_I_8_0_1),
    .I_8_0_2(n88_I_8_0_2),
    .I_9_0_0(n88_I_9_0_0),
    .I_9_0_1(n88_I_9_0_1),
    .I_9_0_2(n88_I_9_0_2),
    .I_10_0_0(n88_I_10_0_0),
    .I_10_0_1(n88_I_10_0_1),
    .I_10_0_2(n88_I_10_0_2),
    .I_11_0_0(n88_I_11_0_0),
    .I_11_0_1(n88_I_11_0_1),
    .I_11_0_2(n88_I_11_0_2),
    .I_12_0_0(n88_I_12_0_0),
    .I_12_0_1(n88_I_12_0_1),
    .I_12_0_2(n88_I_12_0_2),
    .I_13_0_0(n88_I_13_0_0),
    .I_13_0_1(n88_I_13_0_1),
    .I_13_0_2(n88_I_13_0_2),
    .I_14_0_0(n88_I_14_0_0),
    .I_14_0_1(n88_I_14_0_1),
    .I_14_0_2(n88_I_14_0_2),
    .I_15_0_0(n88_I_15_0_0),
    .I_15_0_1(n88_I_15_0_1),
    .I_15_0_2(n88_I_15_0_2),
    .O_0_0(n88_O_0_0),
    .O_0_1(n88_O_0_1),
    .O_0_2(n88_O_0_2),
    .O_1_0(n88_O_1_0),
    .O_1_1(n88_O_1_1),
    .O_1_2(n88_O_1_2),
    .O_2_0(n88_O_2_0),
    .O_2_1(n88_O_2_1),
    .O_2_2(n88_O_2_2),
    .O_3_0(n88_O_3_0),
    .O_3_1(n88_O_3_1),
    .O_3_2(n88_O_3_2),
    .O_4_0(n88_O_4_0),
    .O_4_1(n88_O_4_1),
    .O_4_2(n88_O_4_2),
    .O_5_0(n88_O_5_0),
    .O_5_1(n88_O_5_1),
    .O_5_2(n88_O_5_2),
    .O_6_0(n88_O_6_0),
    .O_6_1(n88_O_6_1),
    .O_6_2(n88_O_6_2),
    .O_7_0(n88_O_7_0),
    .O_7_1(n88_O_7_1),
    .O_7_2(n88_O_7_2),
    .O_8_0(n88_O_8_0),
    .O_8_1(n88_O_8_1),
    .O_8_2(n88_O_8_2),
    .O_9_0(n88_O_9_0),
    .O_9_1(n88_O_9_1),
    .O_9_2(n88_O_9_2),
    .O_10_0(n88_O_10_0),
    .O_10_1(n88_O_10_1),
    .O_10_2(n88_O_10_2),
    .O_11_0(n88_O_11_0),
    .O_11_1(n88_O_11_1),
    .O_11_2(n88_O_11_2),
    .O_12_0(n88_O_12_0),
    .O_12_1(n88_O_12_1),
    .O_12_2(n88_O_12_2),
    .O_13_0(n88_O_13_0),
    .O_13_1(n88_O_13_1),
    .O_13_2(n88_O_13_2),
    .O_14_0(n88_O_14_0),
    .O_14_1(n88_O_14_1),
    .O_14_2(n88_O_14_2),
    .O_15_0(n88_O_15_0),
    .O_15_1(n88_O_15_1),
    .O_15_2(n88_O_15_2)
  );
  Map2T_7 n89 ( // @[Top.scala 147:21]
    .valid_up(n89_valid_up),
    .valid_down(n89_valid_down),
    .I0_0_0_0(n89_I0_0_0_0),
    .I0_0_0_1(n89_I0_0_0_1),
    .I0_0_0_2(n89_I0_0_0_2),
    .I0_0_1_0(n89_I0_0_1_0),
    .I0_0_1_1(n89_I0_0_1_1),
    .I0_0_1_2(n89_I0_0_1_2),
    .I0_1_0_0(n89_I0_1_0_0),
    .I0_1_0_1(n89_I0_1_0_1),
    .I0_1_0_2(n89_I0_1_0_2),
    .I0_1_1_0(n89_I0_1_1_0),
    .I0_1_1_1(n89_I0_1_1_1),
    .I0_1_1_2(n89_I0_1_1_2),
    .I0_2_0_0(n89_I0_2_0_0),
    .I0_2_0_1(n89_I0_2_0_1),
    .I0_2_0_2(n89_I0_2_0_2),
    .I0_2_1_0(n89_I0_2_1_0),
    .I0_2_1_1(n89_I0_2_1_1),
    .I0_2_1_2(n89_I0_2_1_2),
    .I0_3_0_0(n89_I0_3_0_0),
    .I0_3_0_1(n89_I0_3_0_1),
    .I0_3_0_2(n89_I0_3_0_2),
    .I0_3_1_0(n89_I0_3_1_0),
    .I0_3_1_1(n89_I0_3_1_1),
    .I0_3_1_2(n89_I0_3_1_2),
    .I0_4_0_0(n89_I0_4_0_0),
    .I0_4_0_1(n89_I0_4_0_1),
    .I0_4_0_2(n89_I0_4_0_2),
    .I0_4_1_0(n89_I0_4_1_0),
    .I0_4_1_1(n89_I0_4_1_1),
    .I0_4_1_2(n89_I0_4_1_2),
    .I0_5_0_0(n89_I0_5_0_0),
    .I0_5_0_1(n89_I0_5_0_1),
    .I0_5_0_2(n89_I0_5_0_2),
    .I0_5_1_0(n89_I0_5_1_0),
    .I0_5_1_1(n89_I0_5_1_1),
    .I0_5_1_2(n89_I0_5_1_2),
    .I0_6_0_0(n89_I0_6_0_0),
    .I0_6_0_1(n89_I0_6_0_1),
    .I0_6_0_2(n89_I0_6_0_2),
    .I0_6_1_0(n89_I0_6_1_0),
    .I0_6_1_1(n89_I0_6_1_1),
    .I0_6_1_2(n89_I0_6_1_2),
    .I0_7_0_0(n89_I0_7_0_0),
    .I0_7_0_1(n89_I0_7_0_1),
    .I0_7_0_2(n89_I0_7_0_2),
    .I0_7_1_0(n89_I0_7_1_0),
    .I0_7_1_1(n89_I0_7_1_1),
    .I0_7_1_2(n89_I0_7_1_2),
    .I0_8_0_0(n89_I0_8_0_0),
    .I0_8_0_1(n89_I0_8_0_1),
    .I0_8_0_2(n89_I0_8_0_2),
    .I0_8_1_0(n89_I0_8_1_0),
    .I0_8_1_1(n89_I0_8_1_1),
    .I0_8_1_2(n89_I0_8_1_2),
    .I0_9_0_0(n89_I0_9_0_0),
    .I0_9_0_1(n89_I0_9_0_1),
    .I0_9_0_2(n89_I0_9_0_2),
    .I0_9_1_0(n89_I0_9_1_0),
    .I0_9_1_1(n89_I0_9_1_1),
    .I0_9_1_2(n89_I0_9_1_2),
    .I0_10_0_0(n89_I0_10_0_0),
    .I0_10_0_1(n89_I0_10_0_1),
    .I0_10_0_2(n89_I0_10_0_2),
    .I0_10_1_0(n89_I0_10_1_0),
    .I0_10_1_1(n89_I0_10_1_1),
    .I0_10_1_2(n89_I0_10_1_2),
    .I0_11_0_0(n89_I0_11_0_0),
    .I0_11_0_1(n89_I0_11_0_1),
    .I0_11_0_2(n89_I0_11_0_2),
    .I0_11_1_0(n89_I0_11_1_0),
    .I0_11_1_1(n89_I0_11_1_1),
    .I0_11_1_2(n89_I0_11_1_2),
    .I0_12_0_0(n89_I0_12_0_0),
    .I0_12_0_1(n89_I0_12_0_1),
    .I0_12_0_2(n89_I0_12_0_2),
    .I0_12_1_0(n89_I0_12_1_0),
    .I0_12_1_1(n89_I0_12_1_1),
    .I0_12_1_2(n89_I0_12_1_2),
    .I0_13_0_0(n89_I0_13_0_0),
    .I0_13_0_1(n89_I0_13_0_1),
    .I0_13_0_2(n89_I0_13_0_2),
    .I0_13_1_0(n89_I0_13_1_0),
    .I0_13_1_1(n89_I0_13_1_1),
    .I0_13_1_2(n89_I0_13_1_2),
    .I0_14_0_0(n89_I0_14_0_0),
    .I0_14_0_1(n89_I0_14_0_1),
    .I0_14_0_2(n89_I0_14_0_2),
    .I0_14_1_0(n89_I0_14_1_0),
    .I0_14_1_1(n89_I0_14_1_1),
    .I0_14_1_2(n89_I0_14_1_2),
    .I0_15_0_0(n89_I0_15_0_0),
    .I0_15_0_1(n89_I0_15_0_1),
    .I0_15_0_2(n89_I0_15_0_2),
    .I0_15_1_0(n89_I0_15_1_0),
    .I0_15_1_1(n89_I0_15_1_1),
    .I0_15_1_2(n89_I0_15_1_2),
    .I1_0_0(n89_I1_0_0),
    .I1_0_1(n89_I1_0_1),
    .I1_0_2(n89_I1_0_2),
    .I1_1_0(n89_I1_1_0),
    .I1_1_1(n89_I1_1_1),
    .I1_1_2(n89_I1_1_2),
    .I1_2_0(n89_I1_2_0),
    .I1_2_1(n89_I1_2_1),
    .I1_2_2(n89_I1_2_2),
    .I1_3_0(n89_I1_3_0),
    .I1_3_1(n89_I1_3_1),
    .I1_3_2(n89_I1_3_2),
    .I1_4_0(n89_I1_4_0),
    .I1_4_1(n89_I1_4_1),
    .I1_4_2(n89_I1_4_2),
    .I1_5_0(n89_I1_5_0),
    .I1_5_1(n89_I1_5_1),
    .I1_5_2(n89_I1_5_2),
    .I1_6_0(n89_I1_6_0),
    .I1_6_1(n89_I1_6_1),
    .I1_6_2(n89_I1_6_2),
    .I1_7_0(n89_I1_7_0),
    .I1_7_1(n89_I1_7_1),
    .I1_7_2(n89_I1_7_2),
    .I1_8_0(n89_I1_8_0),
    .I1_8_1(n89_I1_8_1),
    .I1_8_2(n89_I1_8_2),
    .I1_9_0(n89_I1_9_0),
    .I1_9_1(n89_I1_9_1),
    .I1_9_2(n89_I1_9_2),
    .I1_10_0(n89_I1_10_0),
    .I1_10_1(n89_I1_10_1),
    .I1_10_2(n89_I1_10_2),
    .I1_11_0(n89_I1_11_0),
    .I1_11_1(n89_I1_11_1),
    .I1_11_2(n89_I1_11_2),
    .I1_12_0(n89_I1_12_0),
    .I1_12_1(n89_I1_12_1),
    .I1_12_2(n89_I1_12_2),
    .I1_13_0(n89_I1_13_0),
    .I1_13_1(n89_I1_13_1),
    .I1_13_2(n89_I1_13_2),
    .I1_14_0(n89_I1_14_0),
    .I1_14_1(n89_I1_14_1),
    .I1_14_2(n89_I1_14_2),
    .I1_15_0(n89_I1_15_0),
    .I1_15_1(n89_I1_15_1),
    .I1_15_2(n89_I1_15_2),
    .O_0_0_0(n89_O_0_0_0),
    .O_0_0_1(n89_O_0_0_1),
    .O_0_0_2(n89_O_0_0_2),
    .O_0_1_0(n89_O_0_1_0),
    .O_0_1_1(n89_O_0_1_1),
    .O_0_1_2(n89_O_0_1_2),
    .O_0_2_0(n89_O_0_2_0),
    .O_0_2_1(n89_O_0_2_1),
    .O_0_2_2(n89_O_0_2_2),
    .O_1_0_0(n89_O_1_0_0),
    .O_1_0_1(n89_O_1_0_1),
    .O_1_0_2(n89_O_1_0_2),
    .O_1_1_0(n89_O_1_1_0),
    .O_1_1_1(n89_O_1_1_1),
    .O_1_1_2(n89_O_1_1_2),
    .O_1_2_0(n89_O_1_2_0),
    .O_1_2_1(n89_O_1_2_1),
    .O_1_2_2(n89_O_1_2_2),
    .O_2_0_0(n89_O_2_0_0),
    .O_2_0_1(n89_O_2_0_1),
    .O_2_0_2(n89_O_2_0_2),
    .O_2_1_0(n89_O_2_1_0),
    .O_2_1_1(n89_O_2_1_1),
    .O_2_1_2(n89_O_2_1_2),
    .O_2_2_0(n89_O_2_2_0),
    .O_2_2_1(n89_O_2_2_1),
    .O_2_2_2(n89_O_2_2_2),
    .O_3_0_0(n89_O_3_0_0),
    .O_3_0_1(n89_O_3_0_1),
    .O_3_0_2(n89_O_3_0_2),
    .O_3_1_0(n89_O_3_1_0),
    .O_3_1_1(n89_O_3_1_1),
    .O_3_1_2(n89_O_3_1_2),
    .O_3_2_0(n89_O_3_2_0),
    .O_3_2_1(n89_O_3_2_1),
    .O_3_2_2(n89_O_3_2_2),
    .O_4_0_0(n89_O_4_0_0),
    .O_4_0_1(n89_O_4_0_1),
    .O_4_0_2(n89_O_4_0_2),
    .O_4_1_0(n89_O_4_1_0),
    .O_4_1_1(n89_O_4_1_1),
    .O_4_1_2(n89_O_4_1_2),
    .O_4_2_0(n89_O_4_2_0),
    .O_4_2_1(n89_O_4_2_1),
    .O_4_2_2(n89_O_4_2_2),
    .O_5_0_0(n89_O_5_0_0),
    .O_5_0_1(n89_O_5_0_1),
    .O_5_0_2(n89_O_5_0_2),
    .O_5_1_0(n89_O_5_1_0),
    .O_5_1_1(n89_O_5_1_1),
    .O_5_1_2(n89_O_5_1_2),
    .O_5_2_0(n89_O_5_2_0),
    .O_5_2_1(n89_O_5_2_1),
    .O_5_2_2(n89_O_5_2_2),
    .O_6_0_0(n89_O_6_0_0),
    .O_6_0_1(n89_O_6_0_1),
    .O_6_0_2(n89_O_6_0_2),
    .O_6_1_0(n89_O_6_1_0),
    .O_6_1_1(n89_O_6_1_1),
    .O_6_1_2(n89_O_6_1_2),
    .O_6_2_0(n89_O_6_2_0),
    .O_6_2_1(n89_O_6_2_1),
    .O_6_2_2(n89_O_6_2_2),
    .O_7_0_0(n89_O_7_0_0),
    .O_7_0_1(n89_O_7_0_1),
    .O_7_0_2(n89_O_7_0_2),
    .O_7_1_0(n89_O_7_1_0),
    .O_7_1_1(n89_O_7_1_1),
    .O_7_1_2(n89_O_7_1_2),
    .O_7_2_0(n89_O_7_2_0),
    .O_7_2_1(n89_O_7_2_1),
    .O_7_2_2(n89_O_7_2_2),
    .O_8_0_0(n89_O_8_0_0),
    .O_8_0_1(n89_O_8_0_1),
    .O_8_0_2(n89_O_8_0_2),
    .O_8_1_0(n89_O_8_1_0),
    .O_8_1_1(n89_O_8_1_1),
    .O_8_1_2(n89_O_8_1_2),
    .O_8_2_0(n89_O_8_2_0),
    .O_8_2_1(n89_O_8_2_1),
    .O_8_2_2(n89_O_8_2_2),
    .O_9_0_0(n89_O_9_0_0),
    .O_9_0_1(n89_O_9_0_1),
    .O_9_0_2(n89_O_9_0_2),
    .O_9_1_0(n89_O_9_1_0),
    .O_9_1_1(n89_O_9_1_1),
    .O_9_1_2(n89_O_9_1_2),
    .O_9_2_0(n89_O_9_2_0),
    .O_9_2_1(n89_O_9_2_1),
    .O_9_2_2(n89_O_9_2_2),
    .O_10_0_0(n89_O_10_0_0),
    .O_10_0_1(n89_O_10_0_1),
    .O_10_0_2(n89_O_10_0_2),
    .O_10_1_0(n89_O_10_1_0),
    .O_10_1_1(n89_O_10_1_1),
    .O_10_1_2(n89_O_10_1_2),
    .O_10_2_0(n89_O_10_2_0),
    .O_10_2_1(n89_O_10_2_1),
    .O_10_2_2(n89_O_10_2_2),
    .O_11_0_0(n89_O_11_0_0),
    .O_11_0_1(n89_O_11_0_1),
    .O_11_0_2(n89_O_11_0_2),
    .O_11_1_0(n89_O_11_1_0),
    .O_11_1_1(n89_O_11_1_1),
    .O_11_1_2(n89_O_11_1_2),
    .O_11_2_0(n89_O_11_2_0),
    .O_11_2_1(n89_O_11_2_1),
    .O_11_2_2(n89_O_11_2_2),
    .O_12_0_0(n89_O_12_0_0),
    .O_12_0_1(n89_O_12_0_1),
    .O_12_0_2(n89_O_12_0_2),
    .O_12_1_0(n89_O_12_1_0),
    .O_12_1_1(n89_O_12_1_1),
    .O_12_1_2(n89_O_12_1_2),
    .O_12_2_0(n89_O_12_2_0),
    .O_12_2_1(n89_O_12_2_1),
    .O_12_2_2(n89_O_12_2_2),
    .O_13_0_0(n89_O_13_0_0),
    .O_13_0_1(n89_O_13_0_1),
    .O_13_0_2(n89_O_13_0_2),
    .O_13_1_0(n89_O_13_1_0),
    .O_13_1_1(n89_O_13_1_1),
    .O_13_1_2(n89_O_13_1_2),
    .O_13_2_0(n89_O_13_2_0),
    .O_13_2_1(n89_O_13_2_1),
    .O_13_2_2(n89_O_13_2_2),
    .O_14_0_0(n89_O_14_0_0),
    .O_14_0_1(n89_O_14_0_1),
    .O_14_0_2(n89_O_14_0_2),
    .O_14_1_0(n89_O_14_1_0),
    .O_14_1_1(n89_O_14_1_1),
    .O_14_1_2(n89_O_14_1_2),
    .O_14_2_0(n89_O_14_2_0),
    .O_14_2_1(n89_O_14_2_1),
    .O_14_2_2(n89_O_14_2_2),
    .O_15_0_0(n89_O_15_0_0),
    .O_15_0_1(n89_O_15_0_1),
    .O_15_0_2(n89_O_15_0_2),
    .O_15_1_0(n89_O_15_1_0),
    .O_15_1_1(n89_O_15_1_1),
    .O_15_1_2(n89_O_15_1_2),
    .O_15_2_0(n89_O_15_2_0),
    .O_15_2_1(n89_O_15_2_1),
    .O_15_2_2(n89_O_15_2_2)
  );
  MapT_6 n98 ( // @[Top.scala 151:21]
    .valid_up(n98_valid_up),
    .valid_down(n98_valid_down),
    .I_0_0_0(n98_I_0_0_0),
    .I_0_0_1(n98_I_0_0_1),
    .I_0_0_2(n98_I_0_0_2),
    .I_0_1_0(n98_I_0_1_0),
    .I_0_1_1(n98_I_0_1_1),
    .I_0_1_2(n98_I_0_1_2),
    .I_0_2_0(n98_I_0_2_0),
    .I_0_2_1(n98_I_0_2_1),
    .I_0_2_2(n98_I_0_2_2),
    .I_1_0_0(n98_I_1_0_0),
    .I_1_0_1(n98_I_1_0_1),
    .I_1_0_2(n98_I_1_0_2),
    .I_1_1_0(n98_I_1_1_0),
    .I_1_1_1(n98_I_1_1_1),
    .I_1_1_2(n98_I_1_1_2),
    .I_1_2_0(n98_I_1_2_0),
    .I_1_2_1(n98_I_1_2_1),
    .I_1_2_2(n98_I_1_2_2),
    .I_2_0_0(n98_I_2_0_0),
    .I_2_0_1(n98_I_2_0_1),
    .I_2_0_2(n98_I_2_0_2),
    .I_2_1_0(n98_I_2_1_0),
    .I_2_1_1(n98_I_2_1_1),
    .I_2_1_2(n98_I_2_1_2),
    .I_2_2_0(n98_I_2_2_0),
    .I_2_2_1(n98_I_2_2_1),
    .I_2_2_2(n98_I_2_2_2),
    .I_3_0_0(n98_I_3_0_0),
    .I_3_0_1(n98_I_3_0_1),
    .I_3_0_2(n98_I_3_0_2),
    .I_3_1_0(n98_I_3_1_0),
    .I_3_1_1(n98_I_3_1_1),
    .I_3_1_2(n98_I_3_1_2),
    .I_3_2_0(n98_I_3_2_0),
    .I_3_2_1(n98_I_3_2_1),
    .I_3_2_2(n98_I_3_2_2),
    .I_4_0_0(n98_I_4_0_0),
    .I_4_0_1(n98_I_4_0_1),
    .I_4_0_2(n98_I_4_0_2),
    .I_4_1_0(n98_I_4_1_0),
    .I_4_1_1(n98_I_4_1_1),
    .I_4_1_2(n98_I_4_1_2),
    .I_4_2_0(n98_I_4_2_0),
    .I_4_2_1(n98_I_4_2_1),
    .I_4_2_2(n98_I_4_2_2),
    .I_5_0_0(n98_I_5_0_0),
    .I_5_0_1(n98_I_5_0_1),
    .I_5_0_2(n98_I_5_0_2),
    .I_5_1_0(n98_I_5_1_0),
    .I_5_1_1(n98_I_5_1_1),
    .I_5_1_2(n98_I_5_1_2),
    .I_5_2_0(n98_I_5_2_0),
    .I_5_2_1(n98_I_5_2_1),
    .I_5_2_2(n98_I_5_2_2),
    .I_6_0_0(n98_I_6_0_0),
    .I_6_0_1(n98_I_6_0_1),
    .I_6_0_2(n98_I_6_0_2),
    .I_6_1_0(n98_I_6_1_0),
    .I_6_1_1(n98_I_6_1_1),
    .I_6_1_2(n98_I_6_1_2),
    .I_6_2_0(n98_I_6_2_0),
    .I_6_2_1(n98_I_6_2_1),
    .I_6_2_2(n98_I_6_2_2),
    .I_7_0_0(n98_I_7_0_0),
    .I_7_0_1(n98_I_7_0_1),
    .I_7_0_2(n98_I_7_0_2),
    .I_7_1_0(n98_I_7_1_0),
    .I_7_1_1(n98_I_7_1_1),
    .I_7_1_2(n98_I_7_1_2),
    .I_7_2_0(n98_I_7_2_0),
    .I_7_2_1(n98_I_7_2_1),
    .I_7_2_2(n98_I_7_2_2),
    .I_8_0_0(n98_I_8_0_0),
    .I_8_0_1(n98_I_8_0_1),
    .I_8_0_2(n98_I_8_0_2),
    .I_8_1_0(n98_I_8_1_0),
    .I_8_1_1(n98_I_8_1_1),
    .I_8_1_2(n98_I_8_1_2),
    .I_8_2_0(n98_I_8_2_0),
    .I_8_2_1(n98_I_8_2_1),
    .I_8_2_2(n98_I_8_2_2),
    .I_9_0_0(n98_I_9_0_0),
    .I_9_0_1(n98_I_9_0_1),
    .I_9_0_2(n98_I_9_0_2),
    .I_9_1_0(n98_I_9_1_0),
    .I_9_1_1(n98_I_9_1_1),
    .I_9_1_2(n98_I_9_1_2),
    .I_9_2_0(n98_I_9_2_0),
    .I_9_2_1(n98_I_9_2_1),
    .I_9_2_2(n98_I_9_2_2),
    .I_10_0_0(n98_I_10_0_0),
    .I_10_0_1(n98_I_10_0_1),
    .I_10_0_2(n98_I_10_0_2),
    .I_10_1_0(n98_I_10_1_0),
    .I_10_1_1(n98_I_10_1_1),
    .I_10_1_2(n98_I_10_1_2),
    .I_10_2_0(n98_I_10_2_0),
    .I_10_2_1(n98_I_10_2_1),
    .I_10_2_2(n98_I_10_2_2),
    .I_11_0_0(n98_I_11_0_0),
    .I_11_0_1(n98_I_11_0_1),
    .I_11_0_2(n98_I_11_0_2),
    .I_11_1_0(n98_I_11_1_0),
    .I_11_1_1(n98_I_11_1_1),
    .I_11_1_2(n98_I_11_1_2),
    .I_11_2_0(n98_I_11_2_0),
    .I_11_2_1(n98_I_11_2_1),
    .I_11_2_2(n98_I_11_2_2),
    .I_12_0_0(n98_I_12_0_0),
    .I_12_0_1(n98_I_12_0_1),
    .I_12_0_2(n98_I_12_0_2),
    .I_12_1_0(n98_I_12_1_0),
    .I_12_1_1(n98_I_12_1_1),
    .I_12_1_2(n98_I_12_1_2),
    .I_12_2_0(n98_I_12_2_0),
    .I_12_2_1(n98_I_12_2_1),
    .I_12_2_2(n98_I_12_2_2),
    .I_13_0_0(n98_I_13_0_0),
    .I_13_0_1(n98_I_13_0_1),
    .I_13_0_2(n98_I_13_0_2),
    .I_13_1_0(n98_I_13_1_0),
    .I_13_1_1(n98_I_13_1_1),
    .I_13_1_2(n98_I_13_1_2),
    .I_13_2_0(n98_I_13_2_0),
    .I_13_2_1(n98_I_13_2_1),
    .I_13_2_2(n98_I_13_2_2),
    .I_14_0_0(n98_I_14_0_0),
    .I_14_0_1(n98_I_14_0_1),
    .I_14_0_2(n98_I_14_0_2),
    .I_14_1_0(n98_I_14_1_0),
    .I_14_1_1(n98_I_14_1_1),
    .I_14_1_2(n98_I_14_1_2),
    .I_14_2_0(n98_I_14_2_0),
    .I_14_2_1(n98_I_14_2_1),
    .I_14_2_2(n98_I_14_2_2),
    .I_15_0_0(n98_I_15_0_0),
    .I_15_0_1(n98_I_15_0_1),
    .I_15_0_2(n98_I_15_0_2),
    .I_15_1_0(n98_I_15_1_0),
    .I_15_1_1(n98_I_15_1_1),
    .I_15_1_2(n98_I_15_1_2),
    .I_15_2_0(n98_I_15_2_0),
    .I_15_2_1(n98_I_15_2_1),
    .I_15_2_2(n98_I_15_2_2),
    .O_0_0_0_0(n98_O_0_0_0_0),
    .O_0_0_0_1(n98_O_0_0_0_1),
    .O_0_0_0_2(n98_O_0_0_0_2),
    .O_0_0_1_0(n98_O_0_0_1_0),
    .O_0_0_1_1(n98_O_0_0_1_1),
    .O_0_0_1_2(n98_O_0_0_1_2),
    .O_0_0_2_0(n98_O_0_0_2_0),
    .O_0_0_2_1(n98_O_0_0_2_1),
    .O_0_0_2_2(n98_O_0_0_2_2),
    .O_1_0_0_0(n98_O_1_0_0_0),
    .O_1_0_0_1(n98_O_1_0_0_1),
    .O_1_0_0_2(n98_O_1_0_0_2),
    .O_1_0_1_0(n98_O_1_0_1_0),
    .O_1_0_1_1(n98_O_1_0_1_1),
    .O_1_0_1_2(n98_O_1_0_1_2),
    .O_1_0_2_0(n98_O_1_0_2_0),
    .O_1_0_2_1(n98_O_1_0_2_1),
    .O_1_0_2_2(n98_O_1_0_2_2),
    .O_2_0_0_0(n98_O_2_0_0_0),
    .O_2_0_0_1(n98_O_2_0_0_1),
    .O_2_0_0_2(n98_O_2_0_0_2),
    .O_2_0_1_0(n98_O_2_0_1_0),
    .O_2_0_1_1(n98_O_2_0_1_1),
    .O_2_0_1_2(n98_O_2_0_1_2),
    .O_2_0_2_0(n98_O_2_0_2_0),
    .O_2_0_2_1(n98_O_2_0_2_1),
    .O_2_0_2_2(n98_O_2_0_2_2),
    .O_3_0_0_0(n98_O_3_0_0_0),
    .O_3_0_0_1(n98_O_3_0_0_1),
    .O_3_0_0_2(n98_O_3_0_0_2),
    .O_3_0_1_0(n98_O_3_0_1_0),
    .O_3_0_1_1(n98_O_3_0_1_1),
    .O_3_0_1_2(n98_O_3_0_1_2),
    .O_3_0_2_0(n98_O_3_0_2_0),
    .O_3_0_2_1(n98_O_3_0_2_1),
    .O_3_0_2_2(n98_O_3_0_2_2),
    .O_4_0_0_0(n98_O_4_0_0_0),
    .O_4_0_0_1(n98_O_4_0_0_1),
    .O_4_0_0_2(n98_O_4_0_0_2),
    .O_4_0_1_0(n98_O_4_0_1_0),
    .O_4_0_1_1(n98_O_4_0_1_1),
    .O_4_0_1_2(n98_O_4_0_1_2),
    .O_4_0_2_0(n98_O_4_0_2_0),
    .O_4_0_2_1(n98_O_4_0_2_1),
    .O_4_0_2_2(n98_O_4_0_2_2),
    .O_5_0_0_0(n98_O_5_0_0_0),
    .O_5_0_0_1(n98_O_5_0_0_1),
    .O_5_0_0_2(n98_O_5_0_0_2),
    .O_5_0_1_0(n98_O_5_0_1_0),
    .O_5_0_1_1(n98_O_5_0_1_1),
    .O_5_0_1_2(n98_O_5_0_1_2),
    .O_5_0_2_0(n98_O_5_0_2_0),
    .O_5_0_2_1(n98_O_5_0_2_1),
    .O_5_0_2_2(n98_O_5_0_2_2),
    .O_6_0_0_0(n98_O_6_0_0_0),
    .O_6_0_0_1(n98_O_6_0_0_1),
    .O_6_0_0_2(n98_O_6_0_0_2),
    .O_6_0_1_0(n98_O_6_0_1_0),
    .O_6_0_1_1(n98_O_6_0_1_1),
    .O_6_0_1_2(n98_O_6_0_1_2),
    .O_6_0_2_0(n98_O_6_0_2_0),
    .O_6_0_2_1(n98_O_6_0_2_1),
    .O_6_0_2_2(n98_O_6_0_2_2),
    .O_7_0_0_0(n98_O_7_0_0_0),
    .O_7_0_0_1(n98_O_7_0_0_1),
    .O_7_0_0_2(n98_O_7_0_0_2),
    .O_7_0_1_0(n98_O_7_0_1_0),
    .O_7_0_1_1(n98_O_7_0_1_1),
    .O_7_0_1_2(n98_O_7_0_1_2),
    .O_7_0_2_0(n98_O_7_0_2_0),
    .O_7_0_2_1(n98_O_7_0_2_1),
    .O_7_0_2_2(n98_O_7_0_2_2),
    .O_8_0_0_0(n98_O_8_0_0_0),
    .O_8_0_0_1(n98_O_8_0_0_1),
    .O_8_0_0_2(n98_O_8_0_0_2),
    .O_8_0_1_0(n98_O_8_0_1_0),
    .O_8_0_1_1(n98_O_8_0_1_1),
    .O_8_0_1_2(n98_O_8_0_1_2),
    .O_8_0_2_0(n98_O_8_0_2_0),
    .O_8_0_2_1(n98_O_8_0_2_1),
    .O_8_0_2_2(n98_O_8_0_2_2),
    .O_9_0_0_0(n98_O_9_0_0_0),
    .O_9_0_0_1(n98_O_9_0_0_1),
    .O_9_0_0_2(n98_O_9_0_0_2),
    .O_9_0_1_0(n98_O_9_0_1_0),
    .O_9_0_1_1(n98_O_9_0_1_1),
    .O_9_0_1_2(n98_O_9_0_1_2),
    .O_9_0_2_0(n98_O_9_0_2_0),
    .O_9_0_2_1(n98_O_9_0_2_1),
    .O_9_0_2_2(n98_O_9_0_2_2),
    .O_10_0_0_0(n98_O_10_0_0_0),
    .O_10_0_0_1(n98_O_10_0_0_1),
    .O_10_0_0_2(n98_O_10_0_0_2),
    .O_10_0_1_0(n98_O_10_0_1_0),
    .O_10_0_1_1(n98_O_10_0_1_1),
    .O_10_0_1_2(n98_O_10_0_1_2),
    .O_10_0_2_0(n98_O_10_0_2_0),
    .O_10_0_2_1(n98_O_10_0_2_1),
    .O_10_0_2_2(n98_O_10_0_2_2),
    .O_11_0_0_0(n98_O_11_0_0_0),
    .O_11_0_0_1(n98_O_11_0_0_1),
    .O_11_0_0_2(n98_O_11_0_0_2),
    .O_11_0_1_0(n98_O_11_0_1_0),
    .O_11_0_1_1(n98_O_11_0_1_1),
    .O_11_0_1_2(n98_O_11_0_1_2),
    .O_11_0_2_0(n98_O_11_0_2_0),
    .O_11_0_2_1(n98_O_11_0_2_1),
    .O_11_0_2_2(n98_O_11_0_2_2),
    .O_12_0_0_0(n98_O_12_0_0_0),
    .O_12_0_0_1(n98_O_12_0_0_1),
    .O_12_0_0_2(n98_O_12_0_0_2),
    .O_12_0_1_0(n98_O_12_0_1_0),
    .O_12_0_1_1(n98_O_12_0_1_1),
    .O_12_0_1_2(n98_O_12_0_1_2),
    .O_12_0_2_0(n98_O_12_0_2_0),
    .O_12_0_2_1(n98_O_12_0_2_1),
    .O_12_0_2_2(n98_O_12_0_2_2),
    .O_13_0_0_0(n98_O_13_0_0_0),
    .O_13_0_0_1(n98_O_13_0_0_1),
    .O_13_0_0_2(n98_O_13_0_0_2),
    .O_13_0_1_0(n98_O_13_0_1_0),
    .O_13_0_1_1(n98_O_13_0_1_1),
    .O_13_0_1_2(n98_O_13_0_1_2),
    .O_13_0_2_0(n98_O_13_0_2_0),
    .O_13_0_2_1(n98_O_13_0_2_1),
    .O_13_0_2_2(n98_O_13_0_2_2),
    .O_14_0_0_0(n98_O_14_0_0_0),
    .O_14_0_0_1(n98_O_14_0_0_1),
    .O_14_0_0_2(n98_O_14_0_0_2),
    .O_14_0_1_0(n98_O_14_0_1_0),
    .O_14_0_1_1(n98_O_14_0_1_1),
    .O_14_0_1_2(n98_O_14_0_1_2),
    .O_14_0_2_0(n98_O_14_0_2_0),
    .O_14_0_2_1(n98_O_14_0_2_1),
    .O_14_0_2_2(n98_O_14_0_2_2),
    .O_15_0_0_0(n98_O_15_0_0_0),
    .O_15_0_0_1(n98_O_15_0_0_1),
    .O_15_0_0_2(n98_O_15_0_0_2),
    .O_15_0_1_0(n98_O_15_0_1_0),
    .O_15_0_1_1(n98_O_15_0_1_1),
    .O_15_0_1_2(n98_O_15_0_1_2),
    .O_15_0_2_0(n98_O_15_0_2_0),
    .O_15_0_2_1(n98_O_15_0_2_1),
    .O_15_0_2_2(n98_O_15_0_2_2)
  );
  MapT_7 n105 ( // @[Top.scala 154:22]
    .valid_up(n105_valid_up),
    .valid_down(n105_valid_down),
    .I_0_0_0_0(n105_I_0_0_0_0),
    .I_0_0_0_1(n105_I_0_0_0_1),
    .I_0_0_0_2(n105_I_0_0_0_2),
    .I_0_0_1_0(n105_I_0_0_1_0),
    .I_0_0_1_1(n105_I_0_0_1_1),
    .I_0_0_1_2(n105_I_0_0_1_2),
    .I_0_0_2_0(n105_I_0_0_2_0),
    .I_0_0_2_1(n105_I_0_0_2_1),
    .I_0_0_2_2(n105_I_0_0_2_2),
    .I_1_0_0_0(n105_I_1_0_0_0),
    .I_1_0_0_1(n105_I_1_0_0_1),
    .I_1_0_0_2(n105_I_1_0_0_2),
    .I_1_0_1_0(n105_I_1_0_1_0),
    .I_1_0_1_1(n105_I_1_0_1_1),
    .I_1_0_1_2(n105_I_1_0_1_2),
    .I_1_0_2_0(n105_I_1_0_2_0),
    .I_1_0_2_1(n105_I_1_0_2_1),
    .I_1_0_2_2(n105_I_1_0_2_2),
    .I_2_0_0_0(n105_I_2_0_0_0),
    .I_2_0_0_1(n105_I_2_0_0_1),
    .I_2_0_0_2(n105_I_2_0_0_2),
    .I_2_0_1_0(n105_I_2_0_1_0),
    .I_2_0_1_1(n105_I_2_0_1_1),
    .I_2_0_1_2(n105_I_2_0_1_2),
    .I_2_0_2_0(n105_I_2_0_2_0),
    .I_2_0_2_1(n105_I_2_0_2_1),
    .I_2_0_2_2(n105_I_2_0_2_2),
    .I_3_0_0_0(n105_I_3_0_0_0),
    .I_3_0_0_1(n105_I_3_0_0_1),
    .I_3_0_0_2(n105_I_3_0_0_2),
    .I_3_0_1_0(n105_I_3_0_1_0),
    .I_3_0_1_1(n105_I_3_0_1_1),
    .I_3_0_1_2(n105_I_3_0_1_2),
    .I_3_0_2_0(n105_I_3_0_2_0),
    .I_3_0_2_1(n105_I_3_0_2_1),
    .I_3_0_2_2(n105_I_3_0_2_2),
    .I_4_0_0_0(n105_I_4_0_0_0),
    .I_4_0_0_1(n105_I_4_0_0_1),
    .I_4_0_0_2(n105_I_4_0_0_2),
    .I_4_0_1_0(n105_I_4_0_1_0),
    .I_4_0_1_1(n105_I_4_0_1_1),
    .I_4_0_1_2(n105_I_4_0_1_2),
    .I_4_0_2_0(n105_I_4_0_2_0),
    .I_4_0_2_1(n105_I_4_0_2_1),
    .I_4_0_2_2(n105_I_4_0_2_2),
    .I_5_0_0_0(n105_I_5_0_0_0),
    .I_5_0_0_1(n105_I_5_0_0_1),
    .I_5_0_0_2(n105_I_5_0_0_2),
    .I_5_0_1_0(n105_I_5_0_1_0),
    .I_5_0_1_1(n105_I_5_0_1_1),
    .I_5_0_1_2(n105_I_5_0_1_2),
    .I_5_0_2_0(n105_I_5_0_2_0),
    .I_5_0_2_1(n105_I_5_0_2_1),
    .I_5_0_2_2(n105_I_5_0_2_2),
    .I_6_0_0_0(n105_I_6_0_0_0),
    .I_6_0_0_1(n105_I_6_0_0_1),
    .I_6_0_0_2(n105_I_6_0_0_2),
    .I_6_0_1_0(n105_I_6_0_1_0),
    .I_6_0_1_1(n105_I_6_0_1_1),
    .I_6_0_1_2(n105_I_6_0_1_2),
    .I_6_0_2_0(n105_I_6_0_2_0),
    .I_6_0_2_1(n105_I_6_0_2_1),
    .I_6_0_2_2(n105_I_6_0_2_2),
    .I_7_0_0_0(n105_I_7_0_0_0),
    .I_7_0_0_1(n105_I_7_0_0_1),
    .I_7_0_0_2(n105_I_7_0_0_2),
    .I_7_0_1_0(n105_I_7_0_1_0),
    .I_7_0_1_1(n105_I_7_0_1_1),
    .I_7_0_1_2(n105_I_7_0_1_2),
    .I_7_0_2_0(n105_I_7_0_2_0),
    .I_7_0_2_1(n105_I_7_0_2_1),
    .I_7_0_2_2(n105_I_7_0_2_2),
    .I_8_0_0_0(n105_I_8_0_0_0),
    .I_8_0_0_1(n105_I_8_0_0_1),
    .I_8_0_0_2(n105_I_8_0_0_2),
    .I_8_0_1_0(n105_I_8_0_1_0),
    .I_8_0_1_1(n105_I_8_0_1_1),
    .I_8_0_1_2(n105_I_8_0_1_2),
    .I_8_0_2_0(n105_I_8_0_2_0),
    .I_8_0_2_1(n105_I_8_0_2_1),
    .I_8_0_2_2(n105_I_8_0_2_2),
    .I_9_0_0_0(n105_I_9_0_0_0),
    .I_9_0_0_1(n105_I_9_0_0_1),
    .I_9_0_0_2(n105_I_9_0_0_2),
    .I_9_0_1_0(n105_I_9_0_1_0),
    .I_9_0_1_1(n105_I_9_0_1_1),
    .I_9_0_1_2(n105_I_9_0_1_2),
    .I_9_0_2_0(n105_I_9_0_2_0),
    .I_9_0_2_1(n105_I_9_0_2_1),
    .I_9_0_2_2(n105_I_9_0_2_2),
    .I_10_0_0_0(n105_I_10_0_0_0),
    .I_10_0_0_1(n105_I_10_0_0_1),
    .I_10_0_0_2(n105_I_10_0_0_2),
    .I_10_0_1_0(n105_I_10_0_1_0),
    .I_10_0_1_1(n105_I_10_0_1_1),
    .I_10_0_1_2(n105_I_10_0_1_2),
    .I_10_0_2_0(n105_I_10_0_2_0),
    .I_10_0_2_1(n105_I_10_0_2_1),
    .I_10_0_2_2(n105_I_10_0_2_2),
    .I_11_0_0_0(n105_I_11_0_0_0),
    .I_11_0_0_1(n105_I_11_0_0_1),
    .I_11_0_0_2(n105_I_11_0_0_2),
    .I_11_0_1_0(n105_I_11_0_1_0),
    .I_11_0_1_1(n105_I_11_0_1_1),
    .I_11_0_1_2(n105_I_11_0_1_2),
    .I_11_0_2_0(n105_I_11_0_2_0),
    .I_11_0_2_1(n105_I_11_0_2_1),
    .I_11_0_2_2(n105_I_11_0_2_2),
    .I_12_0_0_0(n105_I_12_0_0_0),
    .I_12_0_0_1(n105_I_12_0_0_1),
    .I_12_0_0_2(n105_I_12_0_0_2),
    .I_12_0_1_0(n105_I_12_0_1_0),
    .I_12_0_1_1(n105_I_12_0_1_1),
    .I_12_0_1_2(n105_I_12_0_1_2),
    .I_12_0_2_0(n105_I_12_0_2_0),
    .I_12_0_2_1(n105_I_12_0_2_1),
    .I_12_0_2_2(n105_I_12_0_2_2),
    .I_13_0_0_0(n105_I_13_0_0_0),
    .I_13_0_0_1(n105_I_13_0_0_1),
    .I_13_0_0_2(n105_I_13_0_0_2),
    .I_13_0_1_0(n105_I_13_0_1_0),
    .I_13_0_1_1(n105_I_13_0_1_1),
    .I_13_0_1_2(n105_I_13_0_1_2),
    .I_13_0_2_0(n105_I_13_0_2_0),
    .I_13_0_2_1(n105_I_13_0_2_1),
    .I_13_0_2_2(n105_I_13_0_2_2),
    .I_14_0_0_0(n105_I_14_0_0_0),
    .I_14_0_0_1(n105_I_14_0_0_1),
    .I_14_0_0_2(n105_I_14_0_0_2),
    .I_14_0_1_0(n105_I_14_0_1_0),
    .I_14_0_1_1(n105_I_14_0_1_1),
    .I_14_0_1_2(n105_I_14_0_1_2),
    .I_14_0_2_0(n105_I_14_0_2_0),
    .I_14_0_2_1(n105_I_14_0_2_1),
    .I_14_0_2_2(n105_I_14_0_2_2),
    .I_15_0_0_0(n105_I_15_0_0_0),
    .I_15_0_0_1(n105_I_15_0_0_1),
    .I_15_0_0_2(n105_I_15_0_0_2),
    .I_15_0_1_0(n105_I_15_0_1_0),
    .I_15_0_1_1(n105_I_15_0_1_1),
    .I_15_0_1_2(n105_I_15_0_1_2),
    .I_15_0_2_0(n105_I_15_0_2_0),
    .I_15_0_2_1(n105_I_15_0_2_1),
    .I_15_0_2_2(n105_I_15_0_2_2),
    .O_0_0_0(n105_O_0_0_0),
    .O_0_0_1(n105_O_0_0_1),
    .O_0_0_2(n105_O_0_0_2),
    .O_0_1_0(n105_O_0_1_0),
    .O_0_1_1(n105_O_0_1_1),
    .O_0_1_2(n105_O_0_1_2),
    .O_0_2_0(n105_O_0_2_0),
    .O_0_2_1(n105_O_0_2_1),
    .O_0_2_2(n105_O_0_2_2),
    .O_1_0_0(n105_O_1_0_0),
    .O_1_0_1(n105_O_1_0_1),
    .O_1_0_2(n105_O_1_0_2),
    .O_1_1_0(n105_O_1_1_0),
    .O_1_1_1(n105_O_1_1_1),
    .O_1_1_2(n105_O_1_1_2),
    .O_1_2_0(n105_O_1_2_0),
    .O_1_2_1(n105_O_1_2_1),
    .O_1_2_2(n105_O_1_2_2),
    .O_2_0_0(n105_O_2_0_0),
    .O_2_0_1(n105_O_2_0_1),
    .O_2_0_2(n105_O_2_0_2),
    .O_2_1_0(n105_O_2_1_0),
    .O_2_1_1(n105_O_2_1_1),
    .O_2_1_2(n105_O_2_1_2),
    .O_2_2_0(n105_O_2_2_0),
    .O_2_2_1(n105_O_2_2_1),
    .O_2_2_2(n105_O_2_2_2),
    .O_3_0_0(n105_O_3_0_0),
    .O_3_0_1(n105_O_3_0_1),
    .O_3_0_2(n105_O_3_0_2),
    .O_3_1_0(n105_O_3_1_0),
    .O_3_1_1(n105_O_3_1_1),
    .O_3_1_2(n105_O_3_1_2),
    .O_3_2_0(n105_O_3_2_0),
    .O_3_2_1(n105_O_3_2_1),
    .O_3_2_2(n105_O_3_2_2),
    .O_4_0_0(n105_O_4_0_0),
    .O_4_0_1(n105_O_4_0_1),
    .O_4_0_2(n105_O_4_0_2),
    .O_4_1_0(n105_O_4_1_0),
    .O_4_1_1(n105_O_4_1_1),
    .O_4_1_2(n105_O_4_1_2),
    .O_4_2_0(n105_O_4_2_0),
    .O_4_2_1(n105_O_4_2_1),
    .O_4_2_2(n105_O_4_2_2),
    .O_5_0_0(n105_O_5_0_0),
    .O_5_0_1(n105_O_5_0_1),
    .O_5_0_2(n105_O_5_0_2),
    .O_5_1_0(n105_O_5_1_0),
    .O_5_1_1(n105_O_5_1_1),
    .O_5_1_2(n105_O_5_1_2),
    .O_5_2_0(n105_O_5_2_0),
    .O_5_2_1(n105_O_5_2_1),
    .O_5_2_2(n105_O_5_2_2),
    .O_6_0_0(n105_O_6_0_0),
    .O_6_0_1(n105_O_6_0_1),
    .O_6_0_2(n105_O_6_0_2),
    .O_6_1_0(n105_O_6_1_0),
    .O_6_1_1(n105_O_6_1_1),
    .O_6_1_2(n105_O_6_1_2),
    .O_6_2_0(n105_O_6_2_0),
    .O_6_2_1(n105_O_6_2_1),
    .O_6_2_2(n105_O_6_2_2),
    .O_7_0_0(n105_O_7_0_0),
    .O_7_0_1(n105_O_7_0_1),
    .O_7_0_2(n105_O_7_0_2),
    .O_7_1_0(n105_O_7_1_0),
    .O_7_1_1(n105_O_7_1_1),
    .O_7_1_2(n105_O_7_1_2),
    .O_7_2_0(n105_O_7_2_0),
    .O_7_2_1(n105_O_7_2_1),
    .O_7_2_2(n105_O_7_2_2),
    .O_8_0_0(n105_O_8_0_0),
    .O_8_0_1(n105_O_8_0_1),
    .O_8_0_2(n105_O_8_0_2),
    .O_8_1_0(n105_O_8_1_0),
    .O_8_1_1(n105_O_8_1_1),
    .O_8_1_2(n105_O_8_1_2),
    .O_8_2_0(n105_O_8_2_0),
    .O_8_2_1(n105_O_8_2_1),
    .O_8_2_2(n105_O_8_2_2),
    .O_9_0_0(n105_O_9_0_0),
    .O_9_0_1(n105_O_9_0_1),
    .O_9_0_2(n105_O_9_0_2),
    .O_9_1_0(n105_O_9_1_0),
    .O_9_1_1(n105_O_9_1_1),
    .O_9_1_2(n105_O_9_1_2),
    .O_9_2_0(n105_O_9_2_0),
    .O_9_2_1(n105_O_9_2_1),
    .O_9_2_2(n105_O_9_2_2),
    .O_10_0_0(n105_O_10_0_0),
    .O_10_0_1(n105_O_10_0_1),
    .O_10_0_2(n105_O_10_0_2),
    .O_10_1_0(n105_O_10_1_0),
    .O_10_1_1(n105_O_10_1_1),
    .O_10_1_2(n105_O_10_1_2),
    .O_10_2_0(n105_O_10_2_0),
    .O_10_2_1(n105_O_10_2_1),
    .O_10_2_2(n105_O_10_2_2),
    .O_11_0_0(n105_O_11_0_0),
    .O_11_0_1(n105_O_11_0_1),
    .O_11_0_2(n105_O_11_0_2),
    .O_11_1_0(n105_O_11_1_0),
    .O_11_1_1(n105_O_11_1_1),
    .O_11_1_2(n105_O_11_1_2),
    .O_11_2_0(n105_O_11_2_0),
    .O_11_2_1(n105_O_11_2_1),
    .O_11_2_2(n105_O_11_2_2),
    .O_12_0_0(n105_O_12_0_0),
    .O_12_0_1(n105_O_12_0_1),
    .O_12_0_2(n105_O_12_0_2),
    .O_12_1_0(n105_O_12_1_0),
    .O_12_1_1(n105_O_12_1_1),
    .O_12_1_2(n105_O_12_1_2),
    .O_12_2_0(n105_O_12_2_0),
    .O_12_2_1(n105_O_12_2_1),
    .O_12_2_2(n105_O_12_2_2),
    .O_13_0_0(n105_O_13_0_0),
    .O_13_0_1(n105_O_13_0_1),
    .O_13_0_2(n105_O_13_0_2),
    .O_13_1_0(n105_O_13_1_0),
    .O_13_1_1(n105_O_13_1_1),
    .O_13_1_2(n105_O_13_1_2),
    .O_13_2_0(n105_O_13_2_0),
    .O_13_2_1(n105_O_13_2_1),
    .O_13_2_2(n105_O_13_2_2),
    .O_14_0_0(n105_O_14_0_0),
    .O_14_0_1(n105_O_14_0_1),
    .O_14_0_2(n105_O_14_0_2),
    .O_14_1_0(n105_O_14_1_0),
    .O_14_1_1(n105_O_14_1_1),
    .O_14_1_2(n105_O_14_1_2),
    .O_14_2_0(n105_O_14_2_0),
    .O_14_2_1(n105_O_14_2_1),
    .O_14_2_2(n105_O_14_2_2),
    .O_15_0_0(n105_O_15_0_0),
    .O_15_0_1(n105_O_15_0_1),
    .O_15_0_2(n105_O_15_0_2),
    .O_15_1_0(n105_O_15_1_0),
    .O_15_1_1(n105_O_15_1_1),
    .O_15_1_2(n105_O_15_1_2),
    .O_15_2_0(n105_O_15_2_0),
    .O_15_2_1(n105_O_15_2_1),
    .O_15_2_2(n105_O_15_2_2)
  );
  MapT_8 n147 ( // @[Top.scala 157:22]
    .clock(n147_clock),
    .reset(n147_reset),
    .valid_up(n147_valid_up),
    .valid_down(n147_valid_down),
    .I_0_0_0(n147_I_0_0_0),
    .I_0_0_1(n147_I_0_0_1),
    .I_0_0_2(n147_I_0_0_2),
    .I_0_1_0(n147_I_0_1_0),
    .I_0_1_1(n147_I_0_1_1),
    .I_0_1_2(n147_I_0_1_2),
    .I_0_2_0(n147_I_0_2_0),
    .I_0_2_1(n147_I_0_2_1),
    .I_0_2_2(n147_I_0_2_2),
    .I_1_0_0(n147_I_1_0_0),
    .I_1_0_1(n147_I_1_0_1),
    .I_1_0_2(n147_I_1_0_2),
    .I_1_1_0(n147_I_1_1_0),
    .I_1_1_1(n147_I_1_1_1),
    .I_1_1_2(n147_I_1_1_2),
    .I_1_2_0(n147_I_1_2_0),
    .I_1_2_1(n147_I_1_2_1),
    .I_1_2_2(n147_I_1_2_2),
    .I_2_0_0(n147_I_2_0_0),
    .I_2_0_1(n147_I_2_0_1),
    .I_2_0_2(n147_I_2_0_2),
    .I_2_1_0(n147_I_2_1_0),
    .I_2_1_1(n147_I_2_1_1),
    .I_2_1_2(n147_I_2_1_2),
    .I_2_2_0(n147_I_2_2_0),
    .I_2_2_1(n147_I_2_2_1),
    .I_2_2_2(n147_I_2_2_2),
    .I_3_0_0(n147_I_3_0_0),
    .I_3_0_1(n147_I_3_0_1),
    .I_3_0_2(n147_I_3_0_2),
    .I_3_1_0(n147_I_3_1_0),
    .I_3_1_1(n147_I_3_1_1),
    .I_3_1_2(n147_I_3_1_2),
    .I_3_2_0(n147_I_3_2_0),
    .I_3_2_1(n147_I_3_2_1),
    .I_3_2_2(n147_I_3_2_2),
    .I_4_0_0(n147_I_4_0_0),
    .I_4_0_1(n147_I_4_0_1),
    .I_4_0_2(n147_I_4_0_2),
    .I_4_1_0(n147_I_4_1_0),
    .I_4_1_1(n147_I_4_1_1),
    .I_4_1_2(n147_I_4_1_2),
    .I_4_2_0(n147_I_4_2_0),
    .I_4_2_1(n147_I_4_2_1),
    .I_4_2_2(n147_I_4_2_2),
    .I_5_0_0(n147_I_5_0_0),
    .I_5_0_1(n147_I_5_0_1),
    .I_5_0_2(n147_I_5_0_2),
    .I_5_1_0(n147_I_5_1_0),
    .I_5_1_1(n147_I_5_1_1),
    .I_5_1_2(n147_I_5_1_2),
    .I_5_2_0(n147_I_5_2_0),
    .I_5_2_1(n147_I_5_2_1),
    .I_5_2_2(n147_I_5_2_2),
    .I_6_0_0(n147_I_6_0_0),
    .I_6_0_1(n147_I_6_0_1),
    .I_6_0_2(n147_I_6_0_2),
    .I_6_1_0(n147_I_6_1_0),
    .I_6_1_1(n147_I_6_1_1),
    .I_6_1_2(n147_I_6_1_2),
    .I_6_2_0(n147_I_6_2_0),
    .I_6_2_1(n147_I_6_2_1),
    .I_6_2_2(n147_I_6_2_2),
    .I_7_0_0(n147_I_7_0_0),
    .I_7_0_1(n147_I_7_0_1),
    .I_7_0_2(n147_I_7_0_2),
    .I_7_1_0(n147_I_7_1_0),
    .I_7_1_1(n147_I_7_1_1),
    .I_7_1_2(n147_I_7_1_2),
    .I_7_2_0(n147_I_7_2_0),
    .I_7_2_1(n147_I_7_2_1),
    .I_7_2_2(n147_I_7_2_2),
    .I_8_0_0(n147_I_8_0_0),
    .I_8_0_1(n147_I_8_0_1),
    .I_8_0_2(n147_I_8_0_2),
    .I_8_1_0(n147_I_8_1_0),
    .I_8_1_1(n147_I_8_1_1),
    .I_8_1_2(n147_I_8_1_2),
    .I_8_2_0(n147_I_8_2_0),
    .I_8_2_1(n147_I_8_2_1),
    .I_8_2_2(n147_I_8_2_2),
    .I_9_0_0(n147_I_9_0_0),
    .I_9_0_1(n147_I_9_0_1),
    .I_9_0_2(n147_I_9_0_2),
    .I_9_1_0(n147_I_9_1_0),
    .I_9_1_1(n147_I_9_1_1),
    .I_9_1_2(n147_I_9_1_2),
    .I_9_2_0(n147_I_9_2_0),
    .I_9_2_1(n147_I_9_2_1),
    .I_9_2_2(n147_I_9_2_2),
    .I_10_0_0(n147_I_10_0_0),
    .I_10_0_1(n147_I_10_0_1),
    .I_10_0_2(n147_I_10_0_2),
    .I_10_1_0(n147_I_10_1_0),
    .I_10_1_1(n147_I_10_1_1),
    .I_10_1_2(n147_I_10_1_2),
    .I_10_2_0(n147_I_10_2_0),
    .I_10_2_1(n147_I_10_2_1),
    .I_10_2_2(n147_I_10_2_2),
    .I_11_0_0(n147_I_11_0_0),
    .I_11_0_1(n147_I_11_0_1),
    .I_11_0_2(n147_I_11_0_2),
    .I_11_1_0(n147_I_11_1_0),
    .I_11_1_1(n147_I_11_1_1),
    .I_11_1_2(n147_I_11_1_2),
    .I_11_2_0(n147_I_11_2_0),
    .I_11_2_1(n147_I_11_2_1),
    .I_11_2_2(n147_I_11_2_2),
    .I_12_0_0(n147_I_12_0_0),
    .I_12_0_1(n147_I_12_0_1),
    .I_12_0_2(n147_I_12_0_2),
    .I_12_1_0(n147_I_12_1_0),
    .I_12_1_1(n147_I_12_1_1),
    .I_12_1_2(n147_I_12_1_2),
    .I_12_2_0(n147_I_12_2_0),
    .I_12_2_1(n147_I_12_2_1),
    .I_12_2_2(n147_I_12_2_2),
    .I_13_0_0(n147_I_13_0_0),
    .I_13_0_1(n147_I_13_0_1),
    .I_13_0_2(n147_I_13_0_2),
    .I_13_1_0(n147_I_13_1_0),
    .I_13_1_1(n147_I_13_1_1),
    .I_13_1_2(n147_I_13_1_2),
    .I_13_2_0(n147_I_13_2_0),
    .I_13_2_1(n147_I_13_2_1),
    .I_13_2_2(n147_I_13_2_2),
    .I_14_0_0(n147_I_14_0_0),
    .I_14_0_1(n147_I_14_0_1),
    .I_14_0_2(n147_I_14_0_2),
    .I_14_1_0(n147_I_14_1_0),
    .I_14_1_1(n147_I_14_1_1),
    .I_14_1_2(n147_I_14_1_2),
    .I_14_2_0(n147_I_14_2_0),
    .I_14_2_1(n147_I_14_2_1),
    .I_14_2_2(n147_I_14_2_2),
    .I_15_0_0(n147_I_15_0_0),
    .I_15_0_1(n147_I_15_0_1),
    .I_15_0_2(n147_I_15_0_2),
    .I_15_1_0(n147_I_15_1_0),
    .I_15_1_1(n147_I_15_1_1),
    .I_15_1_2(n147_I_15_1_2),
    .I_15_2_0(n147_I_15_2_0),
    .I_15_2_1(n147_I_15_2_1),
    .I_15_2_2(n147_I_15_2_2),
    .O_0_0_0(n147_O_0_0_0),
    .O_1_0_0(n147_O_1_0_0),
    .O_2_0_0(n147_O_2_0_0),
    .O_3_0_0(n147_O_3_0_0),
    .O_4_0_0(n147_O_4_0_0),
    .O_5_0_0(n147_O_5_0_0),
    .O_6_0_0(n147_O_6_0_0),
    .O_7_0_0(n147_O_7_0_0),
    .O_8_0_0(n147_O_8_0_0),
    .O_9_0_0(n147_O_9_0_0),
    .O_10_0_0(n147_O_10_0_0),
    .O_11_0_0(n147_O_11_0_0),
    .O_12_0_0(n147_O_12_0_0),
    .O_13_0_0(n147_O_13_0_0),
    .O_14_0_0(n147_O_14_0_0),
    .O_15_0_0(n147_O_15_0_0)
  );
  Passthrough n148 ( // @[Top.scala 160:22]
    .valid_up(n148_valid_up),
    .valid_down(n148_valid_down),
    .I_0_0_0(n148_I_0_0_0),
    .I_1_0_0(n148_I_1_0_0),
    .I_2_0_0(n148_I_2_0_0),
    .I_3_0_0(n148_I_3_0_0),
    .I_4_0_0(n148_I_4_0_0),
    .I_5_0_0(n148_I_5_0_0),
    .I_6_0_0(n148_I_6_0_0),
    .I_7_0_0(n148_I_7_0_0),
    .I_8_0_0(n148_I_8_0_0),
    .I_9_0_0(n148_I_9_0_0),
    .I_10_0_0(n148_I_10_0_0),
    .I_11_0_0(n148_I_11_0_0),
    .I_12_0_0(n148_I_12_0_0),
    .I_13_0_0(n148_I_13_0_0),
    .I_14_0_0(n148_I_14_0_0),
    .I_15_0_0(n148_I_15_0_0),
    .O_0_0(n148_O_0_0),
    .O_1_0(n148_O_1_0),
    .O_2_0(n148_O_2_0),
    .O_3_0(n148_O_3_0),
    .O_4_0(n148_O_4_0),
    .O_5_0(n148_O_5_0),
    .O_6_0(n148_O_6_0),
    .O_7_0(n148_O_7_0),
    .O_8_0(n148_O_8_0),
    .O_9_0(n148_O_9_0),
    .O_10_0(n148_O_10_0),
    .O_11_0(n148_O_11_0),
    .O_12_0(n148_O_12_0),
    .O_13_0(n148_O_13_0),
    .O_14_0(n148_O_14_0),
    .O_15_0(n148_O_15_0)
  );
  Passthrough_1 n149 ( // @[Top.scala 163:22]
    .valid_up(n149_valid_up),
    .valid_down(n149_valid_down),
    .I_0_0(n149_I_0_0),
    .I_1_0(n149_I_1_0),
    .I_2_0(n149_I_2_0),
    .I_3_0(n149_I_3_0),
    .I_4_0(n149_I_4_0),
    .I_5_0(n149_I_5_0),
    .I_6_0(n149_I_6_0),
    .I_7_0(n149_I_7_0),
    .I_8_0(n149_I_8_0),
    .I_9_0(n149_I_9_0),
    .I_10_0(n149_I_10_0),
    .I_11_0(n149_I_11_0),
    .I_12_0(n149_I_12_0),
    .I_13_0(n149_I_13_0),
    .I_14_0(n149_I_14_0),
    .I_15_0(n149_I_15_0),
    .O_0(n149_O_0),
    .O_1(n149_O_1),
    .O_2(n149_O_2),
    .O_3(n149_O_3),
    .O_4(n149_O_4),
    .O_5(n149_O_5),
    .O_6(n149_O_6),
    .O_7(n149_O_7),
    .O_8(n149_O_8),
    .O_9(n149_O_9),
    .O_10(n149_O_10),
    .O_11(n149_O_11),
    .O_12(n149_O_12),
    .O_13(n149_O_13),
    .O_14(n149_O_14),
    .O_15(n149_O_15)
  );
  ShiftTS n150 ( // @[Top.scala 166:22]
    .clock(n150_clock),
    .reset(n150_reset),
    .valid_up(n150_valid_up),
    .valid_down(n150_valid_down),
    .I_0(n150_I_0),
    .I_1(n150_I_1),
    .I_2(n150_I_2),
    .I_3(n150_I_3),
    .I_4(n150_I_4),
    .I_5(n150_I_5),
    .I_6(n150_I_6),
    .I_7(n150_I_7),
    .I_8(n150_I_8),
    .I_9(n150_I_9),
    .I_10(n150_I_10),
    .I_11(n150_I_11),
    .I_12(n150_I_12),
    .I_13(n150_I_13),
    .I_14(n150_I_14),
    .I_15(n150_I_15),
    .O_0(n150_O_0),
    .O_1(n150_O_1),
    .O_2(n150_O_2),
    .O_3(n150_O_3),
    .O_4(n150_O_4),
    .O_5(n150_O_5),
    .O_6(n150_O_6),
    .O_7(n150_O_7),
    .O_8(n150_O_8),
    .O_9(n150_O_9),
    .O_10(n150_O_10),
    .O_11(n150_O_11),
    .O_12(n150_O_12),
    .O_13(n150_O_13),
    .O_14(n150_O_14),
    .O_15(n150_O_15)
  );
  ShiftTS_2 n151 ( // @[Top.scala 169:22]
    .clock(n151_clock),
    .valid_up(n151_valid_up),
    .valid_down(n151_valid_down),
    .I_0(n151_I_0),
    .I_1(n151_I_1),
    .I_2(n151_I_2),
    .I_3(n151_I_3),
    .I_4(n151_I_4),
    .I_5(n151_I_5),
    .I_6(n151_I_6),
    .I_7(n151_I_7),
    .I_8(n151_I_8),
    .I_9(n151_I_9),
    .I_10(n151_I_10),
    .I_11(n151_I_11),
    .I_12(n151_I_12),
    .I_13(n151_I_13),
    .I_14(n151_I_14),
    .I_15(n151_I_15),
    .O_0(n151_O_0),
    .O_1(n151_O_1),
    .O_2(n151_O_2),
    .O_3(n151_O_3),
    .O_4(n151_O_4),
    .O_5(n151_O_5),
    .O_6(n151_O_6),
    .O_7(n151_O_7),
    .O_8(n151_O_8),
    .O_9(n151_O_9),
    .O_10(n151_O_10),
    .O_11(n151_O_11),
    .O_12(n151_O_12),
    .O_13(n151_O_13),
    .O_14(n151_O_14),
    .O_15(n151_O_15)
  );
  Map2T n152 ( // @[Top.scala 172:22]
    .valid_up(n152_valid_up),
    .valid_down(n152_valid_down),
    .I0_0(n152_I0_0),
    .I0_1(n152_I0_1),
    .I0_2(n152_I0_2),
    .I0_3(n152_I0_3),
    .I0_4(n152_I0_4),
    .I0_5(n152_I0_5),
    .I0_6(n152_I0_6),
    .I0_7(n152_I0_7),
    .I0_8(n152_I0_8),
    .I0_9(n152_I0_9),
    .I0_10(n152_I0_10),
    .I0_11(n152_I0_11),
    .I0_12(n152_I0_12),
    .I0_13(n152_I0_13),
    .I0_14(n152_I0_14),
    .I0_15(n152_I0_15),
    .I1_0(n152_I1_0),
    .I1_1(n152_I1_1),
    .I1_2(n152_I1_2),
    .I1_3(n152_I1_3),
    .I1_4(n152_I1_4),
    .I1_5(n152_I1_5),
    .I1_6(n152_I1_6),
    .I1_7(n152_I1_7),
    .I1_8(n152_I1_8),
    .I1_9(n152_I1_9),
    .I1_10(n152_I1_10),
    .I1_11(n152_I1_11),
    .I1_12(n152_I1_12),
    .I1_13(n152_I1_13),
    .I1_14(n152_I1_14),
    .I1_15(n152_I1_15),
    .O_0_0(n152_O_0_0),
    .O_0_1(n152_O_0_1),
    .O_1_0(n152_O_1_0),
    .O_1_1(n152_O_1_1),
    .O_2_0(n152_O_2_0),
    .O_2_1(n152_O_2_1),
    .O_3_0(n152_O_3_0),
    .O_3_1(n152_O_3_1),
    .O_4_0(n152_O_4_0),
    .O_4_1(n152_O_4_1),
    .O_5_0(n152_O_5_0),
    .O_5_1(n152_O_5_1),
    .O_6_0(n152_O_6_0),
    .O_6_1(n152_O_6_1),
    .O_7_0(n152_O_7_0),
    .O_7_1(n152_O_7_1),
    .O_8_0(n152_O_8_0),
    .O_8_1(n152_O_8_1),
    .O_9_0(n152_O_9_0),
    .O_9_1(n152_O_9_1),
    .O_10_0(n152_O_10_0),
    .O_10_1(n152_O_10_1),
    .O_11_0(n152_O_11_0),
    .O_11_1(n152_O_11_1),
    .O_12_0(n152_O_12_0),
    .O_12_1(n152_O_12_1),
    .O_13_0(n152_O_13_0),
    .O_13_1(n152_O_13_1),
    .O_14_0(n152_O_14_0),
    .O_14_1(n152_O_14_1),
    .O_15_0(n152_O_15_0),
    .O_15_1(n152_O_15_1)
  );
  MapT_9 n161 ( // @[Top.scala 176:22]
    .valid_up(n161_valid_up),
    .valid_down(n161_valid_down),
    .I_0_0(n161_I_0_0),
    .I_0_1(n161_I_0_1),
    .I_1_0(n161_I_1_0),
    .I_1_1(n161_I_1_1),
    .I_2_0(n161_I_2_0),
    .I_2_1(n161_I_2_1),
    .I_3_0(n161_I_3_0),
    .I_3_1(n161_I_3_1),
    .I_4_0(n161_I_4_0),
    .I_4_1(n161_I_4_1),
    .I_5_0(n161_I_5_0),
    .I_5_1(n161_I_5_1),
    .I_6_0(n161_I_6_0),
    .I_6_1(n161_I_6_1),
    .I_7_0(n161_I_7_0),
    .I_7_1(n161_I_7_1),
    .I_8_0(n161_I_8_0),
    .I_8_1(n161_I_8_1),
    .I_9_0(n161_I_9_0),
    .I_9_1(n161_I_9_1),
    .I_10_0(n161_I_10_0),
    .I_10_1(n161_I_10_1),
    .I_11_0(n161_I_11_0),
    .I_11_1(n161_I_11_1),
    .I_12_0(n161_I_12_0),
    .I_12_1(n161_I_12_1),
    .I_13_0(n161_I_13_0),
    .I_13_1(n161_I_13_1),
    .I_14_0(n161_I_14_0),
    .I_14_1(n161_I_14_1),
    .I_15_0(n161_I_15_0),
    .I_15_1(n161_I_15_1),
    .O_0_0_0(n161_O_0_0_0),
    .O_0_0_1(n161_O_0_0_1),
    .O_1_0_0(n161_O_1_0_0),
    .O_1_0_1(n161_O_1_0_1),
    .O_2_0_0(n161_O_2_0_0),
    .O_2_0_1(n161_O_2_0_1),
    .O_3_0_0(n161_O_3_0_0),
    .O_3_0_1(n161_O_3_0_1),
    .O_4_0_0(n161_O_4_0_0),
    .O_4_0_1(n161_O_4_0_1),
    .O_5_0_0(n161_O_5_0_0),
    .O_5_0_1(n161_O_5_0_1),
    .O_6_0_0(n161_O_6_0_0),
    .O_6_0_1(n161_O_6_0_1),
    .O_7_0_0(n161_O_7_0_0),
    .O_7_0_1(n161_O_7_0_1),
    .O_8_0_0(n161_O_8_0_0),
    .O_8_0_1(n161_O_8_0_1),
    .O_9_0_0(n161_O_9_0_0),
    .O_9_0_1(n161_O_9_0_1),
    .O_10_0_0(n161_O_10_0_0),
    .O_10_0_1(n161_O_10_0_1),
    .O_11_0_0(n161_O_11_0_0),
    .O_11_0_1(n161_O_11_0_1),
    .O_12_0_0(n161_O_12_0_0),
    .O_12_0_1(n161_O_12_0_1),
    .O_13_0_0(n161_O_13_0_0),
    .O_13_0_1(n161_O_13_0_1),
    .O_14_0_0(n161_O_14_0_0),
    .O_14_0_1(n161_O_14_0_1),
    .O_15_0_0(n161_O_15_0_0),
    .O_15_0_1(n161_O_15_0_1)
  );
  MapT_10 n168 ( // @[Top.scala 179:22]
    .valid_up(n168_valid_up),
    .valid_down(n168_valid_down),
    .I_0_0_0(n168_I_0_0_0),
    .I_0_0_1(n168_I_0_0_1),
    .I_1_0_0(n168_I_1_0_0),
    .I_1_0_1(n168_I_1_0_1),
    .I_2_0_0(n168_I_2_0_0),
    .I_2_0_1(n168_I_2_0_1),
    .I_3_0_0(n168_I_3_0_0),
    .I_3_0_1(n168_I_3_0_1),
    .I_4_0_0(n168_I_4_0_0),
    .I_4_0_1(n168_I_4_0_1),
    .I_5_0_0(n168_I_5_0_0),
    .I_5_0_1(n168_I_5_0_1),
    .I_6_0_0(n168_I_6_0_0),
    .I_6_0_1(n168_I_6_0_1),
    .I_7_0_0(n168_I_7_0_0),
    .I_7_0_1(n168_I_7_0_1),
    .I_8_0_0(n168_I_8_0_0),
    .I_8_0_1(n168_I_8_0_1),
    .I_9_0_0(n168_I_9_0_0),
    .I_9_0_1(n168_I_9_0_1),
    .I_10_0_0(n168_I_10_0_0),
    .I_10_0_1(n168_I_10_0_1),
    .I_11_0_0(n168_I_11_0_0),
    .I_11_0_1(n168_I_11_0_1),
    .I_12_0_0(n168_I_12_0_0),
    .I_12_0_1(n168_I_12_0_1),
    .I_13_0_0(n168_I_13_0_0),
    .I_13_0_1(n168_I_13_0_1),
    .I_14_0_0(n168_I_14_0_0),
    .I_14_0_1(n168_I_14_0_1),
    .I_15_0_0(n168_I_15_0_0),
    .I_15_0_1(n168_I_15_0_1),
    .O_0_0(n168_O_0_0),
    .O_0_1(n168_O_0_1),
    .O_1_0(n168_O_1_0),
    .O_1_1(n168_O_1_1),
    .O_2_0(n168_O_2_0),
    .O_2_1(n168_O_2_1),
    .O_3_0(n168_O_3_0),
    .O_3_1(n168_O_3_1),
    .O_4_0(n168_O_4_0),
    .O_4_1(n168_O_4_1),
    .O_5_0(n168_O_5_0),
    .O_5_1(n168_O_5_1),
    .O_6_0(n168_O_6_0),
    .O_6_1(n168_O_6_1),
    .O_7_0(n168_O_7_0),
    .O_7_1(n168_O_7_1),
    .O_8_0(n168_O_8_0),
    .O_8_1(n168_O_8_1),
    .O_9_0(n168_O_9_0),
    .O_9_1(n168_O_9_1),
    .O_10_0(n168_O_10_0),
    .O_10_1(n168_O_10_1),
    .O_11_0(n168_O_11_0),
    .O_11_1(n168_O_11_1),
    .O_12_0(n168_O_12_0),
    .O_12_1(n168_O_12_1),
    .O_13_0(n168_O_13_0),
    .O_13_1(n168_O_13_1),
    .O_14_0(n168_O_14_0),
    .O_14_1(n168_O_14_1),
    .O_15_0(n168_O_15_0),
    .O_15_1(n168_O_15_1)
  );
  ShiftTS_2 n169 ( // @[Top.scala 182:22]
    .clock(n169_clock),
    .valid_up(n169_valid_up),
    .valid_down(n169_valid_down),
    .I_0(n169_I_0),
    .I_1(n169_I_1),
    .I_2(n169_I_2),
    .I_3(n169_I_3),
    .I_4(n169_I_4),
    .I_5(n169_I_5),
    .I_6(n169_I_6),
    .I_7(n169_I_7),
    .I_8(n169_I_8),
    .I_9(n169_I_9),
    .I_10(n169_I_10),
    .I_11(n169_I_11),
    .I_12(n169_I_12),
    .I_13(n169_I_13),
    .I_14(n169_I_14),
    .I_15(n169_I_15),
    .O_0(n169_O_0),
    .O_1(n169_O_1),
    .O_2(n169_O_2),
    .O_3(n169_O_3),
    .O_4(n169_O_4),
    .O_5(n169_O_5),
    .O_6(n169_O_6),
    .O_7(n169_O_7),
    .O_8(n169_O_8),
    .O_9(n169_O_9),
    .O_10(n169_O_10),
    .O_11(n169_O_11),
    .O_12(n169_O_12),
    .O_13(n169_O_13),
    .O_14(n169_O_14),
    .O_15(n169_O_15)
  );
  Map2T n170 ( // @[Top.scala 185:22]
    .valid_up(n170_valid_up),
    .valid_down(n170_valid_down),
    .I0_0(n170_I0_0),
    .I0_1(n170_I0_1),
    .I0_2(n170_I0_2),
    .I0_3(n170_I0_3),
    .I0_4(n170_I0_4),
    .I0_5(n170_I0_5),
    .I0_6(n170_I0_6),
    .I0_7(n170_I0_7),
    .I0_8(n170_I0_8),
    .I0_9(n170_I0_9),
    .I0_10(n170_I0_10),
    .I0_11(n170_I0_11),
    .I0_12(n170_I0_12),
    .I0_13(n170_I0_13),
    .I0_14(n170_I0_14),
    .I0_15(n170_I0_15),
    .I1_0(n170_I1_0),
    .I1_1(n170_I1_1),
    .I1_2(n170_I1_2),
    .I1_3(n170_I1_3),
    .I1_4(n170_I1_4),
    .I1_5(n170_I1_5),
    .I1_6(n170_I1_6),
    .I1_7(n170_I1_7),
    .I1_8(n170_I1_8),
    .I1_9(n170_I1_9),
    .I1_10(n170_I1_10),
    .I1_11(n170_I1_11),
    .I1_12(n170_I1_12),
    .I1_13(n170_I1_13),
    .I1_14(n170_I1_14),
    .I1_15(n170_I1_15),
    .O_0_0(n170_O_0_0),
    .O_0_1(n170_O_0_1),
    .O_1_0(n170_O_1_0),
    .O_1_1(n170_O_1_1),
    .O_2_0(n170_O_2_0),
    .O_2_1(n170_O_2_1),
    .O_3_0(n170_O_3_0),
    .O_3_1(n170_O_3_1),
    .O_4_0(n170_O_4_0),
    .O_4_1(n170_O_4_1),
    .O_5_0(n170_O_5_0),
    .O_5_1(n170_O_5_1),
    .O_6_0(n170_O_6_0),
    .O_6_1(n170_O_6_1),
    .O_7_0(n170_O_7_0),
    .O_7_1(n170_O_7_1),
    .O_8_0(n170_O_8_0),
    .O_8_1(n170_O_8_1),
    .O_9_0(n170_O_9_0),
    .O_9_1(n170_O_9_1),
    .O_10_0(n170_O_10_0),
    .O_10_1(n170_O_10_1),
    .O_11_0(n170_O_11_0),
    .O_11_1(n170_O_11_1),
    .O_12_0(n170_O_12_0),
    .O_12_1(n170_O_12_1),
    .O_13_0(n170_O_13_0),
    .O_13_1(n170_O_13_1),
    .O_14_0(n170_O_14_0),
    .O_14_1(n170_O_14_1),
    .O_15_0(n170_O_15_0),
    .O_15_1(n170_O_15_1)
  );
  MapT_9 n179 ( // @[Top.scala 189:22]
    .valid_up(n179_valid_up),
    .valid_down(n179_valid_down),
    .I_0_0(n179_I_0_0),
    .I_0_1(n179_I_0_1),
    .I_1_0(n179_I_1_0),
    .I_1_1(n179_I_1_1),
    .I_2_0(n179_I_2_0),
    .I_2_1(n179_I_2_1),
    .I_3_0(n179_I_3_0),
    .I_3_1(n179_I_3_1),
    .I_4_0(n179_I_4_0),
    .I_4_1(n179_I_4_1),
    .I_5_0(n179_I_5_0),
    .I_5_1(n179_I_5_1),
    .I_6_0(n179_I_6_0),
    .I_6_1(n179_I_6_1),
    .I_7_0(n179_I_7_0),
    .I_7_1(n179_I_7_1),
    .I_8_0(n179_I_8_0),
    .I_8_1(n179_I_8_1),
    .I_9_0(n179_I_9_0),
    .I_9_1(n179_I_9_1),
    .I_10_0(n179_I_10_0),
    .I_10_1(n179_I_10_1),
    .I_11_0(n179_I_11_0),
    .I_11_1(n179_I_11_1),
    .I_12_0(n179_I_12_0),
    .I_12_1(n179_I_12_1),
    .I_13_0(n179_I_13_0),
    .I_13_1(n179_I_13_1),
    .I_14_0(n179_I_14_0),
    .I_14_1(n179_I_14_1),
    .I_15_0(n179_I_15_0),
    .I_15_1(n179_I_15_1),
    .O_0_0_0(n179_O_0_0_0),
    .O_0_0_1(n179_O_0_0_1),
    .O_1_0_0(n179_O_1_0_0),
    .O_1_0_1(n179_O_1_0_1),
    .O_2_0_0(n179_O_2_0_0),
    .O_2_0_1(n179_O_2_0_1),
    .O_3_0_0(n179_O_3_0_0),
    .O_3_0_1(n179_O_3_0_1),
    .O_4_0_0(n179_O_4_0_0),
    .O_4_0_1(n179_O_4_0_1),
    .O_5_0_0(n179_O_5_0_0),
    .O_5_0_1(n179_O_5_0_1),
    .O_6_0_0(n179_O_6_0_0),
    .O_6_0_1(n179_O_6_0_1),
    .O_7_0_0(n179_O_7_0_0),
    .O_7_0_1(n179_O_7_0_1),
    .O_8_0_0(n179_O_8_0_0),
    .O_8_0_1(n179_O_8_0_1),
    .O_9_0_0(n179_O_9_0_0),
    .O_9_0_1(n179_O_9_0_1),
    .O_10_0_0(n179_O_10_0_0),
    .O_10_0_1(n179_O_10_0_1),
    .O_11_0_0(n179_O_11_0_0),
    .O_11_0_1(n179_O_11_0_1),
    .O_12_0_0(n179_O_12_0_0),
    .O_12_0_1(n179_O_12_0_1),
    .O_13_0_0(n179_O_13_0_0),
    .O_13_0_1(n179_O_13_0_1),
    .O_14_0_0(n179_O_14_0_0),
    .O_14_0_1(n179_O_14_0_1),
    .O_15_0_0(n179_O_15_0_0),
    .O_15_0_1(n179_O_15_0_1)
  );
  MapT_10 n186 ( // @[Top.scala 192:22]
    .valid_up(n186_valid_up),
    .valid_down(n186_valid_down),
    .I_0_0_0(n186_I_0_0_0),
    .I_0_0_1(n186_I_0_0_1),
    .I_1_0_0(n186_I_1_0_0),
    .I_1_0_1(n186_I_1_0_1),
    .I_2_0_0(n186_I_2_0_0),
    .I_2_0_1(n186_I_2_0_1),
    .I_3_0_0(n186_I_3_0_0),
    .I_3_0_1(n186_I_3_0_1),
    .I_4_0_0(n186_I_4_0_0),
    .I_4_0_1(n186_I_4_0_1),
    .I_5_0_0(n186_I_5_0_0),
    .I_5_0_1(n186_I_5_0_1),
    .I_6_0_0(n186_I_6_0_0),
    .I_6_0_1(n186_I_6_0_1),
    .I_7_0_0(n186_I_7_0_0),
    .I_7_0_1(n186_I_7_0_1),
    .I_8_0_0(n186_I_8_0_0),
    .I_8_0_1(n186_I_8_0_1),
    .I_9_0_0(n186_I_9_0_0),
    .I_9_0_1(n186_I_9_0_1),
    .I_10_0_0(n186_I_10_0_0),
    .I_10_0_1(n186_I_10_0_1),
    .I_11_0_0(n186_I_11_0_0),
    .I_11_0_1(n186_I_11_0_1),
    .I_12_0_0(n186_I_12_0_0),
    .I_12_0_1(n186_I_12_0_1),
    .I_13_0_0(n186_I_13_0_0),
    .I_13_0_1(n186_I_13_0_1),
    .I_14_0_0(n186_I_14_0_0),
    .I_14_0_1(n186_I_14_0_1),
    .I_15_0_0(n186_I_15_0_0),
    .I_15_0_1(n186_I_15_0_1),
    .O_0_0(n186_O_0_0),
    .O_0_1(n186_O_0_1),
    .O_1_0(n186_O_1_0),
    .O_1_1(n186_O_1_1),
    .O_2_0(n186_O_2_0),
    .O_2_1(n186_O_2_1),
    .O_3_0(n186_O_3_0),
    .O_3_1(n186_O_3_1),
    .O_4_0(n186_O_4_0),
    .O_4_1(n186_O_4_1),
    .O_5_0(n186_O_5_0),
    .O_5_1(n186_O_5_1),
    .O_6_0(n186_O_6_0),
    .O_6_1(n186_O_6_1),
    .O_7_0(n186_O_7_0),
    .O_7_1(n186_O_7_1),
    .O_8_0(n186_O_8_0),
    .O_8_1(n186_O_8_1),
    .O_9_0(n186_O_9_0),
    .O_9_1(n186_O_9_1),
    .O_10_0(n186_O_10_0),
    .O_10_1(n186_O_10_1),
    .O_11_0(n186_O_11_0),
    .O_11_1(n186_O_11_1),
    .O_12_0(n186_O_12_0),
    .O_12_1(n186_O_12_1),
    .O_13_0(n186_O_13_0),
    .O_13_1(n186_O_13_1),
    .O_14_0(n186_O_14_0),
    .O_14_1(n186_O_14_1),
    .O_15_0(n186_O_15_0),
    .O_15_1(n186_O_15_1)
  );
  Map2T_10 n187 ( // @[Top.scala 195:22]
    .valid_up(n187_valid_up),
    .valid_down(n187_valid_down),
    .I0_0_0(n187_I0_0_0),
    .I0_0_1(n187_I0_0_1),
    .I0_1_0(n187_I0_1_0),
    .I0_1_1(n187_I0_1_1),
    .I0_2_0(n187_I0_2_0),
    .I0_2_1(n187_I0_2_1),
    .I0_3_0(n187_I0_3_0),
    .I0_3_1(n187_I0_3_1),
    .I0_4_0(n187_I0_4_0),
    .I0_4_1(n187_I0_4_1),
    .I0_5_0(n187_I0_5_0),
    .I0_5_1(n187_I0_5_1),
    .I0_6_0(n187_I0_6_0),
    .I0_6_1(n187_I0_6_1),
    .I0_7_0(n187_I0_7_0),
    .I0_7_1(n187_I0_7_1),
    .I0_8_0(n187_I0_8_0),
    .I0_8_1(n187_I0_8_1),
    .I0_9_0(n187_I0_9_0),
    .I0_9_1(n187_I0_9_1),
    .I0_10_0(n187_I0_10_0),
    .I0_10_1(n187_I0_10_1),
    .I0_11_0(n187_I0_11_0),
    .I0_11_1(n187_I0_11_1),
    .I0_12_0(n187_I0_12_0),
    .I0_12_1(n187_I0_12_1),
    .I0_13_0(n187_I0_13_0),
    .I0_13_1(n187_I0_13_1),
    .I0_14_0(n187_I0_14_0),
    .I0_14_1(n187_I0_14_1),
    .I0_15_0(n187_I0_15_0),
    .I0_15_1(n187_I0_15_1),
    .I1_0_0(n187_I1_0_0),
    .I1_0_1(n187_I1_0_1),
    .I1_1_0(n187_I1_1_0),
    .I1_1_1(n187_I1_1_1),
    .I1_2_0(n187_I1_2_0),
    .I1_2_1(n187_I1_2_1),
    .I1_3_0(n187_I1_3_0),
    .I1_3_1(n187_I1_3_1),
    .I1_4_0(n187_I1_4_0),
    .I1_4_1(n187_I1_4_1),
    .I1_5_0(n187_I1_5_0),
    .I1_5_1(n187_I1_5_1),
    .I1_6_0(n187_I1_6_0),
    .I1_6_1(n187_I1_6_1),
    .I1_7_0(n187_I1_7_0),
    .I1_7_1(n187_I1_7_1),
    .I1_8_0(n187_I1_8_0),
    .I1_8_1(n187_I1_8_1),
    .I1_9_0(n187_I1_9_0),
    .I1_9_1(n187_I1_9_1),
    .I1_10_0(n187_I1_10_0),
    .I1_10_1(n187_I1_10_1),
    .I1_11_0(n187_I1_11_0),
    .I1_11_1(n187_I1_11_1),
    .I1_12_0(n187_I1_12_0),
    .I1_12_1(n187_I1_12_1),
    .I1_13_0(n187_I1_13_0),
    .I1_13_1(n187_I1_13_1),
    .I1_14_0(n187_I1_14_0),
    .I1_14_1(n187_I1_14_1),
    .I1_15_0(n187_I1_15_0),
    .I1_15_1(n187_I1_15_1),
    .O_0_0_0(n187_O_0_0_0),
    .O_0_0_1(n187_O_0_0_1),
    .O_0_1_0(n187_O_0_1_0),
    .O_0_1_1(n187_O_0_1_1),
    .O_1_0_0(n187_O_1_0_0),
    .O_1_0_1(n187_O_1_0_1),
    .O_1_1_0(n187_O_1_1_0),
    .O_1_1_1(n187_O_1_1_1),
    .O_2_0_0(n187_O_2_0_0),
    .O_2_0_1(n187_O_2_0_1),
    .O_2_1_0(n187_O_2_1_0),
    .O_2_1_1(n187_O_2_1_1),
    .O_3_0_0(n187_O_3_0_0),
    .O_3_0_1(n187_O_3_0_1),
    .O_3_1_0(n187_O_3_1_0),
    .O_3_1_1(n187_O_3_1_1),
    .O_4_0_0(n187_O_4_0_0),
    .O_4_0_1(n187_O_4_0_1),
    .O_4_1_0(n187_O_4_1_0),
    .O_4_1_1(n187_O_4_1_1),
    .O_5_0_0(n187_O_5_0_0),
    .O_5_0_1(n187_O_5_0_1),
    .O_5_1_0(n187_O_5_1_0),
    .O_5_1_1(n187_O_5_1_1),
    .O_6_0_0(n187_O_6_0_0),
    .O_6_0_1(n187_O_6_0_1),
    .O_6_1_0(n187_O_6_1_0),
    .O_6_1_1(n187_O_6_1_1),
    .O_7_0_0(n187_O_7_0_0),
    .O_7_0_1(n187_O_7_0_1),
    .O_7_1_0(n187_O_7_1_0),
    .O_7_1_1(n187_O_7_1_1),
    .O_8_0_0(n187_O_8_0_0),
    .O_8_0_1(n187_O_8_0_1),
    .O_8_1_0(n187_O_8_1_0),
    .O_8_1_1(n187_O_8_1_1),
    .O_9_0_0(n187_O_9_0_0),
    .O_9_0_1(n187_O_9_0_1),
    .O_9_1_0(n187_O_9_1_0),
    .O_9_1_1(n187_O_9_1_1),
    .O_10_0_0(n187_O_10_0_0),
    .O_10_0_1(n187_O_10_0_1),
    .O_10_1_0(n187_O_10_1_0),
    .O_10_1_1(n187_O_10_1_1),
    .O_11_0_0(n187_O_11_0_0),
    .O_11_0_1(n187_O_11_0_1),
    .O_11_1_0(n187_O_11_1_0),
    .O_11_1_1(n187_O_11_1_1),
    .O_12_0_0(n187_O_12_0_0),
    .O_12_0_1(n187_O_12_0_1),
    .O_12_1_0(n187_O_12_1_0),
    .O_12_1_1(n187_O_12_1_1),
    .O_13_0_0(n187_O_13_0_0),
    .O_13_0_1(n187_O_13_0_1),
    .O_13_1_0(n187_O_13_1_0),
    .O_13_1_1(n187_O_13_1_1),
    .O_14_0_0(n187_O_14_0_0),
    .O_14_0_1(n187_O_14_0_1),
    .O_14_1_0(n187_O_14_1_0),
    .O_14_1_1(n187_O_14_1_1),
    .O_15_0_0(n187_O_15_0_0),
    .O_15_0_1(n187_O_15_0_1),
    .O_15_1_0(n187_O_15_1_0),
    .O_15_1_1(n187_O_15_1_1)
  );
  MapT_13 n196 ( // @[Top.scala 199:22]
    .valid_up(n196_valid_up),
    .valid_down(n196_valid_down),
    .I_0_0_0(n196_I_0_0_0),
    .I_0_0_1(n196_I_0_0_1),
    .I_0_1_0(n196_I_0_1_0),
    .I_0_1_1(n196_I_0_1_1),
    .I_1_0_0(n196_I_1_0_0),
    .I_1_0_1(n196_I_1_0_1),
    .I_1_1_0(n196_I_1_1_0),
    .I_1_1_1(n196_I_1_1_1),
    .I_2_0_0(n196_I_2_0_0),
    .I_2_0_1(n196_I_2_0_1),
    .I_2_1_0(n196_I_2_1_0),
    .I_2_1_1(n196_I_2_1_1),
    .I_3_0_0(n196_I_3_0_0),
    .I_3_0_1(n196_I_3_0_1),
    .I_3_1_0(n196_I_3_1_0),
    .I_3_1_1(n196_I_3_1_1),
    .I_4_0_0(n196_I_4_0_0),
    .I_4_0_1(n196_I_4_0_1),
    .I_4_1_0(n196_I_4_1_0),
    .I_4_1_1(n196_I_4_1_1),
    .I_5_0_0(n196_I_5_0_0),
    .I_5_0_1(n196_I_5_0_1),
    .I_5_1_0(n196_I_5_1_0),
    .I_5_1_1(n196_I_5_1_1),
    .I_6_0_0(n196_I_6_0_0),
    .I_6_0_1(n196_I_6_0_1),
    .I_6_1_0(n196_I_6_1_0),
    .I_6_1_1(n196_I_6_1_1),
    .I_7_0_0(n196_I_7_0_0),
    .I_7_0_1(n196_I_7_0_1),
    .I_7_1_0(n196_I_7_1_0),
    .I_7_1_1(n196_I_7_1_1),
    .I_8_0_0(n196_I_8_0_0),
    .I_8_0_1(n196_I_8_0_1),
    .I_8_1_0(n196_I_8_1_0),
    .I_8_1_1(n196_I_8_1_1),
    .I_9_0_0(n196_I_9_0_0),
    .I_9_0_1(n196_I_9_0_1),
    .I_9_1_0(n196_I_9_1_0),
    .I_9_1_1(n196_I_9_1_1),
    .I_10_0_0(n196_I_10_0_0),
    .I_10_0_1(n196_I_10_0_1),
    .I_10_1_0(n196_I_10_1_0),
    .I_10_1_1(n196_I_10_1_1),
    .I_11_0_0(n196_I_11_0_0),
    .I_11_0_1(n196_I_11_0_1),
    .I_11_1_0(n196_I_11_1_0),
    .I_11_1_1(n196_I_11_1_1),
    .I_12_0_0(n196_I_12_0_0),
    .I_12_0_1(n196_I_12_0_1),
    .I_12_1_0(n196_I_12_1_0),
    .I_12_1_1(n196_I_12_1_1),
    .I_13_0_0(n196_I_13_0_0),
    .I_13_0_1(n196_I_13_0_1),
    .I_13_1_0(n196_I_13_1_0),
    .I_13_1_1(n196_I_13_1_1),
    .I_14_0_0(n196_I_14_0_0),
    .I_14_0_1(n196_I_14_0_1),
    .I_14_1_0(n196_I_14_1_0),
    .I_14_1_1(n196_I_14_1_1),
    .I_15_0_0(n196_I_15_0_0),
    .I_15_0_1(n196_I_15_0_1),
    .I_15_1_0(n196_I_15_1_0),
    .I_15_1_1(n196_I_15_1_1),
    .O_0_0_0_0(n196_O_0_0_0_0),
    .O_0_0_0_1(n196_O_0_0_0_1),
    .O_0_0_1_0(n196_O_0_0_1_0),
    .O_0_0_1_1(n196_O_0_0_1_1),
    .O_1_0_0_0(n196_O_1_0_0_0),
    .O_1_0_0_1(n196_O_1_0_0_1),
    .O_1_0_1_0(n196_O_1_0_1_0),
    .O_1_0_1_1(n196_O_1_0_1_1),
    .O_2_0_0_0(n196_O_2_0_0_0),
    .O_2_0_0_1(n196_O_2_0_0_1),
    .O_2_0_1_0(n196_O_2_0_1_0),
    .O_2_0_1_1(n196_O_2_0_1_1),
    .O_3_0_0_0(n196_O_3_0_0_0),
    .O_3_0_0_1(n196_O_3_0_0_1),
    .O_3_0_1_0(n196_O_3_0_1_0),
    .O_3_0_1_1(n196_O_3_0_1_1),
    .O_4_0_0_0(n196_O_4_0_0_0),
    .O_4_0_0_1(n196_O_4_0_0_1),
    .O_4_0_1_0(n196_O_4_0_1_0),
    .O_4_0_1_1(n196_O_4_0_1_1),
    .O_5_0_0_0(n196_O_5_0_0_0),
    .O_5_0_0_1(n196_O_5_0_0_1),
    .O_5_0_1_0(n196_O_5_0_1_0),
    .O_5_0_1_1(n196_O_5_0_1_1),
    .O_6_0_0_0(n196_O_6_0_0_0),
    .O_6_0_0_1(n196_O_6_0_0_1),
    .O_6_0_1_0(n196_O_6_0_1_0),
    .O_6_0_1_1(n196_O_6_0_1_1),
    .O_7_0_0_0(n196_O_7_0_0_0),
    .O_7_0_0_1(n196_O_7_0_0_1),
    .O_7_0_1_0(n196_O_7_0_1_0),
    .O_7_0_1_1(n196_O_7_0_1_1),
    .O_8_0_0_0(n196_O_8_0_0_0),
    .O_8_0_0_1(n196_O_8_0_0_1),
    .O_8_0_1_0(n196_O_8_0_1_0),
    .O_8_0_1_1(n196_O_8_0_1_1),
    .O_9_0_0_0(n196_O_9_0_0_0),
    .O_9_0_0_1(n196_O_9_0_0_1),
    .O_9_0_1_0(n196_O_9_0_1_0),
    .O_9_0_1_1(n196_O_9_0_1_1),
    .O_10_0_0_0(n196_O_10_0_0_0),
    .O_10_0_0_1(n196_O_10_0_0_1),
    .O_10_0_1_0(n196_O_10_0_1_0),
    .O_10_0_1_1(n196_O_10_0_1_1),
    .O_11_0_0_0(n196_O_11_0_0_0),
    .O_11_0_0_1(n196_O_11_0_0_1),
    .O_11_0_1_0(n196_O_11_0_1_0),
    .O_11_0_1_1(n196_O_11_0_1_1),
    .O_12_0_0_0(n196_O_12_0_0_0),
    .O_12_0_0_1(n196_O_12_0_0_1),
    .O_12_0_1_0(n196_O_12_0_1_0),
    .O_12_0_1_1(n196_O_12_0_1_1),
    .O_13_0_0_0(n196_O_13_0_0_0),
    .O_13_0_0_1(n196_O_13_0_0_1),
    .O_13_0_1_0(n196_O_13_0_1_0),
    .O_13_0_1_1(n196_O_13_0_1_1),
    .O_14_0_0_0(n196_O_14_0_0_0),
    .O_14_0_0_1(n196_O_14_0_0_1),
    .O_14_0_1_0(n196_O_14_0_1_0),
    .O_14_0_1_1(n196_O_14_0_1_1),
    .O_15_0_0_0(n196_O_15_0_0_0),
    .O_15_0_0_1(n196_O_15_0_0_1),
    .O_15_0_1_0(n196_O_15_0_1_0),
    .O_15_0_1_1(n196_O_15_0_1_1)
  );
  MapT_14 n203 ( // @[Top.scala 202:22]
    .valid_up(n203_valid_up),
    .valid_down(n203_valid_down),
    .I_0_0_0_0(n203_I_0_0_0_0),
    .I_0_0_0_1(n203_I_0_0_0_1),
    .I_0_0_1_0(n203_I_0_0_1_0),
    .I_0_0_1_1(n203_I_0_0_1_1),
    .I_1_0_0_0(n203_I_1_0_0_0),
    .I_1_0_0_1(n203_I_1_0_0_1),
    .I_1_0_1_0(n203_I_1_0_1_0),
    .I_1_0_1_1(n203_I_1_0_1_1),
    .I_2_0_0_0(n203_I_2_0_0_0),
    .I_2_0_0_1(n203_I_2_0_0_1),
    .I_2_0_1_0(n203_I_2_0_1_0),
    .I_2_0_1_1(n203_I_2_0_1_1),
    .I_3_0_0_0(n203_I_3_0_0_0),
    .I_3_0_0_1(n203_I_3_0_0_1),
    .I_3_0_1_0(n203_I_3_0_1_0),
    .I_3_0_1_1(n203_I_3_0_1_1),
    .I_4_0_0_0(n203_I_4_0_0_0),
    .I_4_0_0_1(n203_I_4_0_0_1),
    .I_4_0_1_0(n203_I_4_0_1_0),
    .I_4_0_1_1(n203_I_4_0_1_1),
    .I_5_0_0_0(n203_I_5_0_0_0),
    .I_5_0_0_1(n203_I_5_0_0_1),
    .I_5_0_1_0(n203_I_5_0_1_0),
    .I_5_0_1_1(n203_I_5_0_1_1),
    .I_6_0_0_0(n203_I_6_0_0_0),
    .I_6_0_0_1(n203_I_6_0_0_1),
    .I_6_0_1_0(n203_I_6_0_1_0),
    .I_6_0_1_1(n203_I_6_0_1_1),
    .I_7_0_0_0(n203_I_7_0_0_0),
    .I_7_0_0_1(n203_I_7_0_0_1),
    .I_7_0_1_0(n203_I_7_0_1_0),
    .I_7_0_1_1(n203_I_7_0_1_1),
    .I_8_0_0_0(n203_I_8_0_0_0),
    .I_8_0_0_1(n203_I_8_0_0_1),
    .I_8_0_1_0(n203_I_8_0_1_0),
    .I_8_0_1_1(n203_I_8_0_1_1),
    .I_9_0_0_0(n203_I_9_0_0_0),
    .I_9_0_0_1(n203_I_9_0_0_1),
    .I_9_0_1_0(n203_I_9_0_1_0),
    .I_9_0_1_1(n203_I_9_0_1_1),
    .I_10_0_0_0(n203_I_10_0_0_0),
    .I_10_0_0_1(n203_I_10_0_0_1),
    .I_10_0_1_0(n203_I_10_0_1_0),
    .I_10_0_1_1(n203_I_10_0_1_1),
    .I_11_0_0_0(n203_I_11_0_0_0),
    .I_11_0_0_1(n203_I_11_0_0_1),
    .I_11_0_1_0(n203_I_11_0_1_0),
    .I_11_0_1_1(n203_I_11_0_1_1),
    .I_12_0_0_0(n203_I_12_0_0_0),
    .I_12_0_0_1(n203_I_12_0_0_1),
    .I_12_0_1_0(n203_I_12_0_1_0),
    .I_12_0_1_1(n203_I_12_0_1_1),
    .I_13_0_0_0(n203_I_13_0_0_0),
    .I_13_0_0_1(n203_I_13_0_0_1),
    .I_13_0_1_0(n203_I_13_0_1_0),
    .I_13_0_1_1(n203_I_13_0_1_1),
    .I_14_0_0_0(n203_I_14_0_0_0),
    .I_14_0_0_1(n203_I_14_0_0_1),
    .I_14_0_1_0(n203_I_14_0_1_0),
    .I_14_0_1_1(n203_I_14_0_1_1),
    .I_15_0_0_0(n203_I_15_0_0_0),
    .I_15_0_0_1(n203_I_15_0_0_1),
    .I_15_0_1_0(n203_I_15_0_1_0),
    .I_15_0_1_1(n203_I_15_0_1_1),
    .O_0_0_0(n203_O_0_0_0),
    .O_0_0_1(n203_O_0_0_1),
    .O_0_1_0(n203_O_0_1_0),
    .O_0_1_1(n203_O_0_1_1),
    .O_1_0_0(n203_O_1_0_0),
    .O_1_0_1(n203_O_1_0_1),
    .O_1_1_0(n203_O_1_1_0),
    .O_1_1_1(n203_O_1_1_1),
    .O_2_0_0(n203_O_2_0_0),
    .O_2_0_1(n203_O_2_0_1),
    .O_2_1_0(n203_O_2_1_0),
    .O_2_1_1(n203_O_2_1_1),
    .O_3_0_0(n203_O_3_0_0),
    .O_3_0_1(n203_O_3_0_1),
    .O_3_1_0(n203_O_3_1_0),
    .O_3_1_1(n203_O_3_1_1),
    .O_4_0_0(n203_O_4_0_0),
    .O_4_0_1(n203_O_4_0_1),
    .O_4_1_0(n203_O_4_1_0),
    .O_4_1_1(n203_O_4_1_1),
    .O_5_0_0(n203_O_5_0_0),
    .O_5_0_1(n203_O_5_0_1),
    .O_5_1_0(n203_O_5_1_0),
    .O_5_1_1(n203_O_5_1_1),
    .O_6_0_0(n203_O_6_0_0),
    .O_6_0_1(n203_O_6_0_1),
    .O_6_1_0(n203_O_6_1_0),
    .O_6_1_1(n203_O_6_1_1),
    .O_7_0_0(n203_O_7_0_0),
    .O_7_0_1(n203_O_7_0_1),
    .O_7_1_0(n203_O_7_1_0),
    .O_7_1_1(n203_O_7_1_1),
    .O_8_0_0(n203_O_8_0_0),
    .O_8_0_1(n203_O_8_0_1),
    .O_8_1_0(n203_O_8_1_0),
    .O_8_1_1(n203_O_8_1_1),
    .O_9_0_0(n203_O_9_0_0),
    .O_9_0_1(n203_O_9_0_1),
    .O_9_1_0(n203_O_9_1_0),
    .O_9_1_1(n203_O_9_1_1),
    .O_10_0_0(n203_O_10_0_0),
    .O_10_0_1(n203_O_10_0_1),
    .O_10_1_0(n203_O_10_1_0),
    .O_10_1_1(n203_O_10_1_1),
    .O_11_0_0(n203_O_11_0_0),
    .O_11_0_1(n203_O_11_0_1),
    .O_11_1_0(n203_O_11_1_0),
    .O_11_1_1(n203_O_11_1_1),
    .O_12_0_0(n203_O_12_0_0),
    .O_12_0_1(n203_O_12_0_1),
    .O_12_1_0(n203_O_12_1_0),
    .O_12_1_1(n203_O_12_1_1),
    .O_13_0_0(n203_O_13_0_0),
    .O_13_0_1(n203_O_13_0_1),
    .O_13_1_0(n203_O_13_1_0),
    .O_13_1_1(n203_O_13_1_1),
    .O_14_0_0(n203_O_14_0_0),
    .O_14_0_1(n203_O_14_0_1),
    .O_14_1_0(n203_O_14_1_0),
    .O_14_1_1(n203_O_14_1_1),
    .O_15_0_0(n203_O_15_0_0),
    .O_15_0_1(n203_O_15_0_1),
    .O_15_1_0(n203_O_15_1_0),
    .O_15_1_1(n203_O_15_1_1)
  );
  MapT_15 n245 ( // @[Top.scala 205:22]
    .clock(n245_clock),
    .reset(n245_reset),
    .valid_up(n245_valid_up),
    .valid_down(n245_valid_down),
    .I_0_0_0(n245_I_0_0_0),
    .I_0_0_1(n245_I_0_0_1),
    .I_0_1_0(n245_I_0_1_0),
    .I_0_1_1(n245_I_0_1_1),
    .I_1_0_0(n245_I_1_0_0),
    .I_1_0_1(n245_I_1_0_1),
    .I_1_1_0(n245_I_1_1_0),
    .I_1_1_1(n245_I_1_1_1),
    .I_2_0_0(n245_I_2_0_0),
    .I_2_0_1(n245_I_2_0_1),
    .I_2_1_0(n245_I_2_1_0),
    .I_2_1_1(n245_I_2_1_1),
    .I_3_0_0(n245_I_3_0_0),
    .I_3_0_1(n245_I_3_0_1),
    .I_3_1_0(n245_I_3_1_0),
    .I_3_1_1(n245_I_3_1_1),
    .I_4_0_0(n245_I_4_0_0),
    .I_4_0_1(n245_I_4_0_1),
    .I_4_1_0(n245_I_4_1_0),
    .I_4_1_1(n245_I_4_1_1),
    .I_5_0_0(n245_I_5_0_0),
    .I_5_0_1(n245_I_5_0_1),
    .I_5_1_0(n245_I_5_1_0),
    .I_5_1_1(n245_I_5_1_1),
    .I_6_0_0(n245_I_6_0_0),
    .I_6_0_1(n245_I_6_0_1),
    .I_6_1_0(n245_I_6_1_0),
    .I_6_1_1(n245_I_6_1_1),
    .I_7_0_0(n245_I_7_0_0),
    .I_7_0_1(n245_I_7_0_1),
    .I_7_1_0(n245_I_7_1_0),
    .I_7_1_1(n245_I_7_1_1),
    .I_8_0_0(n245_I_8_0_0),
    .I_8_0_1(n245_I_8_0_1),
    .I_8_1_0(n245_I_8_1_0),
    .I_8_1_1(n245_I_8_1_1),
    .I_9_0_0(n245_I_9_0_0),
    .I_9_0_1(n245_I_9_0_1),
    .I_9_1_0(n245_I_9_1_0),
    .I_9_1_1(n245_I_9_1_1),
    .I_10_0_0(n245_I_10_0_0),
    .I_10_0_1(n245_I_10_0_1),
    .I_10_1_0(n245_I_10_1_0),
    .I_10_1_1(n245_I_10_1_1),
    .I_11_0_0(n245_I_11_0_0),
    .I_11_0_1(n245_I_11_0_1),
    .I_11_1_0(n245_I_11_1_0),
    .I_11_1_1(n245_I_11_1_1),
    .I_12_0_0(n245_I_12_0_0),
    .I_12_0_1(n245_I_12_0_1),
    .I_12_1_0(n245_I_12_1_0),
    .I_12_1_1(n245_I_12_1_1),
    .I_13_0_0(n245_I_13_0_0),
    .I_13_0_1(n245_I_13_0_1),
    .I_13_1_0(n245_I_13_1_0),
    .I_13_1_1(n245_I_13_1_1),
    .I_14_0_0(n245_I_14_0_0),
    .I_14_0_1(n245_I_14_0_1),
    .I_14_1_0(n245_I_14_1_0),
    .I_14_1_1(n245_I_14_1_1),
    .I_15_0_0(n245_I_15_0_0),
    .I_15_0_1(n245_I_15_0_1),
    .I_15_1_0(n245_I_15_1_0),
    .I_15_1_1(n245_I_15_1_1),
    .O_0_0_0(n245_O_0_0_0),
    .O_1_0_0(n245_O_1_0_0),
    .O_2_0_0(n245_O_2_0_0),
    .O_3_0_0(n245_O_3_0_0),
    .O_4_0_0(n245_O_4_0_0),
    .O_5_0_0(n245_O_5_0_0),
    .O_6_0_0(n245_O_6_0_0),
    .O_7_0_0(n245_O_7_0_0),
    .O_8_0_0(n245_O_8_0_0),
    .O_9_0_0(n245_O_9_0_0),
    .O_10_0_0(n245_O_10_0_0),
    .O_11_0_0(n245_O_11_0_0),
    .O_12_0_0(n245_O_12_0_0),
    .O_13_0_0(n245_O_13_0_0),
    .O_14_0_0(n245_O_14_0_0),
    .O_15_0_0(n245_O_15_0_0)
  );
  Passthrough n246 ( // @[Top.scala 208:22]
    .valid_up(n246_valid_up),
    .valid_down(n246_valid_down),
    .I_0_0_0(n246_I_0_0_0),
    .I_1_0_0(n246_I_1_0_0),
    .I_2_0_0(n246_I_2_0_0),
    .I_3_0_0(n246_I_3_0_0),
    .I_4_0_0(n246_I_4_0_0),
    .I_5_0_0(n246_I_5_0_0),
    .I_6_0_0(n246_I_6_0_0),
    .I_7_0_0(n246_I_7_0_0),
    .I_8_0_0(n246_I_8_0_0),
    .I_9_0_0(n246_I_9_0_0),
    .I_10_0_0(n246_I_10_0_0),
    .I_11_0_0(n246_I_11_0_0),
    .I_12_0_0(n246_I_12_0_0),
    .I_13_0_0(n246_I_13_0_0),
    .I_14_0_0(n246_I_14_0_0),
    .I_15_0_0(n246_I_15_0_0),
    .O_0_0(n246_O_0_0),
    .O_1_0(n246_O_1_0),
    .O_2_0(n246_O_2_0),
    .O_3_0(n246_O_3_0),
    .O_4_0(n246_O_4_0),
    .O_5_0(n246_O_5_0),
    .O_6_0(n246_O_6_0),
    .O_7_0(n246_O_7_0),
    .O_8_0(n246_O_8_0),
    .O_9_0(n246_O_9_0),
    .O_10_0(n246_O_10_0),
    .O_11_0(n246_O_11_0),
    .O_12_0(n246_O_12_0),
    .O_13_0(n246_O_13_0),
    .O_14_0(n246_O_14_0),
    .O_15_0(n246_O_15_0)
  );
  Passthrough_1 n247 ( // @[Top.scala 211:22]
    .valid_up(n247_valid_up),
    .valid_down(n247_valid_down),
    .I_0_0(n247_I_0_0),
    .I_1_0(n247_I_1_0),
    .I_2_0(n247_I_2_0),
    .I_3_0(n247_I_3_0),
    .I_4_0(n247_I_4_0),
    .I_5_0(n247_I_5_0),
    .I_6_0(n247_I_6_0),
    .I_7_0(n247_I_7_0),
    .I_8_0(n247_I_8_0),
    .I_9_0(n247_I_9_0),
    .I_10_0(n247_I_10_0),
    .I_11_0(n247_I_11_0),
    .I_12_0(n247_I_12_0),
    .I_13_0(n247_I_13_0),
    .I_14_0(n247_I_14_0),
    .I_15_0(n247_I_15_0),
    .O_0(n247_O_0),
    .O_1(n247_O_1),
    .O_2(n247_O_2),
    .O_3(n247_O_3),
    .O_4(n247_O_4),
    .O_5(n247_O_5),
    .O_6(n247_O_6),
    .O_7(n247_O_7),
    .O_8(n247_O_8),
    .O_9(n247_O_9),
    .O_10(n247_O_10),
    .O_11(n247_O_11),
    .O_12(n247_O_12),
    .O_13(n247_O_13),
    .O_14(n247_O_14),
    .O_15(n247_O_15)
  );
  FIFO n248 ( // @[Top.scala 214:22]
    .clock(n248_clock),
    .reset(n248_reset),
    .valid_up(n248_valid_up),
    .valid_down(n248_valid_down),
    .I_0(n248_I_0),
    .I_1(n248_I_1),
    .I_2(n248_I_2),
    .I_3(n248_I_3),
    .I_4(n248_I_4),
    .I_5(n248_I_5),
    .I_6(n248_I_6),
    .I_7(n248_I_7),
    .I_8(n248_I_8),
    .I_9(n248_I_9),
    .I_10(n248_I_10),
    .I_11(n248_I_11),
    .I_12(n248_I_12),
    .I_13(n248_I_13),
    .I_14(n248_I_14),
    .I_15(n248_I_15),
    .O_0(n248_O_0),
    .O_1(n248_O_1),
    .O_2(n248_O_2),
    .O_3(n248_O_3),
    .O_4(n248_O_4),
    .O_5(n248_O_5),
    .O_6(n248_O_6),
    .O_7(n248_O_7),
    .O_8(n248_O_8),
    .O_9(n248_O_9),
    .O_10(n248_O_10),
    .O_11(n248_O_11),
    .O_12(n248_O_12),
    .O_13(n248_O_13),
    .O_14(n248_O_14),
    .O_15(n248_O_15)
  );
  FIFO n249 ( // @[Top.scala 217:22]
    .clock(n249_clock),
    .reset(n249_reset),
    .valid_up(n249_valid_up),
    .valid_down(n249_valid_down),
    .I_0(n249_I_0),
    .I_1(n249_I_1),
    .I_2(n249_I_2),
    .I_3(n249_I_3),
    .I_4(n249_I_4),
    .I_5(n249_I_5),
    .I_6(n249_I_6),
    .I_7(n249_I_7),
    .I_8(n249_I_8),
    .I_9(n249_I_9),
    .I_10(n249_I_10),
    .I_11(n249_I_11),
    .I_12(n249_I_12),
    .I_13(n249_I_13),
    .I_14(n249_I_14),
    .I_15(n249_I_15),
    .O_0(n249_O_0),
    .O_1(n249_O_1),
    .O_2(n249_O_2),
    .O_3(n249_O_3),
    .O_4(n249_O_4),
    .O_5(n249_O_5),
    .O_6(n249_O_6),
    .O_7(n249_O_7),
    .O_8(n249_O_8),
    .O_9(n249_O_9),
    .O_10(n249_O_10),
    .O_11(n249_O_11),
    .O_12(n249_O_12),
    .O_13(n249_O_13),
    .O_14(n249_O_14),
    .O_15(n249_O_15)
  );
  FIFO n250 ( // @[Top.scala 220:22]
    .clock(n250_clock),
    .reset(n250_reset),
    .valid_up(n250_valid_up),
    .valid_down(n250_valid_down),
    .I_0(n250_I_0),
    .I_1(n250_I_1),
    .I_2(n250_I_2),
    .I_3(n250_I_3),
    .I_4(n250_I_4),
    .I_5(n250_I_5),
    .I_6(n250_I_6),
    .I_7(n250_I_7),
    .I_8(n250_I_8),
    .I_9(n250_I_9),
    .I_10(n250_I_10),
    .I_11(n250_I_11),
    .I_12(n250_I_12),
    .I_13(n250_I_13),
    .I_14(n250_I_14),
    .I_15(n250_I_15),
    .O_0(n250_O_0),
    .O_1(n250_O_1),
    .O_2(n250_O_2),
    .O_3(n250_O_3),
    .O_4(n250_O_4),
    .O_5(n250_O_5),
    .O_6(n250_O_6),
    .O_7(n250_O_7),
    .O_8(n250_O_8),
    .O_9(n250_O_9),
    .O_10(n250_O_10),
    .O_11(n250_O_11),
    .O_12(n250_O_12),
    .O_13(n250_O_13),
    .O_14(n250_O_14),
    .O_15(n250_O_15)
  );
  assign valid_down = n250_valid_down; // @[Top.scala 224:16]
  assign O_0 = n250_O_0; // @[Top.scala 223:7]
  assign O_1 = n250_O_1; // @[Top.scala 223:7]
  assign O_2 = n250_O_2; // @[Top.scala 223:7]
  assign O_3 = n250_O_3; // @[Top.scala 223:7]
  assign O_4 = n250_O_4; // @[Top.scala 223:7]
  assign O_5 = n250_O_5; // @[Top.scala 223:7]
  assign O_6 = n250_O_6; // @[Top.scala 223:7]
  assign O_7 = n250_O_7; // @[Top.scala 223:7]
  assign O_8 = n250_O_8; // @[Top.scala 223:7]
  assign O_9 = n250_O_9; // @[Top.scala 223:7]
  assign O_10 = n250_O_10; // @[Top.scala 223:7]
  assign O_11 = n250_O_11; // @[Top.scala 223:7]
  assign O_12 = n250_O_12; // @[Top.scala 223:7]
  assign O_13 = n250_O_13; // @[Top.scala 223:7]
  assign O_14 = n250_O_14; // @[Top.scala 223:7]
  assign O_15 = n250_O_15; // @[Top.scala 223:7]
  assign n1_clock = clock;
  assign n1_reset = reset;
  assign n1_valid_up = valid_up; // @[Top.scala 76:17]
  assign n1_I_0 = I_0; // @[Top.scala 75:10]
  assign n1_I_1 = I_1; // @[Top.scala 75:10]
  assign n1_I_2 = I_2; // @[Top.scala 75:10]
  assign n1_I_3 = I_3; // @[Top.scala 75:10]
  assign n1_I_4 = I_4; // @[Top.scala 75:10]
  assign n1_I_5 = I_5; // @[Top.scala 75:10]
  assign n1_I_6 = I_6; // @[Top.scala 75:10]
  assign n1_I_7 = I_7; // @[Top.scala 75:10]
  assign n1_I_8 = I_8; // @[Top.scala 75:10]
  assign n1_I_9 = I_9; // @[Top.scala 75:10]
  assign n1_I_10 = I_10; // @[Top.scala 75:10]
  assign n1_I_11 = I_11; // @[Top.scala 75:10]
  assign n1_I_12 = I_12; // @[Top.scala 75:10]
  assign n1_I_13 = I_13; // @[Top.scala 75:10]
  assign n1_I_14 = I_14; // @[Top.scala 75:10]
  assign n1_I_15 = I_15; // @[Top.scala 75:10]
  assign n2_clock = clock;
  assign n2_reset = reset;
  assign n2_valid_up = n1_valid_down; // @[Top.scala 79:17]
  assign n2_I_0 = n1_O_0; // @[Top.scala 78:10]
  assign n2_I_1 = n1_O_1; // @[Top.scala 78:10]
  assign n2_I_2 = n1_O_2; // @[Top.scala 78:10]
  assign n2_I_3 = n1_O_3; // @[Top.scala 78:10]
  assign n2_I_4 = n1_O_4; // @[Top.scala 78:10]
  assign n2_I_5 = n1_O_5; // @[Top.scala 78:10]
  assign n2_I_6 = n1_O_6; // @[Top.scala 78:10]
  assign n2_I_7 = n1_O_7; // @[Top.scala 78:10]
  assign n2_I_8 = n1_O_8; // @[Top.scala 78:10]
  assign n2_I_9 = n1_O_9; // @[Top.scala 78:10]
  assign n2_I_10 = n1_O_10; // @[Top.scala 78:10]
  assign n2_I_11 = n1_O_11; // @[Top.scala 78:10]
  assign n2_I_12 = n1_O_12; // @[Top.scala 78:10]
  assign n2_I_13 = n1_O_13; // @[Top.scala 78:10]
  assign n2_I_14 = n1_O_14; // @[Top.scala 78:10]
  assign n2_I_15 = n1_O_15; // @[Top.scala 78:10]
  assign n3_clock = clock;
  assign n3_reset = reset;
  assign n3_valid_up = n2_valid_down; // @[Top.scala 82:17]
  assign n3_I_0 = n2_O_0; // @[Top.scala 81:10]
  assign n3_I_1 = n2_O_1; // @[Top.scala 81:10]
  assign n3_I_2 = n2_O_2; // @[Top.scala 81:10]
  assign n3_I_3 = n2_O_3; // @[Top.scala 81:10]
  assign n3_I_4 = n2_O_4; // @[Top.scala 81:10]
  assign n3_I_5 = n2_O_5; // @[Top.scala 81:10]
  assign n3_I_6 = n2_O_6; // @[Top.scala 81:10]
  assign n3_I_7 = n2_O_7; // @[Top.scala 81:10]
  assign n3_I_8 = n2_O_8; // @[Top.scala 81:10]
  assign n3_I_9 = n2_O_9; // @[Top.scala 81:10]
  assign n3_I_10 = n2_O_10; // @[Top.scala 81:10]
  assign n3_I_11 = n2_O_11; // @[Top.scala 81:10]
  assign n3_I_12 = n2_O_12; // @[Top.scala 81:10]
  assign n3_I_13 = n2_O_13; // @[Top.scala 81:10]
  assign n3_I_14 = n2_O_14; // @[Top.scala 81:10]
  assign n3_I_15 = n2_O_15; // @[Top.scala 81:10]
  assign n4_clock = clock;
  assign n4_valid_up = n3_valid_down; // @[Top.scala 85:17]
  assign n4_I_0 = n3_O_0; // @[Top.scala 84:10]
  assign n4_I_1 = n3_O_1; // @[Top.scala 84:10]
  assign n4_I_2 = n3_O_2; // @[Top.scala 84:10]
  assign n4_I_3 = n3_O_3; // @[Top.scala 84:10]
  assign n4_I_4 = n3_O_4; // @[Top.scala 84:10]
  assign n4_I_5 = n3_O_5; // @[Top.scala 84:10]
  assign n4_I_6 = n3_O_6; // @[Top.scala 84:10]
  assign n4_I_7 = n3_O_7; // @[Top.scala 84:10]
  assign n4_I_8 = n3_O_8; // @[Top.scala 84:10]
  assign n4_I_9 = n3_O_9; // @[Top.scala 84:10]
  assign n4_I_10 = n3_O_10; // @[Top.scala 84:10]
  assign n4_I_11 = n3_O_11; // @[Top.scala 84:10]
  assign n4_I_12 = n3_O_12; // @[Top.scala 84:10]
  assign n4_I_13 = n3_O_13; // @[Top.scala 84:10]
  assign n4_I_14 = n3_O_14; // @[Top.scala 84:10]
  assign n4_I_15 = n3_O_15; // @[Top.scala 84:10]
  assign n5_clock = clock;
  assign n5_valid_up = n4_valid_down; // @[Top.scala 88:17]
  assign n5_I_0 = n4_O_0; // @[Top.scala 87:10]
  assign n5_I_1 = n4_O_1; // @[Top.scala 87:10]
  assign n5_I_2 = n4_O_2; // @[Top.scala 87:10]
  assign n5_I_3 = n4_O_3; // @[Top.scala 87:10]
  assign n5_I_4 = n4_O_4; // @[Top.scala 87:10]
  assign n5_I_5 = n4_O_5; // @[Top.scala 87:10]
  assign n5_I_6 = n4_O_6; // @[Top.scala 87:10]
  assign n5_I_7 = n4_O_7; // @[Top.scala 87:10]
  assign n5_I_8 = n4_O_8; // @[Top.scala 87:10]
  assign n5_I_9 = n4_O_9; // @[Top.scala 87:10]
  assign n5_I_10 = n4_O_10; // @[Top.scala 87:10]
  assign n5_I_11 = n4_O_11; // @[Top.scala 87:10]
  assign n5_I_12 = n4_O_12; // @[Top.scala 87:10]
  assign n5_I_13 = n4_O_13; // @[Top.scala 87:10]
  assign n5_I_14 = n4_O_14; // @[Top.scala 87:10]
  assign n5_I_15 = n4_O_15; // @[Top.scala 87:10]
  assign n6_valid_up = n5_valid_down & n4_valid_down; // @[Top.scala 92:17]
  assign n6_I0_0 = n5_O_0; // @[Top.scala 90:11]
  assign n6_I0_1 = n5_O_1; // @[Top.scala 90:11]
  assign n6_I0_2 = n5_O_2; // @[Top.scala 90:11]
  assign n6_I0_3 = n5_O_3; // @[Top.scala 90:11]
  assign n6_I0_4 = n5_O_4; // @[Top.scala 90:11]
  assign n6_I0_5 = n5_O_5; // @[Top.scala 90:11]
  assign n6_I0_6 = n5_O_6; // @[Top.scala 90:11]
  assign n6_I0_7 = n5_O_7; // @[Top.scala 90:11]
  assign n6_I0_8 = n5_O_8; // @[Top.scala 90:11]
  assign n6_I0_9 = n5_O_9; // @[Top.scala 90:11]
  assign n6_I0_10 = n5_O_10; // @[Top.scala 90:11]
  assign n6_I0_11 = n5_O_11; // @[Top.scala 90:11]
  assign n6_I0_12 = n5_O_12; // @[Top.scala 90:11]
  assign n6_I0_13 = n5_O_13; // @[Top.scala 90:11]
  assign n6_I0_14 = n5_O_14; // @[Top.scala 90:11]
  assign n6_I0_15 = n5_O_15; // @[Top.scala 90:11]
  assign n6_I1_0 = n4_O_0; // @[Top.scala 91:11]
  assign n6_I1_1 = n4_O_1; // @[Top.scala 91:11]
  assign n6_I1_2 = n4_O_2; // @[Top.scala 91:11]
  assign n6_I1_3 = n4_O_3; // @[Top.scala 91:11]
  assign n6_I1_4 = n4_O_4; // @[Top.scala 91:11]
  assign n6_I1_5 = n4_O_5; // @[Top.scala 91:11]
  assign n6_I1_6 = n4_O_6; // @[Top.scala 91:11]
  assign n6_I1_7 = n4_O_7; // @[Top.scala 91:11]
  assign n6_I1_8 = n4_O_8; // @[Top.scala 91:11]
  assign n6_I1_9 = n4_O_9; // @[Top.scala 91:11]
  assign n6_I1_10 = n4_O_10; // @[Top.scala 91:11]
  assign n6_I1_11 = n4_O_11; // @[Top.scala 91:11]
  assign n6_I1_12 = n4_O_12; // @[Top.scala 91:11]
  assign n6_I1_13 = n4_O_13; // @[Top.scala 91:11]
  assign n6_I1_14 = n4_O_14; // @[Top.scala 91:11]
  assign n6_I1_15 = n4_O_15; // @[Top.scala 91:11]
  assign n13_valid_up = n6_valid_down & n3_valid_down; // @[Top.scala 96:18]
  assign n13_I0_0_0 = n6_O_0_0; // @[Top.scala 94:12]
  assign n13_I0_0_1 = n6_O_0_1; // @[Top.scala 94:12]
  assign n13_I0_1_0 = n6_O_1_0; // @[Top.scala 94:12]
  assign n13_I0_1_1 = n6_O_1_1; // @[Top.scala 94:12]
  assign n13_I0_2_0 = n6_O_2_0; // @[Top.scala 94:12]
  assign n13_I0_2_1 = n6_O_2_1; // @[Top.scala 94:12]
  assign n13_I0_3_0 = n6_O_3_0; // @[Top.scala 94:12]
  assign n13_I0_3_1 = n6_O_3_1; // @[Top.scala 94:12]
  assign n13_I0_4_0 = n6_O_4_0; // @[Top.scala 94:12]
  assign n13_I0_4_1 = n6_O_4_1; // @[Top.scala 94:12]
  assign n13_I0_5_0 = n6_O_5_0; // @[Top.scala 94:12]
  assign n13_I0_5_1 = n6_O_5_1; // @[Top.scala 94:12]
  assign n13_I0_6_0 = n6_O_6_0; // @[Top.scala 94:12]
  assign n13_I0_6_1 = n6_O_6_1; // @[Top.scala 94:12]
  assign n13_I0_7_0 = n6_O_7_0; // @[Top.scala 94:12]
  assign n13_I0_7_1 = n6_O_7_1; // @[Top.scala 94:12]
  assign n13_I0_8_0 = n6_O_8_0; // @[Top.scala 94:12]
  assign n13_I0_8_1 = n6_O_8_1; // @[Top.scala 94:12]
  assign n13_I0_9_0 = n6_O_9_0; // @[Top.scala 94:12]
  assign n13_I0_9_1 = n6_O_9_1; // @[Top.scala 94:12]
  assign n13_I0_10_0 = n6_O_10_0; // @[Top.scala 94:12]
  assign n13_I0_10_1 = n6_O_10_1; // @[Top.scala 94:12]
  assign n13_I0_11_0 = n6_O_11_0; // @[Top.scala 94:12]
  assign n13_I0_11_1 = n6_O_11_1; // @[Top.scala 94:12]
  assign n13_I0_12_0 = n6_O_12_0; // @[Top.scala 94:12]
  assign n13_I0_12_1 = n6_O_12_1; // @[Top.scala 94:12]
  assign n13_I0_13_0 = n6_O_13_0; // @[Top.scala 94:12]
  assign n13_I0_13_1 = n6_O_13_1; // @[Top.scala 94:12]
  assign n13_I0_14_0 = n6_O_14_0; // @[Top.scala 94:12]
  assign n13_I0_14_1 = n6_O_14_1; // @[Top.scala 94:12]
  assign n13_I0_15_0 = n6_O_15_0; // @[Top.scala 94:12]
  assign n13_I0_15_1 = n6_O_15_1; // @[Top.scala 94:12]
  assign n13_I1_0 = n3_O_0; // @[Top.scala 95:12]
  assign n13_I1_1 = n3_O_1; // @[Top.scala 95:12]
  assign n13_I1_2 = n3_O_2; // @[Top.scala 95:12]
  assign n13_I1_3 = n3_O_3; // @[Top.scala 95:12]
  assign n13_I1_4 = n3_O_4; // @[Top.scala 95:12]
  assign n13_I1_5 = n3_O_5; // @[Top.scala 95:12]
  assign n13_I1_6 = n3_O_6; // @[Top.scala 95:12]
  assign n13_I1_7 = n3_O_7; // @[Top.scala 95:12]
  assign n13_I1_8 = n3_O_8; // @[Top.scala 95:12]
  assign n13_I1_9 = n3_O_9; // @[Top.scala 95:12]
  assign n13_I1_10 = n3_O_10; // @[Top.scala 95:12]
  assign n13_I1_11 = n3_O_11; // @[Top.scala 95:12]
  assign n13_I1_12 = n3_O_12; // @[Top.scala 95:12]
  assign n13_I1_13 = n3_O_13; // @[Top.scala 95:12]
  assign n13_I1_14 = n3_O_14; // @[Top.scala 95:12]
  assign n13_I1_15 = n3_O_15; // @[Top.scala 95:12]
  assign n22_valid_up = n13_valid_down; // @[Top.scala 99:18]
  assign n22_I_0_0 = n13_O_0_0; // @[Top.scala 98:11]
  assign n22_I_0_1 = n13_O_0_1; // @[Top.scala 98:11]
  assign n22_I_0_2 = n13_O_0_2; // @[Top.scala 98:11]
  assign n22_I_1_0 = n13_O_1_0; // @[Top.scala 98:11]
  assign n22_I_1_1 = n13_O_1_1; // @[Top.scala 98:11]
  assign n22_I_1_2 = n13_O_1_2; // @[Top.scala 98:11]
  assign n22_I_2_0 = n13_O_2_0; // @[Top.scala 98:11]
  assign n22_I_2_1 = n13_O_2_1; // @[Top.scala 98:11]
  assign n22_I_2_2 = n13_O_2_2; // @[Top.scala 98:11]
  assign n22_I_3_0 = n13_O_3_0; // @[Top.scala 98:11]
  assign n22_I_3_1 = n13_O_3_1; // @[Top.scala 98:11]
  assign n22_I_3_2 = n13_O_3_2; // @[Top.scala 98:11]
  assign n22_I_4_0 = n13_O_4_0; // @[Top.scala 98:11]
  assign n22_I_4_1 = n13_O_4_1; // @[Top.scala 98:11]
  assign n22_I_4_2 = n13_O_4_2; // @[Top.scala 98:11]
  assign n22_I_5_0 = n13_O_5_0; // @[Top.scala 98:11]
  assign n22_I_5_1 = n13_O_5_1; // @[Top.scala 98:11]
  assign n22_I_5_2 = n13_O_5_2; // @[Top.scala 98:11]
  assign n22_I_6_0 = n13_O_6_0; // @[Top.scala 98:11]
  assign n22_I_6_1 = n13_O_6_1; // @[Top.scala 98:11]
  assign n22_I_6_2 = n13_O_6_2; // @[Top.scala 98:11]
  assign n22_I_7_0 = n13_O_7_0; // @[Top.scala 98:11]
  assign n22_I_7_1 = n13_O_7_1; // @[Top.scala 98:11]
  assign n22_I_7_2 = n13_O_7_2; // @[Top.scala 98:11]
  assign n22_I_8_0 = n13_O_8_0; // @[Top.scala 98:11]
  assign n22_I_8_1 = n13_O_8_1; // @[Top.scala 98:11]
  assign n22_I_8_2 = n13_O_8_2; // @[Top.scala 98:11]
  assign n22_I_9_0 = n13_O_9_0; // @[Top.scala 98:11]
  assign n22_I_9_1 = n13_O_9_1; // @[Top.scala 98:11]
  assign n22_I_9_2 = n13_O_9_2; // @[Top.scala 98:11]
  assign n22_I_10_0 = n13_O_10_0; // @[Top.scala 98:11]
  assign n22_I_10_1 = n13_O_10_1; // @[Top.scala 98:11]
  assign n22_I_10_2 = n13_O_10_2; // @[Top.scala 98:11]
  assign n22_I_11_0 = n13_O_11_0; // @[Top.scala 98:11]
  assign n22_I_11_1 = n13_O_11_1; // @[Top.scala 98:11]
  assign n22_I_11_2 = n13_O_11_2; // @[Top.scala 98:11]
  assign n22_I_12_0 = n13_O_12_0; // @[Top.scala 98:11]
  assign n22_I_12_1 = n13_O_12_1; // @[Top.scala 98:11]
  assign n22_I_12_2 = n13_O_12_2; // @[Top.scala 98:11]
  assign n22_I_13_0 = n13_O_13_0; // @[Top.scala 98:11]
  assign n22_I_13_1 = n13_O_13_1; // @[Top.scala 98:11]
  assign n22_I_13_2 = n13_O_13_2; // @[Top.scala 98:11]
  assign n22_I_14_0 = n13_O_14_0; // @[Top.scala 98:11]
  assign n22_I_14_1 = n13_O_14_1; // @[Top.scala 98:11]
  assign n22_I_14_2 = n13_O_14_2; // @[Top.scala 98:11]
  assign n22_I_15_0 = n13_O_15_0; // @[Top.scala 98:11]
  assign n22_I_15_1 = n13_O_15_1; // @[Top.scala 98:11]
  assign n22_I_15_2 = n13_O_15_2; // @[Top.scala 98:11]
  assign n29_valid_up = n22_valid_down; // @[Top.scala 102:18]
  assign n29_I_0_0_0 = n22_O_0_0_0; // @[Top.scala 101:11]
  assign n29_I_0_0_1 = n22_O_0_0_1; // @[Top.scala 101:11]
  assign n29_I_0_0_2 = n22_O_0_0_2; // @[Top.scala 101:11]
  assign n29_I_1_0_0 = n22_O_1_0_0; // @[Top.scala 101:11]
  assign n29_I_1_0_1 = n22_O_1_0_1; // @[Top.scala 101:11]
  assign n29_I_1_0_2 = n22_O_1_0_2; // @[Top.scala 101:11]
  assign n29_I_2_0_0 = n22_O_2_0_0; // @[Top.scala 101:11]
  assign n29_I_2_0_1 = n22_O_2_0_1; // @[Top.scala 101:11]
  assign n29_I_2_0_2 = n22_O_2_0_2; // @[Top.scala 101:11]
  assign n29_I_3_0_0 = n22_O_3_0_0; // @[Top.scala 101:11]
  assign n29_I_3_0_1 = n22_O_3_0_1; // @[Top.scala 101:11]
  assign n29_I_3_0_2 = n22_O_3_0_2; // @[Top.scala 101:11]
  assign n29_I_4_0_0 = n22_O_4_0_0; // @[Top.scala 101:11]
  assign n29_I_4_0_1 = n22_O_4_0_1; // @[Top.scala 101:11]
  assign n29_I_4_0_2 = n22_O_4_0_2; // @[Top.scala 101:11]
  assign n29_I_5_0_0 = n22_O_5_0_0; // @[Top.scala 101:11]
  assign n29_I_5_0_1 = n22_O_5_0_1; // @[Top.scala 101:11]
  assign n29_I_5_0_2 = n22_O_5_0_2; // @[Top.scala 101:11]
  assign n29_I_6_0_0 = n22_O_6_0_0; // @[Top.scala 101:11]
  assign n29_I_6_0_1 = n22_O_6_0_1; // @[Top.scala 101:11]
  assign n29_I_6_0_2 = n22_O_6_0_2; // @[Top.scala 101:11]
  assign n29_I_7_0_0 = n22_O_7_0_0; // @[Top.scala 101:11]
  assign n29_I_7_0_1 = n22_O_7_0_1; // @[Top.scala 101:11]
  assign n29_I_7_0_2 = n22_O_7_0_2; // @[Top.scala 101:11]
  assign n29_I_8_0_0 = n22_O_8_0_0; // @[Top.scala 101:11]
  assign n29_I_8_0_1 = n22_O_8_0_1; // @[Top.scala 101:11]
  assign n29_I_8_0_2 = n22_O_8_0_2; // @[Top.scala 101:11]
  assign n29_I_9_0_0 = n22_O_9_0_0; // @[Top.scala 101:11]
  assign n29_I_9_0_1 = n22_O_9_0_1; // @[Top.scala 101:11]
  assign n29_I_9_0_2 = n22_O_9_0_2; // @[Top.scala 101:11]
  assign n29_I_10_0_0 = n22_O_10_0_0; // @[Top.scala 101:11]
  assign n29_I_10_0_1 = n22_O_10_0_1; // @[Top.scala 101:11]
  assign n29_I_10_0_2 = n22_O_10_0_2; // @[Top.scala 101:11]
  assign n29_I_11_0_0 = n22_O_11_0_0; // @[Top.scala 101:11]
  assign n29_I_11_0_1 = n22_O_11_0_1; // @[Top.scala 101:11]
  assign n29_I_11_0_2 = n22_O_11_0_2; // @[Top.scala 101:11]
  assign n29_I_12_0_0 = n22_O_12_0_0; // @[Top.scala 101:11]
  assign n29_I_12_0_1 = n22_O_12_0_1; // @[Top.scala 101:11]
  assign n29_I_12_0_2 = n22_O_12_0_2; // @[Top.scala 101:11]
  assign n29_I_13_0_0 = n22_O_13_0_0; // @[Top.scala 101:11]
  assign n29_I_13_0_1 = n22_O_13_0_1; // @[Top.scala 101:11]
  assign n29_I_13_0_2 = n22_O_13_0_2; // @[Top.scala 101:11]
  assign n29_I_14_0_0 = n22_O_14_0_0; // @[Top.scala 101:11]
  assign n29_I_14_0_1 = n22_O_14_0_1; // @[Top.scala 101:11]
  assign n29_I_14_0_2 = n22_O_14_0_2; // @[Top.scala 101:11]
  assign n29_I_15_0_0 = n22_O_15_0_0; // @[Top.scala 101:11]
  assign n29_I_15_0_1 = n22_O_15_0_1; // @[Top.scala 101:11]
  assign n29_I_15_0_2 = n22_O_15_0_2; // @[Top.scala 101:11]
  assign n30_clock = clock;
  assign n30_valid_up = n2_valid_down; // @[Top.scala 105:18]
  assign n30_I_0 = n2_O_0; // @[Top.scala 104:11]
  assign n30_I_1 = n2_O_1; // @[Top.scala 104:11]
  assign n30_I_2 = n2_O_2; // @[Top.scala 104:11]
  assign n30_I_3 = n2_O_3; // @[Top.scala 104:11]
  assign n30_I_4 = n2_O_4; // @[Top.scala 104:11]
  assign n30_I_5 = n2_O_5; // @[Top.scala 104:11]
  assign n30_I_6 = n2_O_6; // @[Top.scala 104:11]
  assign n30_I_7 = n2_O_7; // @[Top.scala 104:11]
  assign n30_I_8 = n2_O_8; // @[Top.scala 104:11]
  assign n30_I_9 = n2_O_9; // @[Top.scala 104:11]
  assign n30_I_10 = n2_O_10; // @[Top.scala 104:11]
  assign n30_I_11 = n2_O_11; // @[Top.scala 104:11]
  assign n30_I_12 = n2_O_12; // @[Top.scala 104:11]
  assign n30_I_13 = n2_O_13; // @[Top.scala 104:11]
  assign n30_I_14 = n2_O_14; // @[Top.scala 104:11]
  assign n30_I_15 = n2_O_15; // @[Top.scala 104:11]
  assign n31_clock = clock;
  assign n31_valid_up = n30_valid_down; // @[Top.scala 108:18]
  assign n31_I_0 = n30_O_0; // @[Top.scala 107:11]
  assign n31_I_1 = n30_O_1; // @[Top.scala 107:11]
  assign n31_I_2 = n30_O_2; // @[Top.scala 107:11]
  assign n31_I_3 = n30_O_3; // @[Top.scala 107:11]
  assign n31_I_4 = n30_O_4; // @[Top.scala 107:11]
  assign n31_I_5 = n30_O_5; // @[Top.scala 107:11]
  assign n31_I_6 = n30_O_6; // @[Top.scala 107:11]
  assign n31_I_7 = n30_O_7; // @[Top.scala 107:11]
  assign n31_I_8 = n30_O_8; // @[Top.scala 107:11]
  assign n31_I_9 = n30_O_9; // @[Top.scala 107:11]
  assign n31_I_10 = n30_O_10; // @[Top.scala 107:11]
  assign n31_I_11 = n30_O_11; // @[Top.scala 107:11]
  assign n31_I_12 = n30_O_12; // @[Top.scala 107:11]
  assign n31_I_13 = n30_O_13; // @[Top.scala 107:11]
  assign n31_I_14 = n30_O_14; // @[Top.scala 107:11]
  assign n31_I_15 = n30_O_15; // @[Top.scala 107:11]
  assign n32_valid_up = n31_valid_down & n30_valid_down; // @[Top.scala 112:18]
  assign n32_I0_0 = n31_O_0; // @[Top.scala 110:12]
  assign n32_I0_1 = n31_O_1; // @[Top.scala 110:12]
  assign n32_I0_2 = n31_O_2; // @[Top.scala 110:12]
  assign n32_I0_3 = n31_O_3; // @[Top.scala 110:12]
  assign n32_I0_4 = n31_O_4; // @[Top.scala 110:12]
  assign n32_I0_5 = n31_O_5; // @[Top.scala 110:12]
  assign n32_I0_6 = n31_O_6; // @[Top.scala 110:12]
  assign n32_I0_7 = n31_O_7; // @[Top.scala 110:12]
  assign n32_I0_8 = n31_O_8; // @[Top.scala 110:12]
  assign n32_I0_9 = n31_O_9; // @[Top.scala 110:12]
  assign n32_I0_10 = n31_O_10; // @[Top.scala 110:12]
  assign n32_I0_11 = n31_O_11; // @[Top.scala 110:12]
  assign n32_I0_12 = n31_O_12; // @[Top.scala 110:12]
  assign n32_I0_13 = n31_O_13; // @[Top.scala 110:12]
  assign n32_I0_14 = n31_O_14; // @[Top.scala 110:12]
  assign n32_I0_15 = n31_O_15; // @[Top.scala 110:12]
  assign n32_I1_0 = n30_O_0; // @[Top.scala 111:12]
  assign n32_I1_1 = n30_O_1; // @[Top.scala 111:12]
  assign n32_I1_2 = n30_O_2; // @[Top.scala 111:12]
  assign n32_I1_3 = n30_O_3; // @[Top.scala 111:12]
  assign n32_I1_4 = n30_O_4; // @[Top.scala 111:12]
  assign n32_I1_5 = n30_O_5; // @[Top.scala 111:12]
  assign n32_I1_6 = n30_O_6; // @[Top.scala 111:12]
  assign n32_I1_7 = n30_O_7; // @[Top.scala 111:12]
  assign n32_I1_8 = n30_O_8; // @[Top.scala 111:12]
  assign n32_I1_9 = n30_O_9; // @[Top.scala 111:12]
  assign n32_I1_10 = n30_O_10; // @[Top.scala 111:12]
  assign n32_I1_11 = n30_O_11; // @[Top.scala 111:12]
  assign n32_I1_12 = n30_O_12; // @[Top.scala 111:12]
  assign n32_I1_13 = n30_O_13; // @[Top.scala 111:12]
  assign n32_I1_14 = n30_O_14; // @[Top.scala 111:12]
  assign n32_I1_15 = n30_O_15; // @[Top.scala 111:12]
  assign n39_valid_up = n32_valid_down & n2_valid_down; // @[Top.scala 116:18]
  assign n39_I0_0_0 = n32_O_0_0; // @[Top.scala 114:12]
  assign n39_I0_0_1 = n32_O_0_1; // @[Top.scala 114:12]
  assign n39_I0_1_0 = n32_O_1_0; // @[Top.scala 114:12]
  assign n39_I0_1_1 = n32_O_1_1; // @[Top.scala 114:12]
  assign n39_I0_2_0 = n32_O_2_0; // @[Top.scala 114:12]
  assign n39_I0_2_1 = n32_O_2_1; // @[Top.scala 114:12]
  assign n39_I0_3_0 = n32_O_3_0; // @[Top.scala 114:12]
  assign n39_I0_3_1 = n32_O_3_1; // @[Top.scala 114:12]
  assign n39_I0_4_0 = n32_O_4_0; // @[Top.scala 114:12]
  assign n39_I0_4_1 = n32_O_4_1; // @[Top.scala 114:12]
  assign n39_I0_5_0 = n32_O_5_0; // @[Top.scala 114:12]
  assign n39_I0_5_1 = n32_O_5_1; // @[Top.scala 114:12]
  assign n39_I0_6_0 = n32_O_6_0; // @[Top.scala 114:12]
  assign n39_I0_6_1 = n32_O_6_1; // @[Top.scala 114:12]
  assign n39_I0_7_0 = n32_O_7_0; // @[Top.scala 114:12]
  assign n39_I0_7_1 = n32_O_7_1; // @[Top.scala 114:12]
  assign n39_I0_8_0 = n32_O_8_0; // @[Top.scala 114:12]
  assign n39_I0_8_1 = n32_O_8_1; // @[Top.scala 114:12]
  assign n39_I0_9_0 = n32_O_9_0; // @[Top.scala 114:12]
  assign n39_I0_9_1 = n32_O_9_1; // @[Top.scala 114:12]
  assign n39_I0_10_0 = n32_O_10_0; // @[Top.scala 114:12]
  assign n39_I0_10_1 = n32_O_10_1; // @[Top.scala 114:12]
  assign n39_I0_11_0 = n32_O_11_0; // @[Top.scala 114:12]
  assign n39_I0_11_1 = n32_O_11_1; // @[Top.scala 114:12]
  assign n39_I0_12_0 = n32_O_12_0; // @[Top.scala 114:12]
  assign n39_I0_12_1 = n32_O_12_1; // @[Top.scala 114:12]
  assign n39_I0_13_0 = n32_O_13_0; // @[Top.scala 114:12]
  assign n39_I0_13_1 = n32_O_13_1; // @[Top.scala 114:12]
  assign n39_I0_14_0 = n32_O_14_0; // @[Top.scala 114:12]
  assign n39_I0_14_1 = n32_O_14_1; // @[Top.scala 114:12]
  assign n39_I0_15_0 = n32_O_15_0; // @[Top.scala 114:12]
  assign n39_I0_15_1 = n32_O_15_1; // @[Top.scala 114:12]
  assign n39_I1_0 = n2_O_0; // @[Top.scala 115:12]
  assign n39_I1_1 = n2_O_1; // @[Top.scala 115:12]
  assign n39_I1_2 = n2_O_2; // @[Top.scala 115:12]
  assign n39_I1_3 = n2_O_3; // @[Top.scala 115:12]
  assign n39_I1_4 = n2_O_4; // @[Top.scala 115:12]
  assign n39_I1_5 = n2_O_5; // @[Top.scala 115:12]
  assign n39_I1_6 = n2_O_6; // @[Top.scala 115:12]
  assign n39_I1_7 = n2_O_7; // @[Top.scala 115:12]
  assign n39_I1_8 = n2_O_8; // @[Top.scala 115:12]
  assign n39_I1_9 = n2_O_9; // @[Top.scala 115:12]
  assign n39_I1_10 = n2_O_10; // @[Top.scala 115:12]
  assign n39_I1_11 = n2_O_11; // @[Top.scala 115:12]
  assign n39_I1_12 = n2_O_12; // @[Top.scala 115:12]
  assign n39_I1_13 = n2_O_13; // @[Top.scala 115:12]
  assign n39_I1_14 = n2_O_14; // @[Top.scala 115:12]
  assign n39_I1_15 = n2_O_15; // @[Top.scala 115:12]
  assign n48_valid_up = n39_valid_down; // @[Top.scala 119:18]
  assign n48_I_0_0 = n39_O_0_0; // @[Top.scala 118:11]
  assign n48_I_0_1 = n39_O_0_1; // @[Top.scala 118:11]
  assign n48_I_0_2 = n39_O_0_2; // @[Top.scala 118:11]
  assign n48_I_1_0 = n39_O_1_0; // @[Top.scala 118:11]
  assign n48_I_1_1 = n39_O_1_1; // @[Top.scala 118:11]
  assign n48_I_1_2 = n39_O_1_2; // @[Top.scala 118:11]
  assign n48_I_2_0 = n39_O_2_0; // @[Top.scala 118:11]
  assign n48_I_2_1 = n39_O_2_1; // @[Top.scala 118:11]
  assign n48_I_2_2 = n39_O_2_2; // @[Top.scala 118:11]
  assign n48_I_3_0 = n39_O_3_0; // @[Top.scala 118:11]
  assign n48_I_3_1 = n39_O_3_1; // @[Top.scala 118:11]
  assign n48_I_3_2 = n39_O_3_2; // @[Top.scala 118:11]
  assign n48_I_4_0 = n39_O_4_0; // @[Top.scala 118:11]
  assign n48_I_4_1 = n39_O_4_1; // @[Top.scala 118:11]
  assign n48_I_4_2 = n39_O_4_2; // @[Top.scala 118:11]
  assign n48_I_5_0 = n39_O_5_0; // @[Top.scala 118:11]
  assign n48_I_5_1 = n39_O_5_1; // @[Top.scala 118:11]
  assign n48_I_5_2 = n39_O_5_2; // @[Top.scala 118:11]
  assign n48_I_6_0 = n39_O_6_0; // @[Top.scala 118:11]
  assign n48_I_6_1 = n39_O_6_1; // @[Top.scala 118:11]
  assign n48_I_6_2 = n39_O_6_2; // @[Top.scala 118:11]
  assign n48_I_7_0 = n39_O_7_0; // @[Top.scala 118:11]
  assign n48_I_7_1 = n39_O_7_1; // @[Top.scala 118:11]
  assign n48_I_7_2 = n39_O_7_2; // @[Top.scala 118:11]
  assign n48_I_8_0 = n39_O_8_0; // @[Top.scala 118:11]
  assign n48_I_8_1 = n39_O_8_1; // @[Top.scala 118:11]
  assign n48_I_8_2 = n39_O_8_2; // @[Top.scala 118:11]
  assign n48_I_9_0 = n39_O_9_0; // @[Top.scala 118:11]
  assign n48_I_9_1 = n39_O_9_1; // @[Top.scala 118:11]
  assign n48_I_9_2 = n39_O_9_2; // @[Top.scala 118:11]
  assign n48_I_10_0 = n39_O_10_0; // @[Top.scala 118:11]
  assign n48_I_10_1 = n39_O_10_1; // @[Top.scala 118:11]
  assign n48_I_10_2 = n39_O_10_2; // @[Top.scala 118:11]
  assign n48_I_11_0 = n39_O_11_0; // @[Top.scala 118:11]
  assign n48_I_11_1 = n39_O_11_1; // @[Top.scala 118:11]
  assign n48_I_11_2 = n39_O_11_2; // @[Top.scala 118:11]
  assign n48_I_12_0 = n39_O_12_0; // @[Top.scala 118:11]
  assign n48_I_12_1 = n39_O_12_1; // @[Top.scala 118:11]
  assign n48_I_12_2 = n39_O_12_2; // @[Top.scala 118:11]
  assign n48_I_13_0 = n39_O_13_0; // @[Top.scala 118:11]
  assign n48_I_13_1 = n39_O_13_1; // @[Top.scala 118:11]
  assign n48_I_13_2 = n39_O_13_2; // @[Top.scala 118:11]
  assign n48_I_14_0 = n39_O_14_0; // @[Top.scala 118:11]
  assign n48_I_14_1 = n39_O_14_1; // @[Top.scala 118:11]
  assign n48_I_14_2 = n39_O_14_2; // @[Top.scala 118:11]
  assign n48_I_15_0 = n39_O_15_0; // @[Top.scala 118:11]
  assign n48_I_15_1 = n39_O_15_1; // @[Top.scala 118:11]
  assign n48_I_15_2 = n39_O_15_2; // @[Top.scala 118:11]
  assign n55_valid_up = n48_valid_down; // @[Top.scala 122:18]
  assign n55_I_0_0_0 = n48_O_0_0_0; // @[Top.scala 121:11]
  assign n55_I_0_0_1 = n48_O_0_0_1; // @[Top.scala 121:11]
  assign n55_I_0_0_2 = n48_O_0_0_2; // @[Top.scala 121:11]
  assign n55_I_1_0_0 = n48_O_1_0_0; // @[Top.scala 121:11]
  assign n55_I_1_0_1 = n48_O_1_0_1; // @[Top.scala 121:11]
  assign n55_I_1_0_2 = n48_O_1_0_2; // @[Top.scala 121:11]
  assign n55_I_2_0_0 = n48_O_2_0_0; // @[Top.scala 121:11]
  assign n55_I_2_0_1 = n48_O_2_0_1; // @[Top.scala 121:11]
  assign n55_I_2_0_2 = n48_O_2_0_2; // @[Top.scala 121:11]
  assign n55_I_3_0_0 = n48_O_3_0_0; // @[Top.scala 121:11]
  assign n55_I_3_0_1 = n48_O_3_0_1; // @[Top.scala 121:11]
  assign n55_I_3_0_2 = n48_O_3_0_2; // @[Top.scala 121:11]
  assign n55_I_4_0_0 = n48_O_4_0_0; // @[Top.scala 121:11]
  assign n55_I_4_0_1 = n48_O_4_0_1; // @[Top.scala 121:11]
  assign n55_I_4_0_2 = n48_O_4_0_2; // @[Top.scala 121:11]
  assign n55_I_5_0_0 = n48_O_5_0_0; // @[Top.scala 121:11]
  assign n55_I_5_0_1 = n48_O_5_0_1; // @[Top.scala 121:11]
  assign n55_I_5_0_2 = n48_O_5_0_2; // @[Top.scala 121:11]
  assign n55_I_6_0_0 = n48_O_6_0_0; // @[Top.scala 121:11]
  assign n55_I_6_0_1 = n48_O_6_0_1; // @[Top.scala 121:11]
  assign n55_I_6_0_2 = n48_O_6_0_2; // @[Top.scala 121:11]
  assign n55_I_7_0_0 = n48_O_7_0_0; // @[Top.scala 121:11]
  assign n55_I_7_0_1 = n48_O_7_0_1; // @[Top.scala 121:11]
  assign n55_I_7_0_2 = n48_O_7_0_2; // @[Top.scala 121:11]
  assign n55_I_8_0_0 = n48_O_8_0_0; // @[Top.scala 121:11]
  assign n55_I_8_0_1 = n48_O_8_0_1; // @[Top.scala 121:11]
  assign n55_I_8_0_2 = n48_O_8_0_2; // @[Top.scala 121:11]
  assign n55_I_9_0_0 = n48_O_9_0_0; // @[Top.scala 121:11]
  assign n55_I_9_0_1 = n48_O_9_0_1; // @[Top.scala 121:11]
  assign n55_I_9_0_2 = n48_O_9_0_2; // @[Top.scala 121:11]
  assign n55_I_10_0_0 = n48_O_10_0_0; // @[Top.scala 121:11]
  assign n55_I_10_0_1 = n48_O_10_0_1; // @[Top.scala 121:11]
  assign n55_I_10_0_2 = n48_O_10_0_2; // @[Top.scala 121:11]
  assign n55_I_11_0_0 = n48_O_11_0_0; // @[Top.scala 121:11]
  assign n55_I_11_0_1 = n48_O_11_0_1; // @[Top.scala 121:11]
  assign n55_I_11_0_2 = n48_O_11_0_2; // @[Top.scala 121:11]
  assign n55_I_12_0_0 = n48_O_12_0_0; // @[Top.scala 121:11]
  assign n55_I_12_0_1 = n48_O_12_0_1; // @[Top.scala 121:11]
  assign n55_I_12_0_2 = n48_O_12_0_2; // @[Top.scala 121:11]
  assign n55_I_13_0_0 = n48_O_13_0_0; // @[Top.scala 121:11]
  assign n55_I_13_0_1 = n48_O_13_0_1; // @[Top.scala 121:11]
  assign n55_I_13_0_2 = n48_O_13_0_2; // @[Top.scala 121:11]
  assign n55_I_14_0_0 = n48_O_14_0_0; // @[Top.scala 121:11]
  assign n55_I_14_0_1 = n48_O_14_0_1; // @[Top.scala 121:11]
  assign n55_I_14_0_2 = n48_O_14_0_2; // @[Top.scala 121:11]
  assign n55_I_15_0_0 = n48_O_15_0_0; // @[Top.scala 121:11]
  assign n55_I_15_0_1 = n48_O_15_0_1; // @[Top.scala 121:11]
  assign n55_I_15_0_2 = n48_O_15_0_2; // @[Top.scala 121:11]
  assign n56_valid_up = n29_valid_down & n55_valid_down; // @[Top.scala 126:18]
  assign n56_I0_0_0 = n29_O_0_0; // @[Top.scala 124:12]
  assign n56_I0_0_1 = n29_O_0_1; // @[Top.scala 124:12]
  assign n56_I0_0_2 = n29_O_0_2; // @[Top.scala 124:12]
  assign n56_I0_1_0 = n29_O_1_0; // @[Top.scala 124:12]
  assign n56_I0_1_1 = n29_O_1_1; // @[Top.scala 124:12]
  assign n56_I0_1_2 = n29_O_1_2; // @[Top.scala 124:12]
  assign n56_I0_2_0 = n29_O_2_0; // @[Top.scala 124:12]
  assign n56_I0_2_1 = n29_O_2_1; // @[Top.scala 124:12]
  assign n56_I0_2_2 = n29_O_2_2; // @[Top.scala 124:12]
  assign n56_I0_3_0 = n29_O_3_0; // @[Top.scala 124:12]
  assign n56_I0_3_1 = n29_O_3_1; // @[Top.scala 124:12]
  assign n56_I0_3_2 = n29_O_3_2; // @[Top.scala 124:12]
  assign n56_I0_4_0 = n29_O_4_0; // @[Top.scala 124:12]
  assign n56_I0_4_1 = n29_O_4_1; // @[Top.scala 124:12]
  assign n56_I0_4_2 = n29_O_4_2; // @[Top.scala 124:12]
  assign n56_I0_5_0 = n29_O_5_0; // @[Top.scala 124:12]
  assign n56_I0_5_1 = n29_O_5_1; // @[Top.scala 124:12]
  assign n56_I0_5_2 = n29_O_5_2; // @[Top.scala 124:12]
  assign n56_I0_6_0 = n29_O_6_0; // @[Top.scala 124:12]
  assign n56_I0_6_1 = n29_O_6_1; // @[Top.scala 124:12]
  assign n56_I0_6_2 = n29_O_6_2; // @[Top.scala 124:12]
  assign n56_I0_7_0 = n29_O_7_0; // @[Top.scala 124:12]
  assign n56_I0_7_1 = n29_O_7_1; // @[Top.scala 124:12]
  assign n56_I0_7_2 = n29_O_7_2; // @[Top.scala 124:12]
  assign n56_I0_8_0 = n29_O_8_0; // @[Top.scala 124:12]
  assign n56_I0_8_1 = n29_O_8_1; // @[Top.scala 124:12]
  assign n56_I0_8_2 = n29_O_8_2; // @[Top.scala 124:12]
  assign n56_I0_9_0 = n29_O_9_0; // @[Top.scala 124:12]
  assign n56_I0_9_1 = n29_O_9_1; // @[Top.scala 124:12]
  assign n56_I0_9_2 = n29_O_9_2; // @[Top.scala 124:12]
  assign n56_I0_10_0 = n29_O_10_0; // @[Top.scala 124:12]
  assign n56_I0_10_1 = n29_O_10_1; // @[Top.scala 124:12]
  assign n56_I0_10_2 = n29_O_10_2; // @[Top.scala 124:12]
  assign n56_I0_11_0 = n29_O_11_0; // @[Top.scala 124:12]
  assign n56_I0_11_1 = n29_O_11_1; // @[Top.scala 124:12]
  assign n56_I0_11_2 = n29_O_11_2; // @[Top.scala 124:12]
  assign n56_I0_12_0 = n29_O_12_0; // @[Top.scala 124:12]
  assign n56_I0_12_1 = n29_O_12_1; // @[Top.scala 124:12]
  assign n56_I0_12_2 = n29_O_12_2; // @[Top.scala 124:12]
  assign n56_I0_13_0 = n29_O_13_0; // @[Top.scala 124:12]
  assign n56_I0_13_1 = n29_O_13_1; // @[Top.scala 124:12]
  assign n56_I0_13_2 = n29_O_13_2; // @[Top.scala 124:12]
  assign n56_I0_14_0 = n29_O_14_0; // @[Top.scala 124:12]
  assign n56_I0_14_1 = n29_O_14_1; // @[Top.scala 124:12]
  assign n56_I0_14_2 = n29_O_14_2; // @[Top.scala 124:12]
  assign n56_I0_15_0 = n29_O_15_0; // @[Top.scala 124:12]
  assign n56_I0_15_1 = n29_O_15_1; // @[Top.scala 124:12]
  assign n56_I0_15_2 = n29_O_15_2; // @[Top.scala 124:12]
  assign n56_I1_0_0 = n55_O_0_0; // @[Top.scala 125:12]
  assign n56_I1_0_1 = n55_O_0_1; // @[Top.scala 125:12]
  assign n56_I1_0_2 = n55_O_0_2; // @[Top.scala 125:12]
  assign n56_I1_1_0 = n55_O_1_0; // @[Top.scala 125:12]
  assign n56_I1_1_1 = n55_O_1_1; // @[Top.scala 125:12]
  assign n56_I1_1_2 = n55_O_1_2; // @[Top.scala 125:12]
  assign n56_I1_2_0 = n55_O_2_0; // @[Top.scala 125:12]
  assign n56_I1_2_1 = n55_O_2_1; // @[Top.scala 125:12]
  assign n56_I1_2_2 = n55_O_2_2; // @[Top.scala 125:12]
  assign n56_I1_3_0 = n55_O_3_0; // @[Top.scala 125:12]
  assign n56_I1_3_1 = n55_O_3_1; // @[Top.scala 125:12]
  assign n56_I1_3_2 = n55_O_3_2; // @[Top.scala 125:12]
  assign n56_I1_4_0 = n55_O_4_0; // @[Top.scala 125:12]
  assign n56_I1_4_1 = n55_O_4_1; // @[Top.scala 125:12]
  assign n56_I1_4_2 = n55_O_4_2; // @[Top.scala 125:12]
  assign n56_I1_5_0 = n55_O_5_0; // @[Top.scala 125:12]
  assign n56_I1_5_1 = n55_O_5_1; // @[Top.scala 125:12]
  assign n56_I1_5_2 = n55_O_5_2; // @[Top.scala 125:12]
  assign n56_I1_6_0 = n55_O_6_0; // @[Top.scala 125:12]
  assign n56_I1_6_1 = n55_O_6_1; // @[Top.scala 125:12]
  assign n56_I1_6_2 = n55_O_6_2; // @[Top.scala 125:12]
  assign n56_I1_7_0 = n55_O_7_0; // @[Top.scala 125:12]
  assign n56_I1_7_1 = n55_O_7_1; // @[Top.scala 125:12]
  assign n56_I1_7_2 = n55_O_7_2; // @[Top.scala 125:12]
  assign n56_I1_8_0 = n55_O_8_0; // @[Top.scala 125:12]
  assign n56_I1_8_1 = n55_O_8_1; // @[Top.scala 125:12]
  assign n56_I1_8_2 = n55_O_8_2; // @[Top.scala 125:12]
  assign n56_I1_9_0 = n55_O_9_0; // @[Top.scala 125:12]
  assign n56_I1_9_1 = n55_O_9_1; // @[Top.scala 125:12]
  assign n56_I1_9_2 = n55_O_9_2; // @[Top.scala 125:12]
  assign n56_I1_10_0 = n55_O_10_0; // @[Top.scala 125:12]
  assign n56_I1_10_1 = n55_O_10_1; // @[Top.scala 125:12]
  assign n56_I1_10_2 = n55_O_10_2; // @[Top.scala 125:12]
  assign n56_I1_11_0 = n55_O_11_0; // @[Top.scala 125:12]
  assign n56_I1_11_1 = n55_O_11_1; // @[Top.scala 125:12]
  assign n56_I1_11_2 = n55_O_11_2; // @[Top.scala 125:12]
  assign n56_I1_12_0 = n55_O_12_0; // @[Top.scala 125:12]
  assign n56_I1_12_1 = n55_O_12_1; // @[Top.scala 125:12]
  assign n56_I1_12_2 = n55_O_12_2; // @[Top.scala 125:12]
  assign n56_I1_13_0 = n55_O_13_0; // @[Top.scala 125:12]
  assign n56_I1_13_1 = n55_O_13_1; // @[Top.scala 125:12]
  assign n56_I1_13_2 = n55_O_13_2; // @[Top.scala 125:12]
  assign n56_I1_14_0 = n55_O_14_0; // @[Top.scala 125:12]
  assign n56_I1_14_1 = n55_O_14_1; // @[Top.scala 125:12]
  assign n56_I1_14_2 = n55_O_14_2; // @[Top.scala 125:12]
  assign n56_I1_15_0 = n55_O_15_0; // @[Top.scala 125:12]
  assign n56_I1_15_1 = n55_O_15_1; // @[Top.scala 125:12]
  assign n56_I1_15_2 = n55_O_15_2; // @[Top.scala 125:12]
  assign n63_clock = clock;
  assign n63_valid_up = n1_valid_down; // @[Top.scala 129:18]
  assign n63_I_0 = n1_O_0; // @[Top.scala 128:11]
  assign n63_I_1 = n1_O_1; // @[Top.scala 128:11]
  assign n63_I_2 = n1_O_2; // @[Top.scala 128:11]
  assign n63_I_3 = n1_O_3; // @[Top.scala 128:11]
  assign n63_I_4 = n1_O_4; // @[Top.scala 128:11]
  assign n63_I_5 = n1_O_5; // @[Top.scala 128:11]
  assign n63_I_6 = n1_O_6; // @[Top.scala 128:11]
  assign n63_I_7 = n1_O_7; // @[Top.scala 128:11]
  assign n63_I_8 = n1_O_8; // @[Top.scala 128:11]
  assign n63_I_9 = n1_O_9; // @[Top.scala 128:11]
  assign n63_I_10 = n1_O_10; // @[Top.scala 128:11]
  assign n63_I_11 = n1_O_11; // @[Top.scala 128:11]
  assign n63_I_12 = n1_O_12; // @[Top.scala 128:11]
  assign n63_I_13 = n1_O_13; // @[Top.scala 128:11]
  assign n63_I_14 = n1_O_14; // @[Top.scala 128:11]
  assign n63_I_15 = n1_O_15; // @[Top.scala 128:11]
  assign n64_clock = clock;
  assign n64_valid_up = n63_valid_down; // @[Top.scala 132:18]
  assign n64_I_0 = n63_O_0; // @[Top.scala 131:11]
  assign n64_I_1 = n63_O_1; // @[Top.scala 131:11]
  assign n64_I_2 = n63_O_2; // @[Top.scala 131:11]
  assign n64_I_3 = n63_O_3; // @[Top.scala 131:11]
  assign n64_I_4 = n63_O_4; // @[Top.scala 131:11]
  assign n64_I_5 = n63_O_5; // @[Top.scala 131:11]
  assign n64_I_6 = n63_O_6; // @[Top.scala 131:11]
  assign n64_I_7 = n63_O_7; // @[Top.scala 131:11]
  assign n64_I_8 = n63_O_8; // @[Top.scala 131:11]
  assign n64_I_9 = n63_O_9; // @[Top.scala 131:11]
  assign n64_I_10 = n63_O_10; // @[Top.scala 131:11]
  assign n64_I_11 = n63_O_11; // @[Top.scala 131:11]
  assign n64_I_12 = n63_O_12; // @[Top.scala 131:11]
  assign n64_I_13 = n63_O_13; // @[Top.scala 131:11]
  assign n64_I_14 = n63_O_14; // @[Top.scala 131:11]
  assign n64_I_15 = n63_O_15; // @[Top.scala 131:11]
  assign n65_valid_up = n64_valid_down & n63_valid_down; // @[Top.scala 136:18]
  assign n65_I0_0 = n64_O_0; // @[Top.scala 134:12]
  assign n65_I0_1 = n64_O_1; // @[Top.scala 134:12]
  assign n65_I0_2 = n64_O_2; // @[Top.scala 134:12]
  assign n65_I0_3 = n64_O_3; // @[Top.scala 134:12]
  assign n65_I0_4 = n64_O_4; // @[Top.scala 134:12]
  assign n65_I0_5 = n64_O_5; // @[Top.scala 134:12]
  assign n65_I0_6 = n64_O_6; // @[Top.scala 134:12]
  assign n65_I0_7 = n64_O_7; // @[Top.scala 134:12]
  assign n65_I0_8 = n64_O_8; // @[Top.scala 134:12]
  assign n65_I0_9 = n64_O_9; // @[Top.scala 134:12]
  assign n65_I0_10 = n64_O_10; // @[Top.scala 134:12]
  assign n65_I0_11 = n64_O_11; // @[Top.scala 134:12]
  assign n65_I0_12 = n64_O_12; // @[Top.scala 134:12]
  assign n65_I0_13 = n64_O_13; // @[Top.scala 134:12]
  assign n65_I0_14 = n64_O_14; // @[Top.scala 134:12]
  assign n65_I0_15 = n64_O_15; // @[Top.scala 134:12]
  assign n65_I1_0 = n63_O_0; // @[Top.scala 135:12]
  assign n65_I1_1 = n63_O_1; // @[Top.scala 135:12]
  assign n65_I1_2 = n63_O_2; // @[Top.scala 135:12]
  assign n65_I1_3 = n63_O_3; // @[Top.scala 135:12]
  assign n65_I1_4 = n63_O_4; // @[Top.scala 135:12]
  assign n65_I1_5 = n63_O_5; // @[Top.scala 135:12]
  assign n65_I1_6 = n63_O_6; // @[Top.scala 135:12]
  assign n65_I1_7 = n63_O_7; // @[Top.scala 135:12]
  assign n65_I1_8 = n63_O_8; // @[Top.scala 135:12]
  assign n65_I1_9 = n63_O_9; // @[Top.scala 135:12]
  assign n65_I1_10 = n63_O_10; // @[Top.scala 135:12]
  assign n65_I1_11 = n63_O_11; // @[Top.scala 135:12]
  assign n65_I1_12 = n63_O_12; // @[Top.scala 135:12]
  assign n65_I1_13 = n63_O_13; // @[Top.scala 135:12]
  assign n65_I1_14 = n63_O_14; // @[Top.scala 135:12]
  assign n65_I1_15 = n63_O_15; // @[Top.scala 135:12]
  assign n72_valid_up = n65_valid_down & n1_valid_down; // @[Top.scala 140:18]
  assign n72_I0_0_0 = n65_O_0_0; // @[Top.scala 138:12]
  assign n72_I0_0_1 = n65_O_0_1; // @[Top.scala 138:12]
  assign n72_I0_1_0 = n65_O_1_0; // @[Top.scala 138:12]
  assign n72_I0_1_1 = n65_O_1_1; // @[Top.scala 138:12]
  assign n72_I0_2_0 = n65_O_2_0; // @[Top.scala 138:12]
  assign n72_I0_2_1 = n65_O_2_1; // @[Top.scala 138:12]
  assign n72_I0_3_0 = n65_O_3_0; // @[Top.scala 138:12]
  assign n72_I0_3_1 = n65_O_3_1; // @[Top.scala 138:12]
  assign n72_I0_4_0 = n65_O_4_0; // @[Top.scala 138:12]
  assign n72_I0_4_1 = n65_O_4_1; // @[Top.scala 138:12]
  assign n72_I0_5_0 = n65_O_5_0; // @[Top.scala 138:12]
  assign n72_I0_5_1 = n65_O_5_1; // @[Top.scala 138:12]
  assign n72_I0_6_0 = n65_O_6_0; // @[Top.scala 138:12]
  assign n72_I0_6_1 = n65_O_6_1; // @[Top.scala 138:12]
  assign n72_I0_7_0 = n65_O_7_0; // @[Top.scala 138:12]
  assign n72_I0_7_1 = n65_O_7_1; // @[Top.scala 138:12]
  assign n72_I0_8_0 = n65_O_8_0; // @[Top.scala 138:12]
  assign n72_I0_8_1 = n65_O_8_1; // @[Top.scala 138:12]
  assign n72_I0_9_0 = n65_O_9_0; // @[Top.scala 138:12]
  assign n72_I0_9_1 = n65_O_9_1; // @[Top.scala 138:12]
  assign n72_I0_10_0 = n65_O_10_0; // @[Top.scala 138:12]
  assign n72_I0_10_1 = n65_O_10_1; // @[Top.scala 138:12]
  assign n72_I0_11_0 = n65_O_11_0; // @[Top.scala 138:12]
  assign n72_I0_11_1 = n65_O_11_1; // @[Top.scala 138:12]
  assign n72_I0_12_0 = n65_O_12_0; // @[Top.scala 138:12]
  assign n72_I0_12_1 = n65_O_12_1; // @[Top.scala 138:12]
  assign n72_I0_13_0 = n65_O_13_0; // @[Top.scala 138:12]
  assign n72_I0_13_1 = n65_O_13_1; // @[Top.scala 138:12]
  assign n72_I0_14_0 = n65_O_14_0; // @[Top.scala 138:12]
  assign n72_I0_14_1 = n65_O_14_1; // @[Top.scala 138:12]
  assign n72_I0_15_0 = n65_O_15_0; // @[Top.scala 138:12]
  assign n72_I0_15_1 = n65_O_15_1; // @[Top.scala 138:12]
  assign n72_I1_0 = n1_O_0; // @[Top.scala 139:12]
  assign n72_I1_1 = n1_O_1; // @[Top.scala 139:12]
  assign n72_I1_2 = n1_O_2; // @[Top.scala 139:12]
  assign n72_I1_3 = n1_O_3; // @[Top.scala 139:12]
  assign n72_I1_4 = n1_O_4; // @[Top.scala 139:12]
  assign n72_I1_5 = n1_O_5; // @[Top.scala 139:12]
  assign n72_I1_6 = n1_O_6; // @[Top.scala 139:12]
  assign n72_I1_7 = n1_O_7; // @[Top.scala 139:12]
  assign n72_I1_8 = n1_O_8; // @[Top.scala 139:12]
  assign n72_I1_9 = n1_O_9; // @[Top.scala 139:12]
  assign n72_I1_10 = n1_O_10; // @[Top.scala 139:12]
  assign n72_I1_11 = n1_O_11; // @[Top.scala 139:12]
  assign n72_I1_12 = n1_O_12; // @[Top.scala 139:12]
  assign n72_I1_13 = n1_O_13; // @[Top.scala 139:12]
  assign n72_I1_14 = n1_O_14; // @[Top.scala 139:12]
  assign n72_I1_15 = n1_O_15; // @[Top.scala 139:12]
  assign n81_valid_up = n72_valid_down; // @[Top.scala 143:18]
  assign n81_I_0_0 = n72_O_0_0; // @[Top.scala 142:11]
  assign n81_I_0_1 = n72_O_0_1; // @[Top.scala 142:11]
  assign n81_I_0_2 = n72_O_0_2; // @[Top.scala 142:11]
  assign n81_I_1_0 = n72_O_1_0; // @[Top.scala 142:11]
  assign n81_I_1_1 = n72_O_1_1; // @[Top.scala 142:11]
  assign n81_I_1_2 = n72_O_1_2; // @[Top.scala 142:11]
  assign n81_I_2_0 = n72_O_2_0; // @[Top.scala 142:11]
  assign n81_I_2_1 = n72_O_2_1; // @[Top.scala 142:11]
  assign n81_I_2_2 = n72_O_2_2; // @[Top.scala 142:11]
  assign n81_I_3_0 = n72_O_3_0; // @[Top.scala 142:11]
  assign n81_I_3_1 = n72_O_3_1; // @[Top.scala 142:11]
  assign n81_I_3_2 = n72_O_3_2; // @[Top.scala 142:11]
  assign n81_I_4_0 = n72_O_4_0; // @[Top.scala 142:11]
  assign n81_I_4_1 = n72_O_4_1; // @[Top.scala 142:11]
  assign n81_I_4_2 = n72_O_4_2; // @[Top.scala 142:11]
  assign n81_I_5_0 = n72_O_5_0; // @[Top.scala 142:11]
  assign n81_I_5_1 = n72_O_5_1; // @[Top.scala 142:11]
  assign n81_I_5_2 = n72_O_5_2; // @[Top.scala 142:11]
  assign n81_I_6_0 = n72_O_6_0; // @[Top.scala 142:11]
  assign n81_I_6_1 = n72_O_6_1; // @[Top.scala 142:11]
  assign n81_I_6_2 = n72_O_6_2; // @[Top.scala 142:11]
  assign n81_I_7_0 = n72_O_7_0; // @[Top.scala 142:11]
  assign n81_I_7_1 = n72_O_7_1; // @[Top.scala 142:11]
  assign n81_I_7_2 = n72_O_7_2; // @[Top.scala 142:11]
  assign n81_I_8_0 = n72_O_8_0; // @[Top.scala 142:11]
  assign n81_I_8_1 = n72_O_8_1; // @[Top.scala 142:11]
  assign n81_I_8_2 = n72_O_8_2; // @[Top.scala 142:11]
  assign n81_I_9_0 = n72_O_9_0; // @[Top.scala 142:11]
  assign n81_I_9_1 = n72_O_9_1; // @[Top.scala 142:11]
  assign n81_I_9_2 = n72_O_9_2; // @[Top.scala 142:11]
  assign n81_I_10_0 = n72_O_10_0; // @[Top.scala 142:11]
  assign n81_I_10_1 = n72_O_10_1; // @[Top.scala 142:11]
  assign n81_I_10_2 = n72_O_10_2; // @[Top.scala 142:11]
  assign n81_I_11_0 = n72_O_11_0; // @[Top.scala 142:11]
  assign n81_I_11_1 = n72_O_11_1; // @[Top.scala 142:11]
  assign n81_I_11_2 = n72_O_11_2; // @[Top.scala 142:11]
  assign n81_I_12_0 = n72_O_12_0; // @[Top.scala 142:11]
  assign n81_I_12_1 = n72_O_12_1; // @[Top.scala 142:11]
  assign n81_I_12_2 = n72_O_12_2; // @[Top.scala 142:11]
  assign n81_I_13_0 = n72_O_13_0; // @[Top.scala 142:11]
  assign n81_I_13_1 = n72_O_13_1; // @[Top.scala 142:11]
  assign n81_I_13_2 = n72_O_13_2; // @[Top.scala 142:11]
  assign n81_I_14_0 = n72_O_14_0; // @[Top.scala 142:11]
  assign n81_I_14_1 = n72_O_14_1; // @[Top.scala 142:11]
  assign n81_I_14_2 = n72_O_14_2; // @[Top.scala 142:11]
  assign n81_I_15_0 = n72_O_15_0; // @[Top.scala 142:11]
  assign n81_I_15_1 = n72_O_15_1; // @[Top.scala 142:11]
  assign n81_I_15_2 = n72_O_15_2; // @[Top.scala 142:11]
  assign n88_valid_up = n81_valid_down; // @[Top.scala 146:18]
  assign n88_I_0_0_0 = n81_O_0_0_0; // @[Top.scala 145:11]
  assign n88_I_0_0_1 = n81_O_0_0_1; // @[Top.scala 145:11]
  assign n88_I_0_0_2 = n81_O_0_0_2; // @[Top.scala 145:11]
  assign n88_I_1_0_0 = n81_O_1_0_0; // @[Top.scala 145:11]
  assign n88_I_1_0_1 = n81_O_1_0_1; // @[Top.scala 145:11]
  assign n88_I_1_0_2 = n81_O_1_0_2; // @[Top.scala 145:11]
  assign n88_I_2_0_0 = n81_O_2_0_0; // @[Top.scala 145:11]
  assign n88_I_2_0_1 = n81_O_2_0_1; // @[Top.scala 145:11]
  assign n88_I_2_0_2 = n81_O_2_0_2; // @[Top.scala 145:11]
  assign n88_I_3_0_0 = n81_O_3_0_0; // @[Top.scala 145:11]
  assign n88_I_3_0_1 = n81_O_3_0_1; // @[Top.scala 145:11]
  assign n88_I_3_0_2 = n81_O_3_0_2; // @[Top.scala 145:11]
  assign n88_I_4_0_0 = n81_O_4_0_0; // @[Top.scala 145:11]
  assign n88_I_4_0_1 = n81_O_4_0_1; // @[Top.scala 145:11]
  assign n88_I_4_0_2 = n81_O_4_0_2; // @[Top.scala 145:11]
  assign n88_I_5_0_0 = n81_O_5_0_0; // @[Top.scala 145:11]
  assign n88_I_5_0_1 = n81_O_5_0_1; // @[Top.scala 145:11]
  assign n88_I_5_0_2 = n81_O_5_0_2; // @[Top.scala 145:11]
  assign n88_I_6_0_0 = n81_O_6_0_0; // @[Top.scala 145:11]
  assign n88_I_6_0_1 = n81_O_6_0_1; // @[Top.scala 145:11]
  assign n88_I_6_0_2 = n81_O_6_0_2; // @[Top.scala 145:11]
  assign n88_I_7_0_0 = n81_O_7_0_0; // @[Top.scala 145:11]
  assign n88_I_7_0_1 = n81_O_7_0_1; // @[Top.scala 145:11]
  assign n88_I_7_0_2 = n81_O_7_0_2; // @[Top.scala 145:11]
  assign n88_I_8_0_0 = n81_O_8_0_0; // @[Top.scala 145:11]
  assign n88_I_8_0_1 = n81_O_8_0_1; // @[Top.scala 145:11]
  assign n88_I_8_0_2 = n81_O_8_0_2; // @[Top.scala 145:11]
  assign n88_I_9_0_0 = n81_O_9_0_0; // @[Top.scala 145:11]
  assign n88_I_9_0_1 = n81_O_9_0_1; // @[Top.scala 145:11]
  assign n88_I_9_0_2 = n81_O_9_0_2; // @[Top.scala 145:11]
  assign n88_I_10_0_0 = n81_O_10_0_0; // @[Top.scala 145:11]
  assign n88_I_10_0_1 = n81_O_10_0_1; // @[Top.scala 145:11]
  assign n88_I_10_0_2 = n81_O_10_0_2; // @[Top.scala 145:11]
  assign n88_I_11_0_0 = n81_O_11_0_0; // @[Top.scala 145:11]
  assign n88_I_11_0_1 = n81_O_11_0_1; // @[Top.scala 145:11]
  assign n88_I_11_0_2 = n81_O_11_0_2; // @[Top.scala 145:11]
  assign n88_I_12_0_0 = n81_O_12_0_0; // @[Top.scala 145:11]
  assign n88_I_12_0_1 = n81_O_12_0_1; // @[Top.scala 145:11]
  assign n88_I_12_0_2 = n81_O_12_0_2; // @[Top.scala 145:11]
  assign n88_I_13_0_0 = n81_O_13_0_0; // @[Top.scala 145:11]
  assign n88_I_13_0_1 = n81_O_13_0_1; // @[Top.scala 145:11]
  assign n88_I_13_0_2 = n81_O_13_0_2; // @[Top.scala 145:11]
  assign n88_I_14_0_0 = n81_O_14_0_0; // @[Top.scala 145:11]
  assign n88_I_14_0_1 = n81_O_14_0_1; // @[Top.scala 145:11]
  assign n88_I_14_0_2 = n81_O_14_0_2; // @[Top.scala 145:11]
  assign n88_I_15_0_0 = n81_O_15_0_0; // @[Top.scala 145:11]
  assign n88_I_15_0_1 = n81_O_15_0_1; // @[Top.scala 145:11]
  assign n88_I_15_0_2 = n81_O_15_0_2; // @[Top.scala 145:11]
  assign n89_valid_up = n56_valid_down & n88_valid_down; // @[Top.scala 150:18]
  assign n89_I0_0_0_0 = n56_O_0_0_0; // @[Top.scala 148:12]
  assign n89_I0_0_0_1 = n56_O_0_0_1; // @[Top.scala 148:12]
  assign n89_I0_0_0_2 = n56_O_0_0_2; // @[Top.scala 148:12]
  assign n89_I0_0_1_0 = n56_O_0_1_0; // @[Top.scala 148:12]
  assign n89_I0_0_1_1 = n56_O_0_1_1; // @[Top.scala 148:12]
  assign n89_I0_0_1_2 = n56_O_0_1_2; // @[Top.scala 148:12]
  assign n89_I0_1_0_0 = n56_O_1_0_0; // @[Top.scala 148:12]
  assign n89_I0_1_0_1 = n56_O_1_0_1; // @[Top.scala 148:12]
  assign n89_I0_1_0_2 = n56_O_1_0_2; // @[Top.scala 148:12]
  assign n89_I0_1_1_0 = n56_O_1_1_0; // @[Top.scala 148:12]
  assign n89_I0_1_1_1 = n56_O_1_1_1; // @[Top.scala 148:12]
  assign n89_I0_1_1_2 = n56_O_1_1_2; // @[Top.scala 148:12]
  assign n89_I0_2_0_0 = n56_O_2_0_0; // @[Top.scala 148:12]
  assign n89_I0_2_0_1 = n56_O_2_0_1; // @[Top.scala 148:12]
  assign n89_I0_2_0_2 = n56_O_2_0_2; // @[Top.scala 148:12]
  assign n89_I0_2_1_0 = n56_O_2_1_0; // @[Top.scala 148:12]
  assign n89_I0_2_1_1 = n56_O_2_1_1; // @[Top.scala 148:12]
  assign n89_I0_2_1_2 = n56_O_2_1_2; // @[Top.scala 148:12]
  assign n89_I0_3_0_0 = n56_O_3_0_0; // @[Top.scala 148:12]
  assign n89_I0_3_0_1 = n56_O_3_0_1; // @[Top.scala 148:12]
  assign n89_I0_3_0_2 = n56_O_3_0_2; // @[Top.scala 148:12]
  assign n89_I0_3_1_0 = n56_O_3_1_0; // @[Top.scala 148:12]
  assign n89_I0_3_1_1 = n56_O_3_1_1; // @[Top.scala 148:12]
  assign n89_I0_3_1_2 = n56_O_3_1_2; // @[Top.scala 148:12]
  assign n89_I0_4_0_0 = n56_O_4_0_0; // @[Top.scala 148:12]
  assign n89_I0_4_0_1 = n56_O_4_0_1; // @[Top.scala 148:12]
  assign n89_I0_4_0_2 = n56_O_4_0_2; // @[Top.scala 148:12]
  assign n89_I0_4_1_0 = n56_O_4_1_0; // @[Top.scala 148:12]
  assign n89_I0_4_1_1 = n56_O_4_1_1; // @[Top.scala 148:12]
  assign n89_I0_4_1_2 = n56_O_4_1_2; // @[Top.scala 148:12]
  assign n89_I0_5_0_0 = n56_O_5_0_0; // @[Top.scala 148:12]
  assign n89_I0_5_0_1 = n56_O_5_0_1; // @[Top.scala 148:12]
  assign n89_I0_5_0_2 = n56_O_5_0_2; // @[Top.scala 148:12]
  assign n89_I0_5_1_0 = n56_O_5_1_0; // @[Top.scala 148:12]
  assign n89_I0_5_1_1 = n56_O_5_1_1; // @[Top.scala 148:12]
  assign n89_I0_5_1_2 = n56_O_5_1_2; // @[Top.scala 148:12]
  assign n89_I0_6_0_0 = n56_O_6_0_0; // @[Top.scala 148:12]
  assign n89_I0_6_0_1 = n56_O_6_0_1; // @[Top.scala 148:12]
  assign n89_I0_6_0_2 = n56_O_6_0_2; // @[Top.scala 148:12]
  assign n89_I0_6_1_0 = n56_O_6_1_0; // @[Top.scala 148:12]
  assign n89_I0_6_1_1 = n56_O_6_1_1; // @[Top.scala 148:12]
  assign n89_I0_6_1_2 = n56_O_6_1_2; // @[Top.scala 148:12]
  assign n89_I0_7_0_0 = n56_O_7_0_0; // @[Top.scala 148:12]
  assign n89_I0_7_0_1 = n56_O_7_0_1; // @[Top.scala 148:12]
  assign n89_I0_7_0_2 = n56_O_7_0_2; // @[Top.scala 148:12]
  assign n89_I0_7_1_0 = n56_O_7_1_0; // @[Top.scala 148:12]
  assign n89_I0_7_1_1 = n56_O_7_1_1; // @[Top.scala 148:12]
  assign n89_I0_7_1_2 = n56_O_7_1_2; // @[Top.scala 148:12]
  assign n89_I0_8_0_0 = n56_O_8_0_0; // @[Top.scala 148:12]
  assign n89_I0_8_0_1 = n56_O_8_0_1; // @[Top.scala 148:12]
  assign n89_I0_8_0_2 = n56_O_8_0_2; // @[Top.scala 148:12]
  assign n89_I0_8_1_0 = n56_O_8_1_0; // @[Top.scala 148:12]
  assign n89_I0_8_1_1 = n56_O_8_1_1; // @[Top.scala 148:12]
  assign n89_I0_8_1_2 = n56_O_8_1_2; // @[Top.scala 148:12]
  assign n89_I0_9_0_0 = n56_O_9_0_0; // @[Top.scala 148:12]
  assign n89_I0_9_0_1 = n56_O_9_0_1; // @[Top.scala 148:12]
  assign n89_I0_9_0_2 = n56_O_9_0_2; // @[Top.scala 148:12]
  assign n89_I0_9_1_0 = n56_O_9_1_0; // @[Top.scala 148:12]
  assign n89_I0_9_1_1 = n56_O_9_1_1; // @[Top.scala 148:12]
  assign n89_I0_9_1_2 = n56_O_9_1_2; // @[Top.scala 148:12]
  assign n89_I0_10_0_0 = n56_O_10_0_0; // @[Top.scala 148:12]
  assign n89_I0_10_0_1 = n56_O_10_0_1; // @[Top.scala 148:12]
  assign n89_I0_10_0_2 = n56_O_10_0_2; // @[Top.scala 148:12]
  assign n89_I0_10_1_0 = n56_O_10_1_0; // @[Top.scala 148:12]
  assign n89_I0_10_1_1 = n56_O_10_1_1; // @[Top.scala 148:12]
  assign n89_I0_10_1_2 = n56_O_10_1_2; // @[Top.scala 148:12]
  assign n89_I0_11_0_0 = n56_O_11_0_0; // @[Top.scala 148:12]
  assign n89_I0_11_0_1 = n56_O_11_0_1; // @[Top.scala 148:12]
  assign n89_I0_11_0_2 = n56_O_11_0_2; // @[Top.scala 148:12]
  assign n89_I0_11_1_0 = n56_O_11_1_0; // @[Top.scala 148:12]
  assign n89_I0_11_1_1 = n56_O_11_1_1; // @[Top.scala 148:12]
  assign n89_I0_11_1_2 = n56_O_11_1_2; // @[Top.scala 148:12]
  assign n89_I0_12_0_0 = n56_O_12_0_0; // @[Top.scala 148:12]
  assign n89_I0_12_0_1 = n56_O_12_0_1; // @[Top.scala 148:12]
  assign n89_I0_12_0_2 = n56_O_12_0_2; // @[Top.scala 148:12]
  assign n89_I0_12_1_0 = n56_O_12_1_0; // @[Top.scala 148:12]
  assign n89_I0_12_1_1 = n56_O_12_1_1; // @[Top.scala 148:12]
  assign n89_I0_12_1_2 = n56_O_12_1_2; // @[Top.scala 148:12]
  assign n89_I0_13_0_0 = n56_O_13_0_0; // @[Top.scala 148:12]
  assign n89_I0_13_0_1 = n56_O_13_0_1; // @[Top.scala 148:12]
  assign n89_I0_13_0_2 = n56_O_13_0_2; // @[Top.scala 148:12]
  assign n89_I0_13_1_0 = n56_O_13_1_0; // @[Top.scala 148:12]
  assign n89_I0_13_1_1 = n56_O_13_1_1; // @[Top.scala 148:12]
  assign n89_I0_13_1_2 = n56_O_13_1_2; // @[Top.scala 148:12]
  assign n89_I0_14_0_0 = n56_O_14_0_0; // @[Top.scala 148:12]
  assign n89_I0_14_0_1 = n56_O_14_0_1; // @[Top.scala 148:12]
  assign n89_I0_14_0_2 = n56_O_14_0_2; // @[Top.scala 148:12]
  assign n89_I0_14_1_0 = n56_O_14_1_0; // @[Top.scala 148:12]
  assign n89_I0_14_1_1 = n56_O_14_1_1; // @[Top.scala 148:12]
  assign n89_I0_14_1_2 = n56_O_14_1_2; // @[Top.scala 148:12]
  assign n89_I0_15_0_0 = n56_O_15_0_0; // @[Top.scala 148:12]
  assign n89_I0_15_0_1 = n56_O_15_0_1; // @[Top.scala 148:12]
  assign n89_I0_15_0_2 = n56_O_15_0_2; // @[Top.scala 148:12]
  assign n89_I0_15_1_0 = n56_O_15_1_0; // @[Top.scala 148:12]
  assign n89_I0_15_1_1 = n56_O_15_1_1; // @[Top.scala 148:12]
  assign n89_I0_15_1_2 = n56_O_15_1_2; // @[Top.scala 148:12]
  assign n89_I1_0_0 = n88_O_0_0; // @[Top.scala 149:12]
  assign n89_I1_0_1 = n88_O_0_1; // @[Top.scala 149:12]
  assign n89_I1_0_2 = n88_O_0_2; // @[Top.scala 149:12]
  assign n89_I1_1_0 = n88_O_1_0; // @[Top.scala 149:12]
  assign n89_I1_1_1 = n88_O_1_1; // @[Top.scala 149:12]
  assign n89_I1_1_2 = n88_O_1_2; // @[Top.scala 149:12]
  assign n89_I1_2_0 = n88_O_2_0; // @[Top.scala 149:12]
  assign n89_I1_2_1 = n88_O_2_1; // @[Top.scala 149:12]
  assign n89_I1_2_2 = n88_O_2_2; // @[Top.scala 149:12]
  assign n89_I1_3_0 = n88_O_3_0; // @[Top.scala 149:12]
  assign n89_I1_3_1 = n88_O_3_1; // @[Top.scala 149:12]
  assign n89_I1_3_2 = n88_O_3_2; // @[Top.scala 149:12]
  assign n89_I1_4_0 = n88_O_4_0; // @[Top.scala 149:12]
  assign n89_I1_4_1 = n88_O_4_1; // @[Top.scala 149:12]
  assign n89_I1_4_2 = n88_O_4_2; // @[Top.scala 149:12]
  assign n89_I1_5_0 = n88_O_5_0; // @[Top.scala 149:12]
  assign n89_I1_5_1 = n88_O_5_1; // @[Top.scala 149:12]
  assign n89_I1_5_2 = n88_O_5_2; // @[Top.scala 149:12]
  assign n89_I1_6_0 = n88_O_6_0; // @[Top.scala 149:12]
  assign n89_I1_6_1 = n88_O_6_1; // @[Top.scala 149:12]
  assign n89_I1_6_2 = n88_O_6_2; // @[Top.scala 149:12]
  assign n89_I1_7_0 = n88_O_7_0; // @[Top.scala 149:12]
  assign n89_I1_7_1 = n88_O_7_1; // @[Top.scala 149:12]
  assign n89_I1_7_2 = n88_O_7_2; // @[Top.scala 149:12]
  assign n89_I1_8_0 = n88_O_8_0; // @[Top.scala 149:12]
  assign n89_I1_8_1 = n88_O_8_1; // @[Top.scala 149:12]
  assign n89_I1_8_2 = n88_O_8_2; // @[Top.scala 149:12]
  assign n89_I1_9_0 = n88_O_9_0; // @[Top.scala 149:12]
  assign n89_I1_9_1 = n88_O_9_1; // @[Top.scala 149:12]
  assign n89_I1_9_2 = n88_O_9_2; // @[Top.scala 149:12]
  assign n89_I1_10_0 = n88_O_10_0; // @[Top.scala 149:12]
  assign n89_I1_10_1 = n88_O_10_1; // @[Top.scala 149:12]
  assign n89_I1_10_2 = n88_O_10_2; // @[Top.scala 149:12]
  assign n89_I1_11_0 = n88_O_11_0; // @[Top.scala 149:12]
  assign n89_I1_11_1 = n88_O_11_1; // @[Top.scala 149:12]
  assign n89_I1_11_2 = n88_O_11_2; // @[Top.scala 149:12]
  assign n89_I1_12_0 = n88_O_12_0; // @[Top.scala 149:12]
  assign n89_I1_12_1 = n88_O_12_1; // @[Top.scala 149:12]
  assign n89_I1_12_2 = n88_O_12_2; // @[Top.scala 149:12]
  assign n89_I1_13_0 = n88_O_13_0; // @[Top.scala 149:12]
  assign n89_I1_13_1 = n88_O_13_1; // @[Top.scala 149:12]
  assign n89_I1_13_2 = n88_O_13_2; // @[Top.scala 149:12]
  assign n89_I1_14_0 = n88_O_14_0; // @[Top.scala 149:12]
  assign n89_I1_14_1 = n88_O_14_1; // @[Top.scala 149:12]
  assign n89_I1_14_2 = n88_O_14_2; // @[Top.scala 149:12]
  assign n89_I1_15_0 = n88_O_15_0; // @[Top.scala 149:12]
  assign n89_I1_15_1 = n88_O_15_1; // @[Top.scala 149:12]
  assign n89_I1_15_2 = n88_O_15_2; // @[Top.scala 149:12]
  assign n98_valid_up = n89_valid_down; // @[Top.scala 153:18]
  assign n98_I_0_0_0 = n89_O_0_0_0; // @[Top.scala 152:11]
  assign n98_I_0_0_1 = n89_O_0_0_1; // @[Top.scala 152:11]
  assign n98_I_0_0_2 = n89_O_0_0_2; // @[Top.scala 152:11]
  assign n98_I_0_1_0 = n89_O_0_1_0; // @[Top.scala 152:11]
  assign n98_I_0_1_1 = n89_O_0_1_1; // @[Top.scala 152:11]
  assign n98_I_0_1_2 = n89_O_0_1_2; // @[Top.scala 152:11]
  assign n98_I_0_2_0 = n89_O_0_2_0; // @[Top.scala 152:11]
  assign n98_I_0_2_1 = n89_O_0_2_1; // @[Top.scala 152:11]
  assign n98_I_0_2_2 = n89_O_0_2_2; // @[Top.scala 152:11]
  assign n98_I_1_0_0 = n89_O_1_0_0; // @[Top.scala 152:11]
  assign n98_I_1_0_1 = n89_O_1_0_1; // @[Top.scala 152:11]
  assign n98_I_1_0_2 = n89_O_1_0_2; // @[Top.scala 152:11]
  assign n98_I_1_1_0 = n89_O_1_1_0; // @[Top.scala 152:11]
  assign n98_I_1_1_1 = n89_O_1_1_1; // @[Top.scala 152:11]
  assign n98_I_1_1_2 = n89_O_1_1_2; // @[Top.scala 152:11]
  assign n98_I_1_2_0 = n89_O_1_2_0; // @[Top.scala 152:11]
  assign n98_I_1_2_1 = n89_O_1_2_1; // @[Top.scala 152:11]
  assign n98_I_1_2_2 = n89_O_1_2_2; // @[Top.scala 152:11]
  assign n98_I_2_0_0 = n89_O_2_0_0; // @[Top.scala 152:11]
  assign n98_I_2_0_1 = n89_O_2_0_1; // @[Top.scala 152:11]
  assign n98_I_2_0_2 = n89_O_2_0_2; // @[Top.scala 152:11]
  assign n98_I_2_1_0 = n89_O_2_1_0; // @[Top.scala 152:11]
  assign n98_I_2_1_1 = n89_O_2_1_1; // @[Top.scala 152:11]
  assign n98_I_2_1_2 = n89_O_2_1_2; // @[Top.scala 152:11]
  assign n98_I_2_2_0 = n89_O_2_2_0; // @[Top.scala 152:11]
  assign n98_I_2_2_1 = n89_O_2_2_1; // @[Top.scala 152:11]
  assign n98_I_2_2_2 = n89_O_2_2_2; // @[Top.scala 152:11]
  assign n98_I_3_0_0 = n89_O_3_0_0; // @[Top.scala 152:11]
  assign n98_I_3_0_1 = n89_O_3_0_1; // @[Top.scala 152:11]
  assign n98_I_3_0_2 = n89_O_3_0_2; // @[Top.scala 152:11]
  assign n98_I_3_1_0 = n89_O_3_1_0; // @[Top.scala 152:11]
  assign n98_I_3_1_1 = n89_O_3_1_1; // @[Top.scala 152:11]
  assign n98_I_3_1_2 = n89_O_3_1_2; // @[Top.scala 152:11]
  assign n98_I_3_2_0 = n89_O_3_2_0; // @[Top.scala 152:11]
  assign n98_I_3_2_1 = n89_O_3_2_1; // @[Top.scala 152:11]
  assign n98_I_3_2_2 = n89_O_3_2_2; // @[Top.scala 152:11]
  assign n98_I_4_0_0 = n89_O_4_0_0; // @[Top.scala 152:11]
  assign n98_I_4_0_1 = n89_O_4_0_1; // @[Top.scala 152:11]
  assign n98_I_4_0_2 = n89_O_4_0_2; // @[Top.scala 152:11]
  assign n98_I_4_1_0 = n89_O_4_1_0; // @[Top.scala 152:11]
  assign n98_I_4_1_1 = n89_O_4_1_1; // @[Top.scala 152:11]
  assign n98_I_4_1_2 = n89_O_4_1_2; // @[Top.scala 152:11]
  assign n98_I_4_2_0 = n89_O_4_2_0; // @[Top.scala 152:11]
  assign n98_I_4_2_1 = n89_O_4_2_1; // @[Top.scala 152:11]
  assign n98_I_4_2_2 = n89_O_4_2_2; // @[Top.scala 152:11]
  assign n98_I_5_0_0 = n89_O_5_0_0; // @[Top.scala 152:11]
  assign n98_I_5_0_1 = n89_O_5_0_1; // @[Top.scala 152:11]
  assign n98_I_5_0_2 = n89_O_5_0_2; // @[Top.scala 152:11]
  assign n98_I_5_1_0 = n89_O_5_1_0; // @[Top.scala 152:11]
  assign n98_I_5_1_1 = n89_O_5_1_1; // @[Top.scala 152:11]
  assign n98_I_5_1_2 = n89_O_5_1_2; // @[Top.scala 152:11]
  assign n98_I_5_2_0 = n89_O_5_2_0; // @[Top.scala 152:11]
  assign n98_I_5_2_1 = n89_O_5_2_1; // @[Top.scala 152:11]
  assign n98_I_5_2_2 = n89_O_5_2_2; // @[Top.scala 152:11]
  assign n98_I_6_0_0 = n89_O_6_0_0; // @[Top.scala 152:11]
  assign n98_I_6_0_1 = n89_O_6_0_1; // @[Top.scala 152:11]
  assign n98_I_6_0_2 = n89_O_6_0_2; // @[Top.scala 152:11]
  assign n98_I_6_1_0 = n89_O_6_1_0; // @[Top.scala 152:11]
  assign n98_I_6_1_1 = n89_O_6_1_1; // @[Top.scala 152:11]
  assign n98_I_6_1_2 = n89_O_6_1_2; // @[Top.scala 152:11]
  assign n98_I_6_2_0 = n89_O_6_2_0; // @[Top.scala 152:11]
  assign n98_I_6_2_1 = n89_O_6_2_1; // @[Top.scala 152:11]
  assign n98_I_6_2_2 = n89_O_6_2_2; // @[Top.scala 152:11]
  assign n98_I_7_0_0 = n89_O_7_0_0; // @[Top.scala 152:11]
  assign n98_I_7_0_1 = n89_O_7_0_1; // @[Top.scala 152:11]
  assign n98_I_7_0_2 = n89_O_7_0_2; // @[Top.scala 152:11]
  assign n98_I_7_1_0 = n89_O_7_1_0; // @[Top.scala 152:11]
  assign n98_I_7_1_1 = n89_O_7_1_1; // @[Top.scala 152:11]
  assign n98_I_7_1_2 = n89_O_7_1_2; // @[Top.scala 152:11]
  assign n98_I_7_2_0 = n89_O_7_2_0; // @[Top.scala 152:11]
  assign n98_I_7_2_1 = n89_O_7_2_1; // @[Top.scala 152:11]
  assign n98_I_7_2_2 = n89_O_7_2_2; // @[Top.scala 152:11]
  assign n98_I_8_0_0 = n89_O_8_0_0; // @[Top.scala 152:11]
  assign n98_I_8_0_1 = n89_O_8_0_1; // @[Top.scala 152:11]
  assign n98_I_8_0_2 = n89_O_8_0_2; // @[Top.scala 152:11]
  assign n98_I_8_1_0 = n89_O_8_1_0; // @[Top.scala 152:11]
  assign n98_I_8_1_1 = n89_O_8_1_1; // @[Top.scala 152:11]
  assign n98_I_8_1_2 = n89_O_8_1_2; // @[Top.scala 152:11]
  assign n98_I_8_2_0 = n89_O_8_2_0; // @[Top.scala 152:11]
  assign n98_I_8_2_1 = n89_O_8_2_1; // @[Top.scala 152:11]
  assign n98_I_8_2_2 = n89_O_8_2_2; // @[Top.scala 152:11]
  assign n98_I_9_0_0 = n89_O_9_0_0; // @[Top.scala 152:11]
  assign n98_I_9_0_1 = n89_O_9_0_1; // @[Top.scala 152:11]
  assign n98_I_9_0_2 = n89_O_9_0_2; // @[Top.scala 152:11]
  assign n98_I_9_1_0 = n89_O_9_1_0; // @[Top.scala 152:11]
  assign n98_I_9_1_1 = n89_O_9_1_1; // @[Top.scala 152:11]
  assign n98_I_9_1_2 = n89_O_9_1_2; // @[Top.scala 152:11]
  assign n98_I_9_2_0 = n89_O_9_2_0; // @[Top.scala 152:11]
  assign n98_I_9_2_1 = n89_O_9_2_1; // @[Top.scala 152:11]
  assign n98_I_9_2_2 = n89_O_9_2_2; // @[Top.scala 152:11]
  assign n98_I_10_0_0 = n89_O_10_0_0; // @[Top.scala 152:11]
  assign n98_I_10_0_1 = n89_O_10_0_1; // @[Top.scala 152:11]
  assign n98_I_10_0_2 = n89_O_10_0_2; // @[Top.scala 152:11]
  assign n98_I_10_1_0 = n89_O_10_1_0; // @[Top.scala 152:11]
  assign n98_I_10_1_1 = n89_O_10_1_1; // @[Top.scala 152:11]
  assign n98_I_10_1_2 = n89_O_10_1_2; // @[Top.scala 152:11]
  assign n98_I_10_2_0 = n89_O_10_2_0; // @[Top.scala 152:11]
  assign n98_I_10_2_1 = n89_O_10_2_1; // @[Top.scala 152:11]
  assign n98_I_10_2_2 = n89_O_10_2_2; // @[Top.scala 152:11]
  assign n98_I_11_0_0 = n89_O_11_0_0; // @[Top.scala 152:11]
  assign n98_I_11_0_1 = n89_O_11_0_1; // @[Top.scala 152:11]
  assign n98_I_11_0_2 = n89_O_11_0_2; // @[Top.scala 152:11]
  assign n98_I_11_1_0 = n89_O_11_1_0; // @[Top.scala 152:11]
  assign n98_I_11_1_1 = n89_O_11_1_1; // @[Top.scala 152:11]
  assign n98_I_11_1_2 = n89_O_11_1_2; // @[Top.scala 152:11]
  assign n98_I_11_2_0 = n89_O_11_2_0; // @[Top.scala 152:11]
  assign n98_I_11_2_1 = n89_O_11_2_1; // @[Top.scala 152:11]
  assign n98_I_11_2_2 = n89_O_11_2_2; // @[Top.scala 152:11]
  assign n98_I_12_0_0 = n89_O_12_0_0; // @[Top.scala 152:11]
  assign n98_I_12_0_1 = n89_O_12_0_1; // @[Top.scala 152:11]
  assign n98_I_12_0_2 = n89_O_12_0_2; // @[Top.scala 152:11]
  assign n98_I_12_1_0 = n89_O_12_1_0; // @[Top.scala 152:11]
  assign n98_I_12_1_1 = n89_O_12_1_1; // @[Top.scala 152:11]
  assign n98_I_12_1_2 = n89_O_12_1_2; // @[Top.scala 152:11]
  assign n98_I_12_2_0 = n89_O_12_2_0; // @[Top.scala 152:11]
  assign n98_I_12_2_1 = n89_O_12_2_1; // @[Top.scala 152:11]
  assign n98_I_12_2_2 = n89_O_12_2_2; // @[Top.scala 152:11]
  assign n98_I_13_0_0 = n89_O_13_0_0; // @[Top.scala 152:11]
  assign n98_I_13_0_1 = n89_O_13_0_1; // @[Top.scala 152:11]
  assign n98_I_13_0_2 = n89_O_13_0_2; // @[Top.scala 152:11]
  assign n98_I_13_1_0 = n89_O_13_1_0; // @[Top.scala 152:11]
  assign n98_I_13_1_1 = n89_O_13_1_1; // @[Top.scala 152:11]
  assign n98_I_13_1_2 = n89_O_13_1_2; // @[Top.scala 152:11]
  assign n98_I_13_2_0 = n89_O_13_2_0; // @[Top.scala 152:11]
  assign n98_I_13_2_1 = n89_O_13_2_1; // @[Top.scala 152:11]
  assign n98_I_13_2_2 = n89_O_13_2_2; // @[Top.scala 152:11]
  assign n98_I_14_0_0 = n89_O_14_0_0; // @[Top.scala 152:11]
  assign n98_I_14_0_1 = n89_O_14_0_1; // @[Top.scala 152:11]
  assign n98_I_14_0_2 = n89_O_14_0_2; // @[Top.scala 152:11]
  assign n98_I_14_1_0 = n89_O_14_1_0; // @[Top.scala 152:11]
  assign n98_I_14_1_1 = n89_O_14_1_1; // @[Top.scala 152:11]
  assign n98_I_14_1_2 = n89_O_14_1_2; // @[Top.scala 152:11]
  assign n98_I_14_2_0 = n89_O_14_2_0; // @[Top.scala 152:11]
  assign n98_I_14_2_1 = n89_O_14_2_1; // @[Top.scala 152:11]
  assign n98_I_14_2_2 = n89_O_14_2_2; // @[Top.scala 152:11]
  assign n98_I_15_0_0 = n89_O_15_0_0; // @[Top.scala 152:11]
  assign n98_I_15_0_1 = n89_O_15_0_1; // @[Top.scala 152:11]
  assign n98_I_15_0_2 = n89_O_15_0_2; // @[Top.scala 152:11]
  assign n98_I_15_1_0 = n89_O_15_1_0; // @[Top.scala 152:11]
  assign n98_I_15_1_1 = n89_O_15_1_1; // @[Top.scala 152:11]
  assign n98_I_15_1_2 = n89_O_15_1_2; // @[Top.scala 152:11]
  assign n98_I_15_2_0 = n89_O_15_2_0; // @[Top.scala 152:11]
  assign n98_I_15_2_1 = n89_O_15_2_1; // @[Top.scala 152:11]
  assign n98_I_15_2_2 = n89_O_15_2_2; // @[Top.scala 152:11]
  assign n105_valid_up = n98_valid_down; // @[Top.scala 156:19]
  assign n105_I_0_0_0_0 = n98_O_0_0_0_0; // @[Top.scala 155:12]
  assign n105_I_0_0_0_1 = n98_O_0_0_0_1; // @[Top.scala 155:12]
  assign n105_I_0_0_0_2 = n98_O_0_0_0_2; // @[Top.scala 155:12]
  assign n105_I_0_0_1_0 = n98_O_0_0_1_0; // @[Top.scala 155:12]
  assign n105_I_0_0_1_1 = n98_O_0_0_1_1; // @[Top.scala 155:12]
  assign n105_I_0_0_1_2 = n98_O_0_0_1_2; // @[Top.scala 155:12]
  assign n105_I_0_0_2_0 = n98_O_0_0_2_0; // @[Top.scala 155:12]
  assign n105_I_0_0_2_1 = n98_O_0_0_2_1; // @[Top.scala 155:12]
  assign n105_I_0_0_2_2 = n98_O_0_0_2_2; // @[Top.scala 155:12]
  assign n105_I_1_0_0_0 = n98_O_1_0_0_0; // @[Top.scala 155:12]
  assign n105_I_1_0_0_1 = n98_O_1_0_0_1; // @[Top.scala 155:12]
  assign n105_I_1_0_0_2 = n98_O_1_0_0_2; // @[Top.scala 155:12]
  assign n105_I_1_0_1_0 = n98_O_1_0_1_0; // @[Top.scala 155:12]
  assign n105_I_1_0_1_1 = n98_O_1_0_1_1; // @[Top.scala 155:12]
  assign n105_I_1_0_1_2 = n98_O_1_0_1_2; // @[Top.scala 155:12]
  assign n105_I_1_0_2_0 = n98_O_1_0_2_0; // @[Top.scala 155:12]
  assign n105_I_1_0_2_1 = n98_O_1_0_2_1; // @[Top.scala 155:12]
  assign n105_I_1_0_2_2 = n98_O_1_0_2_2; // @[Top.scala 155:12]
  assign n105_I_2_0_0_0 = n98_O_2_0_0_0; // @[Top.scala 155:12]
  assign n105_I_2_0_0_1 = n98_O_2_0_0_1; // @[Top.scala 155:12]
  assign n105_I_2_0_0_2 = n98_O_2_0_0_2; // @[Top.scala 155:12]
  assign n105_I_2_0_1_0 = n98_O_2_0_1_0; // @[Top.scala 155:12]
  assign n105_I_2_0_1_1 = n98_O_2_0_1_1; // @[Top.scala 155:12]
  assign n105_I_2_0_1_2 = n98_O_2_0_1_2; // @[Top.scala 155:12]
  assign n105_I_2_0_2_0 = n98_O_2_0_2_0; // @[Top.scala 155:12]
  assign n105_I_2_0_2_1 = n98_O_2_0_2_1; // @[Top.scala 155:12]
  assign n105_I_2_0_2_2 = n98_O_2_0_2_2; // @[Top.scala 155:12]
  assign n105_I_3_0_0_0 = n98_O_3_0_0_0; // @[Top.scala 155:12]
  assign n105_I_3_0_0_1 = n98_O_3_0_0_1; // @[Top.scala 155:12]
  assign n105_I_3_0_0_2 = n98_O_3_0_0_2; // @[Top.scala 155:12]
  assign n105_I_3_0_1_0 = n98_O_3_0_1_0; // @[Top.scala 155:12]
  assign n105_I_3_0_1_1 = n98_O_3_0_1_1; // @[Top.scala 155:12]
  assign n105_I_3_0_1_2 = n98_O_3_0_1_2; // @[Top.scala 155:12]
  assign n105_I_3_0_2_0 = n98_O_3_0_2_0; // @[Top.scala 155:12]
  assign n105_I_3_0_2_1 = n98_O_3_0_2_1; // @[Top.scala 155:12]
  assign n105_I_3_0_2_2 = n98_O_3_0_2_2; // @[Top.scala 155:12]
  assign n105_I_4_0_0_0 = n98_O_4_0_0_0; // @[Top.scala 155:12]
  assign n105_I_4_0_0_1 = n98_O_4_0_0_1; // @[Top.scala 155:12]
  assign n105_I_4_0_0_2 = n98_O_4_0_0_2; // @[Top.scala 155:12]
  assign n105_I_4_0_1_0 = n98_O_4_0_1_0; // @[Top.scala 155:12]
  assign n105_I_4_0_1_1 = n98_O_4_0_1_1; // @[Top.scala 155:12]
  assign n105_I_4_0_1_2 = n98_O_4_0_1_2; // @[Top.scala 155:12]
  assign n105_I_4_0_2_0 = n98_O_4_0_2_0; // @[Top.scala 155:12]
  assign n105_I_4_0_2_1 = n98_O_4_0_2_1; // @[Top.scala 155:12]
  assign n105_I_4_0_2_2 = n98_O_4_0_2_2; // @[Top.scala 155:12]
  assign n105_I_5_0_0_0 = n98_O_5_0_0_0; // @[Top.scala 155:12]
  assign n105_I_5_0_0_1 = n98_O_5_0_0_1; // @[Top.scala 155:12]
  assign n105_I_5_0_0_2 = n98_O_5_0_0_2; // @[Top.scala 155:12]
  assign n105_I_5_0_1_0 = n98_O_5_0_1_0; // @[Top.scala 155:12]
  assign n105_I_5_0_1_1 = n98_O_5_0_1_1; // @[Top.scala 155:12]
  assign n105_I_5_0_1_2 = n98_O_5_0_1_2; // @[Top.scala 155:12]
  assign n105_I_5_0_2_0 = n98_O_5_0_2_0; // @[Top.scala 155:12]
  assign n105_I_5_0_2_1 = n98_O_5_0_2_1; // @[Top.scala 155:12]
  assign n105_I_5_0_2_2 = n98_O_5_0_2_2; // @[Top.scala 155:12]
  assign n105_I_6_0_0_0 = n98_O_6_0_0_0; // @[Top.scala 155:12]
  assign n105_I_6_0_0_1 = n98_O_6_0_0_1; // @[Top.scala 155:12]
  assign n105_I_6_0_0_2 = n98_O_6_0_0_2; // @[Top.scala 155:12]
  assign n105_I_6_0_1_0 = n98_O_6_0_1_0; // @[Top.scala 155:12]
  assign n105_I_6_0_1_1 = n98_O_6_0_1_1; // @[Top.scala 155:12]
  assign n105_I_6_0_1_2 = n98_O_6_0_1_2; // @[Top.scala 155:12]
  assign n105_I_6_0_2_0 = n98_O_6_0_2_0; // @[Top.scala 155:12]
  assign n105_I_6_0_2_1 = n98_O_6_0_2_1; // @[Top.scala 155:12]
  assign n105_I_6_0_2_2 = n98_O_6_0_2_2; // @[Top.scala 155:12]
  assign n105_I_7_0_0_0 = n98_O_7_0_0_0; // @[Top.scala 155:12]
  assign n105_I_7_0_0_1 = n98_O_7_0_0_1; // @[Top.scala 155:12]
  assign n105_I_7_0_0_2 = n98_O_7_0_0_2; // @[Top.scala 155:12]
  assign n105_I_7_0_1_0 = n98_O_7_0_1_0; // @[Top.scala 155:12]
  assign n105_I_7_0_1_1 = n98_O_7_0_1_1; // @[Top.scala 155:12]
  assign n105_I_7_0_1_2 = n98_O_7_0_1_2; // @[Top.scala 155:12]
  assign n105_I_7_0_2_0 = n98_O_7_0_2_0; // @[Top.scala 155:12]
  assign n105_I_7_0_2_1 = n98_O_7_0_2_1; // @[Top.scala 155:12]
  assign n105_I_7_0_2_2 = n98_O_7_0_2_2; // @[Top.scala 155:12]
  assign n105_I_8_0_0_0 = n98_O_8_0_0_0; // @[Top.scala 155:12]
  assign n105_I_8_0_0_1 = n98_O_8_0_0_1; // @[Top.scala 155:12]
  assign n105_I_8_0_0_2 = n98_O_8_0_0_2; // @[Top.scala 155:12]
  assign n105_I_8_0_1_0 = n98_O_8_0_1_0; // @[Top.scala 155:12]
  assign n105_I_8_0_1_1 = n98_O_8_0_1_1; // @[Top.scala 155:12]
  assign n105_I_8_0_1_2 = n98_O_8_0_1_2; // @[Top.scala 155:12]
  assign n105_I_8_0_2_0 = n98_O_8_0_2_0; // @[Top.scala 155:12]
  assign n105_I_8_0_2_1 = n98_O_8_0_2_1; // @[Top.scala 155:12]
  assign n105_I_8_0_2_2 = n98_O_8_0_2_2; // @[Top.scala 155:12]
  assign n105_I_9_0_0_0 = n98_O_9_0_0_0; // @[Top.scala 155:12]
  assign n105_I_9_0_0_1 = n98_O_9_0_0_1; // @[Top.scala 155:12]
  assign n105_I_9_0_0_2 = n98_O_9_0_0_2; // @[Top.scala 155:12]
  assign n105_I_9_0_1_0 = n98_O_9_0_1_0; // @[Top.scala 155:12]
  assign n105_I_9_0_1_1 = n98_O_9_0_1_1; // @[Top.scala 155:12]
  assign n105_I_9_0_1_2 = n98_O_9_0_1_2; // @[Top.scala 155:12]
  assign n105_I_9_0_2_0 = n98_O_9_0_2_0; // @[Top.scala 155:12]
  assign n105_I_9_0_2_1 = n98_O_9_0_2_1; // @[Top.scala 155:12]
  assign n105_I_9_0_2_2 = n98_O_9_0_2_2; // @[Top.scala 155:12]
  assign n105_I_10_0_0_0 = n98_O_10_0_0_0; // @[Top.scala 155:12]
  assign n105_I_10_0_0_1 = n98_O_10_0_0_1; // @[Top.scala 155:12]
  assign n105_I_10_0_0_2 = n98_O_10_0_0_2; // @[Top.scala 155:12]
  assign n105_I_10_0_1_0 = n98_O_10_0_1_0; // @[Top.scala 155:12]
  assign n105_I_10_0_1_1 = n98_O_10_0_1_1; // @[Top.scala 155:12]
  assign n105_I_10_0_1_2 = n98_O_10_0_1_2; // @[Top.scala 155:12]
  assign n105_I_10_0_2_0 = n98_O_10_0_2_0; // @[Top.scala 155:12]
  assign n105_I_10_0_2_1 = n98_O_10_0_2_1; // @[Top.scala 155:12]
  assign n105_I_10_0_2_2 = n98_O_10_0_2_2; // @[Top.scala 155:12]
  assign n105_I_11_0_0_0 = n98_O_11_0_0_0; // @[Top.scala 155:12]
  assign n105_I_11_0_0_1 = n98_O_11_0_0_1; // @[Top.scala 155:12]
  assign n105_I_11_0_0_2 = n98_O_11_0_0_2; // @[Top.scala 155:12]
  assign n105_I_11_0_1_0 = n98_O_11_0_1_0; // @[Top.scala 155:12]
  assign n105_I_11_0_1_1 = n98_O_11_0_1_1; // @[Top.scala 155:12]
  assign n105_I_11_0_1_2 = n98_O_11_0_1_2; // @[Top.scala 155:12]
  assign n105_I_11_0_2_0 = n98_O_11_0_2_0; // @[Top.scala 155:12]
  assign n105_I_11_0_2_1 = n98_O_11_0_2_1; // @[Top.scala 155:12]
  assign n105_I_11_0_2_2 = n98_O_11_0_2_2; // @[Top.scala 155:12]
  assign n105_I_12_0_0_0 = n98_O_12_0_0_0; // @[Top.scala 155:12]
  assign n105_I_12_0_0_1 = n98_O_12_0_0_1; // @[Top.scala 155:12]
  assign n105_I_12_0_0_2 = n98_O_12_0_0_2; // @[Top.scala 155:12]
  assign n105_I_12_0_1_0 = n98_O_12_0_1_0; // @[Top.scala 155:12]
  assign n105_I_12_0_1_1 = n98_O_12_0_1_1; // @[Top.scala 155:12]
  assign n105_I_12_0_1_2 = n98_O_12_0_1_2; // @[Top.scala 155:12]
  assign n105_I_12_0_2_0 = n98_O_12_0_2_0; // @[Top.scala 155:12]
  assign n105_I_12_0_2_1 = n98_O_12_0_2_1; // @[Top.scala 155:12]
  assign n105_I_12_0_2_2 = n98_O_12_0_2_2; // @[Top.scala 155:12]
  assign n105_I_13_0_0_0 = n98_O_13_0_0_0; // @[Top.scala 155:12]
  assign n105_I_13_0_0_1 = n98_O_13_0_0_1; // @[Top.scala 155:12]
  assign n105_I_13_0_0_2 = n98_O_13_0_0_2; // @[Top.scala 155:12]
  assign n105_I_13_0_1_0 = n98_O_13_0_1_0; // @[Top.scala 155:12]
  assign n105_I_13_0_1_1 = n98_O_13_0_1_1; // @[Top.scala 155:12]
  assign n105_I_13_0_1_2 = n98_O_13_0_1_2; // @[Top.scala 155:12]
  assign n105_I_13_0_2_0 = n98_O_13_0_2_0; // @[Top.scala 155:12]
  assign n105_I_13_0_2_1 = n98_O_13_0_2_1; // @[Top.scala 155:12]
  assign n105_I_13_0_2_2 = n98_O_13_0_2_2; // @[Top.scala 155:12]
  assign n105_I_14_0_0_0 = n98_O_14_0_0_0; // @[Top.scala 155:12]
  assign n105_I_14_0_0_1 = n98_O_14_0_0_1; // @[Top.scala 155:12]
  assign n105_I_14_0_0_2 = n98_O_14_0_0_2; // @[Top.scala 155:12]
  assign n105_I_14_0_1_0 = n98_O_14_0_1_0; // @[Top.scala 155:12]
  assign n105_I_14_0_1_1 = n98_O_14_0_1_1; // @[Top.scala 155:12]
  assign n105_I_14_0_1_2 = n98_O_14_0_1_2; // @[Top.scala 155:12]
  assign n105_I_14_0_2_0 = n98_O_14_0_2_0; // @[Top.scala 155:12]
  assign n105_I_14_0_2_1 = n98_O_14_0_2_1; // @[Top.scala 155:12]
  assign n105_I_14_0_2_2 = n98_O_14_0_2_2; // @[Top.scala 155:12]
  assign n105_I_15_0_0_0 = n98_O_15_0_0_0; // @[Top.scala 155:12]
  assign n105_I_15_0_0_1 = n98_O_15_0_0_1; // @[Top.scala 155:12]
  assign n105_I_15_0_0_2 = n98_O_15_0_0_2; // @[Top.scala 155:12]
  assign n105_I_15_0_1_0 = n98_O_15_0_1_0; // @[Top.scala 155:12]
  assign n105_I_15_0_1_1 = n98_O_15_0_1_1; // @[Top.scala 155:12]
  assign n105_I_15_0_1_2 = n98_O_15_0_1_2; // @[Top.scala 155:12]
  assign n105_I_15_0_2_0 = n98_O_15_0_2_0; // @[Top.scala 155:12]
  assign n105_I_15_0_2_1 = n98_O_15_0_2_1; // @[Top.scala 155:12]
  assign n105_I_15_0_2_2 = n98_O_15_0_2_2; // @[Top.scala 155:12]
  assign n147_clock = clock;
  assign n147_reset = reset;
  assign n147_valid_up = n105_valid_down; // @[Top.scala 159:19]
  assign n147_I_0_0_0 = n105_O_0_0_0; // @[Top.scala 158:12]
  assign n147_I_0_0_1 = n105_O_0_0_1; // @[Top.scala 158:12]
  assign n147_I_0_0_2 = n105_O_0_0_2; // @[Top.scala 158:12]
  assign n147_I_0_1_0 = n105_O_0_1_0; // @[Top.scala 158:12]
  assign n147_I_0_1_1 = n105_O_0_1_1; // @[Top.scala 158:12]
  assign n147_I_0_1_2 = n105_O_0_1_2; // @[Top.scala 158:12]
  assign n147_I_0_2_0 = n105_O_0_2_0; // @[Top.scala 158:12]
  assign n147_I_0_2_1 = n105_O_0_2_1; // @[Top.scala 158:12]
  assign n147_I_0_2_2 = n105_O_0_2_2; // @[Top.scala 158:12]
  assign n147_I_1_0_0 = n105_O_1_0_0; // @[Top.scala 158:12]
  assign n147_I_1_0_1 = n105_O_1_0_1; // @[Top.scala 158:12]
  assign n147_I_1_0_2 = n105_O_1_0_2; // @[Top.scala 158:12]
  assign n147_I_1_1_0 = n105_O_1_1_0; // @[Top.scala 158:12]
  assign n147_I_1_1_1 = n105_O_1_1_1; // @[Top.scala 158:12]
  assign n147_I_1_1_2 = n105_O_1_1_2; // @[Top.scala 158:12]
  assign n147_I_1_2_0 = n105_O_1_2_0; // @[Top.scala 158:12]
  assign n147_I_1_2_1 = n105_O_1_2_1; // @[Top.scala 158:12]
  assign n147_I_1_2_2 = n105_O_1_2_2; // @[Top.scala 158:12]
  assign n147_I_2_0_0 = n105_O_2_0_0; // @[Top.scala 158:12]
  assign n147_I_2_0_1 = n105_O_2_0_1; // @[Top.scala 158:12]
  assign n147_I_2_0_2 = n105_O_2_0_2; // @[Top.scala 158:12]
  assign n147_I_2_1_0 = n105_O_2_1_0; // @[Top.scala 158:12]
  assign n147_I_2_1_1 = n105_O_2_1_1; // @[Top.scala 158:12]
  assign n147_I_2_1_2 = n105_O_2_1_2; // @[Top.scala 158:12]
  assign n147_I_2_2_0 = n105_O_2_2_0; // @[Top.scala 158:12]
  assign n147_I_2_2_1 = n105_O_2_2_1; // @[Top.scala 158:12]
  assign n147_I_2_2_2 = n105_O_2_2_2; // @[Top.scala 158:12]
  assign n147_I_3_0_0 = n105_O_3_0_0; // @[Top.scala 158:12]
  assign n147_I_3_0_1 = n105_O_3_0_1; // @[Top.scala 158:12]
  assign n147_I_3_0_2 = n105_O_3_0_2; // @[Top.scala 158:12]
  assign n147_I_3_1_0 = n105_O_3_1_0; // @[Top.scala 158:12]
  assign n147_I_3_1_1 = n105_O_3_1_1; // @[Top.scala 158:12]
  assign n147_I_3_1_2 = n105_O_3_1_2; // @[Top.scala 158:12]
  assign n147_I_3_2_0 = n105_O_3_2_0; // @[Top.scala 158:12]
  assign n147_I_3_2_1 = n105_O_3_2_1; // @[Top.scala 158:12]
  assign n147_I_3_2_2 = n105_O_3_2_2; // @[Top.scala 158:12]
  assign n147_I_4_0_0 = n105_O_4_0_0; // @[Top.scala 158:12]
  assign n147_I_4_0_1 = n105_O_4_0_1; // @[Top.scala 158:12]
  assign n147_I_4_0_2 = n105_O_4_0_2; // @[Top.scala 158:12]
  assign n147_I_4_1_0 = n105_O_4_1_0; // @[Top.scala 158:12]
  assign n147_I_4_1_1 = n105_O_4_1_1; // @[Top.scala 158:12]
  assign n147_I_4_1_2 = n105_O_4_1_2; // @[Top.scala 158:12]
  assign n147_I_4_2_0 = n105_O_4_2_0; // @[Top.scala 158:12]
  assign n147_I_4_2_1 = n105_O_4_2_1; // @[Top.scala 158:12]
  assign n147_I_4_2_2 = n105_O_4_2_2; // @[Top.scala 158:12]
  assign n147_I_5_0_0 = n105_O_5_0_0; // @[Top.scala 158:12]
  assign n147_I_5_0_1 = n105_O_5_0_1; // @[Top.scala 158:12]
  assign n147_I_5_0_2 = n105_O_5_0_2; // @[Top.scala 158:12]
  assign n147_I_5_1_0 = n105_O_5_1_0; // @[Top.scala 158:12]
  assign n147_I_5_1_1 = n105_O_5_1_1; // @[Top.scala 158:12]
  assign n147_I_5_1_2 = n105_O_5_1_2; // @[Top.scala 158:12]
  assign n147_I_5_2_0 = n105_O_5_2_0; // @[Top.scala 158:12]
  assign n147_I_5_2_1 = n105_O_5_2_1; // @[Top.scala 158:12]
  assign n147_I_5_2_2 = n105_O_5_2_2; // @[Top.scala 158:12]
  assign n147_I_6_0_0 = n105_O_6_0_0; // @[Top.scala 158:12]
  assign n147_I_6_0_1 = n105_O_6_0_1; // @[Top.scala 158:12]
  assign n147_I_6_0_2 = n105_O_6_0_2; // @[Top.scala 158:12]
  assign n147_I_6_1_0 = n105_O_6_1_0; // @[Top.scala 158:12]
  assign n147_I_6_1_1 = n105_O_6_1_1; // @[Top.scala 158:12]
  assign n147_I_6_1_2 = n105_O_6_1_2; // @[Top.scala 158:12]
  assign n147_I_6_2_0 = n105_O_6_2_0; // @[Top.scala 158:12]
  assign n147_I_6_2_1 = n105_O_6_2_1; // @[Top.scala 158:12]
  assign n147_I_6_2_2 = n105_O_6_2_2; // @[Top.scala 158:12]
  assign n147_I_7_0_0 = n105_O_7_0_0; // @[Top.scala 158:12]
  assign n147_I_7_0_1 = n105_O_7_0_1; // @[Top.scala 158:12]
  assign n147_I_7_0_2 = n105_O_7_0_2; // @[Top.scala 158:12]
  assign n147_I_7_1_0 = n105_O_7_1_0; // @[Top.scala 158:12]
  assign n147_I_7_1_1 = n105_O_7_1_1; // @[Top.scala 158:12]
  assign n147_I_7_1_2 = n105_O_7_1_2; // @[Top.scala 158:12]
  assign n147_I_7_2_0 = n105_O_7_2_0; // @[Top.scala 158:12]
  assign n147_I_7_2_1 = n105_O_7_2_1; // @[Top.scala 158:12]
  assign n147_I_7_2_2 = n105_O_7_2_2; // @[Top.scala 158:12]
  assign n147_I_8_0_0 = n105_O_8_0_0; // @[Top.scala 158:12]
  assign n147_I_8_0_1 = n105_O_8_0_1; // @[Top.scala 158:12]
  assign n147_I_8_0_2 = n105_O_8_0_2; // @[Top.scala 158:12]
  assign n147_I_8_1_0 = n105_O_8_1_0; // @[Top.scala 158:12]
  assign n147_I_8_1_1 = n105_O_8_1_1; // @[Top.scala 158:12]
  assign n147_I_8_1_2 = n105_O_8_1_2; // @[Top.scala 158:12]
  assign n147_I_8_2_0 = n105_O_8_2_0; // @[Top.scala 158:12]
  assign n147_I_8_2_1 = n105_O_8_2_1; // @[Top.scala 158:12]
  assign n147_I_8_2_2 = n105_O_8_2_2; // @[Top.scala 158:12]
  assign n147_I_9_0_0 = n105_O_9_0_0; // @[Top.scala 158:12]
  assign n147_I_9_0_1 = n105_O_9_0_1; // @[Top.scala 158:12]
  assign n147_I_9_0_2 = n105_O_9_0_2; // @[Top.scala 158:12]
  assign n147_I_9_1_0 = n105_O_9_1_0; // @[Top.scala 158:12]
  assign n147_I_9_1_1 = n105_O_9_1_1; // @[Top.scala 158:12]
  assign n147_I_9_1_2 = n105_O_9_1_2; // @[Top.scala 158:12]
  assign n147_I_9_2_0 = n105_O_9_2_0; // @[Top.scala 158:12]
  assign n147_I_9_2_1 = n105_O_9_2_1; // @[Top.scala 158:12]
  assign n147_I_9_2_2 = n105_O_9_2_2; // @[Top.scala 158:12]
  assign n147_I_10_0_0 = n105_O_10_0_0; // @[Top.scala 158:12]
  assign n147_I_10_0_1 = n105_O_10_0_1; // @[Top.scala 158:12]
  assign n147_I_10_0_2 = n105_O_10_0_2; // @[Top.scala 158:12]
  assign n147_I_10_1_0 = n105_O_10_1_0; // @[Top.scala 158:12]
  assign n147_I_10_1_1 = n105_O_10_1_1; // @[Top.scala 158:12]
  assign n147_I_10_1_2 = n105_O_10_1_2; // @[Top.scala 158:12]
  assign n147_I_10_2_0 = n105_O_10_2_0; // @[Top.scala 158:12]
  assign n147_I_10_2_1 = n105_O_10_2_1; // @[Top.scala 158:12]
  assign n147_I_10_2_2 = n105_O_10_2_2; // @[Top.scala 158:12]
  assign n147_I_11_0_0 = n105_O_11_0_0; // @[Top.scala 158:12]
  assign n147_I_11_0_1 = n105_O_11_0_1; // @[Top.scala 158:12]
  assign n147_I_11_0_2 = n105_O_11_0_2; // @[Top.scala 158:12]
  assign n147_I_11_1_0 = n105_O_11_1_0; // @[Top.scala 158:12]
  assign n147_I_11_1_1 = n105_O_11_1_1; // @[Top.scala 158:12]
  assign n147_I_11_1_2 = n105_O_11_1_2; // @[Top.scala 158:12]
  assign n147_I_11_2_0 = n105_O_11_2_0; // @[Top.scala 158:12]
  assign n147_I_11_2_1 = n105_O_11_2_1; // @[Top.scala 158:12]
  assign n147_I_11_2_2 = n105_O_11_2_2; // @[Top.scala 158:12]
  assign n147_I_12_0_0 = n105_O_12_0_0; // @[Top.scala 158:12]
  assign n147_I_12_0_1 = n105_O_12_0_1; // @[Top.scala 158:12]
  assign n147_I_12_0_2 = n105_O_12_0_2; // @[Top.scala 158:12]
  assign n147_I_12_1_0 = n105_O_12_1_0; // @[Top.scala 158:12]
  assign n147_I_12_1_1 = n105_O_12_1_1; // @[Top.scala 158:12]
  assign n147_I_12_1_2 = n105_O_12_1_2; // @[Top.scala 158:12]
  assign n147_I_12_2_0 = n105_O_12_2_0; // @[Top.scala 158:12]
  assign n147_I_12_2_1 = n105_O_12_2_1; // @[Top.scala 158:12]
  assign n147_I_12_2_2 = n105_O_12_2_2; // @[Top.scala 158:12]
  assign n147_I_13_0_0 = n105_O_13_0_0; // @[Top.scala 158:12]
  assign n147_I_13_0_1 = n105_O_13_0_1; // @[Top.scala 158:12]
  assign n147_I_13_0_2 = n105_O_13_0_2; // @[Top.scala 158:12]
  assign n147_I_13_1_0 = n105_O_13_1_0; // @[Top.scala 158:12]
  assign n147_I_13_1_1 = n105_O_13_1_1; // @[Top.scala 158:12]
  assign n147_I_13_1_2 = n105_O_13_1_2; // @[Top.scala 158:12]
  assign n147_I_13_2_0 = n105_O_13_2_0; // @[Top.scala 158:12]
  assign n147_I_13_2_1 = n105_O_13_2_1; // @[Top.scala 158:12]
  assign n147_I_13_2_2 = n105_O_13_2_2; // @[Top.scala 158:12]
  assign n147_I_14_0_0 = n105_O_14_0_0; // @[Top.scala 158:12]
  assign n147_I_14_0_1 = n105_O_14_0_1; // @[Top.scala 158:12]
  assign n147_I_14_0_2 = n105_O_14_0_2; // @[Top.scala 158:12]
  assign n147_I_14_1_0 = n105_O_14_1_0; // @[Top.scala 158:12]
  assign n147_I_14_1_1 = n105_O_14_1_1; // @[Top.scala 158:12]
  assign n147_I_14_1_2 = n105_O_14_1_2; // @[Top.scala 158:12]
  assign n147_I_14_2_0 = n105_O_14_2_0; // @[Top.scala 158:12]
  assign n147_I_14_2_1 = n105_O_14_2_1; // @[Top.scala 158:12]
  assign n147_I_14_2_2 = n105_O_14_2_2; // @[Top.scala 158:12]
  assign n147_I_15_0_0 = n105_O_15_0_0; // @[Top.scala 158:12]
  assign n147_I_15_0_1 = n105_O_15_0_1; // @[Top.scala 158:12]
  assign n147_I_15_0_2 = n105_O_15_0_2; // @[Top.scala 158:12]
  assign n147_I_15_1_0 = n105_O_15_1_0; // @[Top.scala 158:12]
  assign n147_I_15_1_1 = n105_O_15_1_1; // @[Top.scala 158:12]
  assign n147_I_15_1_2 = n105_O_15_1_2; // @[Top.scala 158:12]
  assign n147_I_15_2_0 = n105_O_15_2_0; // @[Top.scala 158:12]
  assign n147_I_15_2_1 = n105_O_15_2_1; // @[Top.scala 158:12]
  assign n147_I_15_2_2 = n105_O_15_2_2; // @[Top.scala 158:12]
  assign n148_valid_up = n147_valid_down; // @[Top.scala 162:19]
  assign n148_I_0_0_0 = n147_O_0_0_0; // @[Top.scala 161:12]
  assign n148_I_1_0_0 = n147_O_1_0_0; // @[Top.scala 161:12]
  assign n148_I_2_0_0 = n147_O_2_0_0; // @[Top.scala 161:12]
  assign n148_I_3_0_0 = n147_O_3_0_0; // @[Top.scala 161:12]
  assign n148_I_4_0_0 = n147_O_4_0_0; // @[Top.scala 161:12]
  assign n148_I_5_0_0 = n147_O_5_0_0; // @[Top.scala 161:12]
  assign n148_I_6_0_0 = n147_O_6_0_0; // @[Top.scala 161:12]
  assign n148_I_7_0_0 = n147_O_7_0_0; // @[Top.scala 161:12]
  assign n148_I_8_0_0 = n147_O_8_0_0; // @[Top.scala 161:12]
  assign n148_I_9_0_0 = n147_O_9_0_0; // @[Top.scala 161:12]
  assign n148_I_10_0_0 = n147_O_10_0_0; // @[Top.scala 161:12]
  assign n148_I_11_0_0 = n147_O_11_0_0; // @[Top.scala 161:12]
  assign n148_I_12_0_0 = n147_O_12_0_0; // @[Top.scala 161:12]
  assign n148_I_13_0_0 = n147_O_13_0_0; // @[Top.scala 161:12]
  assign n148_I_14_0_0 = n147_O_14_0_0; // @[Top.scala 161:12]
  assign n148_I_15_0_0 = n147_O_15_0_0; // @[Top.scala 161:12]
  assign n149_valid_up = n148_valid_down; // @[Top.scala 165:19]
  assign n149_I_0_0 = n148_O_0_0; // @[Top.scala 164:12]
  assign n149_I_1_0 = n148_O_1_0; // @[Top.scala 164:12]
  assign n149_I_2_0 = n148_O_2_0; // @[Top.scala 164:12]
  assign n149_I_3_0 = n148_O_3_0; // @[Top.scala 164:12]
  assign n149_I_4_0 = n148_O_4_0; // @[Top.scala 164:12]
  assign n149_I_5_0 = n148_O_5_0; // @[Top.scala 164:12]
  assign n149_I_6_0 = n148_O_6_0; // @[Top.scala 164:12]
  assign n149_I_7_0 = n148_O_7_0; // @[Top.scala 164:12]
  assign n149_I_8_0 = n148_O_8_0; // @[Top.scala 164:12]
  assign n149_I_9_0 = n148_O_9_0; // @[Top.scala 164:12]
  assign n149_I_10_0 = n148_O_10_0; // @[Top.scala 164:12]
  assign n149_I_11_0 = n148_O_11_0; // @[Top.scala 164:12]
  assign n149_I_12_0 = n148_O_12_0; // @[Top.scala 164:12]
  assign n149_I_13_0 = n148_O_13_0; // @[Top.scala 164:12]
  assign n149_I_14_0 = n148_O_14_0; // @[Top.scala 164:12]
  assign n149_I_15_0 = n148_O_15_0; // @[Top.scala 164:12]
  assign n150_clock = clock;
  assign n150_reset = reset;
  assign n150_valid_up = n149_valid_down; // @[Top.scala 168:19]
  assign n150_I_0 = n149_O_0; // @[Top.scala 167:12]
  assign n150_I_1 = n149_O_1; // @[Top.scala 167:12]
  assign n150_I_2 = n149_O_2; // @[Top.scala 167:12]
  assign n150_I_3 = n149_O_3; // @[Top.scala 167:12]
  assign n150_I_4 = n149_O_4; // @[Top.scala 167:12]
  assign n150_I_5 = n149_O_5; // @[Top.scala 167:12]
  assign n150_I_6 = n149_O_6; // @[Top.scala 167:12]
  assign n150_I_7 = n149_O_7; // @[Top.scala 167:12]
  assign n150_I_8 = n149_O_8; // @[Top.scala 167:12]
  assign n150_I_9 = n149_O_9; // @[Top.scala 167:12]
  assign n150_I_10 = n149_O_10; // @[Top.scala 167:12]
  assign n150_I_11 = n149_O_11; // @[Top.scala 167:12]
  assign n150_I_12 = n149_O_12; // @[Top.scala 167:12]
  assign n150_I_13 = n149_O_13; // @[Top.scala 167:12]
  assign n150_I_14 = n149_O_14; // @[Top.scala 167:12]
  assign n150_I_15 = n149_O_15; // @[Top.scala 167:12]
  assign n151_clock = clock;
  assign n151_valid_up = n150_valid_down; // @[Top.scala 171:19]
  assign n151_I_0 = n150_O_0; // @[Top.scala 170:12]
  assign n151_I_1 = n150_O_1; // @[Top.scala 170:12]
  assign n151_I_2 = n150_O_2; // @[Top.scala 170:12]
  assign n151_I_3 = n150_O_3; // @[Top.scala 170:12]
  assign n151_I_4 = n150_O_4; // @[Top.scala 170:12]
  assign n151_I_5 = n150_O_5; // @[Top.scala 170:12]
  assign n151_I_6 = n150_O_6; // @[Top.scala 170:12]
  assign n151_I_7 = n150_O_7; // @[Top.scala 170:12]
  assign n151_I_8 = n150_O_8; // @[Top.scala 170:12]
  assign n151_I_9 = n150_O_9; // @[Top.scala 170:12]
  assign n151_I_10 = n150_O_10; // @[Top.scala 170:12]
  assign n151_I_11 = n150_O_11; // @[Top.scala 170:12]
  assign n151_I_12 = n150_O_12; // @[Top.scala 170:12]
  assign n151_I_13 = n150_O_13; // @[Top.scala 170:12]
  assign n151_I_14 = n150_O_14; // @[Top.scala 170:12]
  assign n151_I_15 = n150_O_15; // @[Top.scala 170:12]
  assign n152_valid_up = n151_valid_down & n150_valid_down; // @[Top.scala 175:19]
  assign n152_I0_0 = n151_O_0; // @[Top.scala 173:13]
  assign n152_I0_1 = n151_O_1; // @[Top.scala 173:13]
  assign n152_I0_2 = n151_O_2; // @[Top.scala 173:13]
  assign n152_I0_3 = n151_O_3; // @[Top.scala 173:13]
  assign n152_I0_4 = n151_O_4; // @[Top.scala 173:13]
  assign n152_I0_5 = n151_O_5; // @[Top.scala 173:13]
  assign n152_I0_6 = n151_O_6; // @[Top.scala 173:13]
  assign n152_I0_7 = n151_O_7; // @[Top.scala 173:13]
  assign n152_I0_8 = n151_O_8; // @[Top.scala 173:13]
  assign n152_I0_9 = n151_O_9; // @[Top.scala 173:13]
  assign n152_I0_10 = n151_O_10; // @[Top.scala 173:13]
  assign n152_I0_11 = n151_O_11; // @[Top.scala 173:13]
  assign n152_I0_12 = n151_O_12; // @[Top.scala 173:13]
  assign n152_I0_13 = n151_O_13; // @[Top.scala 173:13]
  assign n152_I0_14 = n151_O_14; // @[Top.scala 173:13]
  assign n152_I0_15 = n151_O_15; // @[Top.scala 173:13]
  assign n152_I1_0 = n150_O_0; // @[Top.scala 174:13]
  assign n152_I1_1 = n150_O_1; // @[Top.scala 174:13]
  assign n152_I1_2 = n150_O_2; // @[Top.scala 174:13]
  assign n152_I1_3 = n150_O_3; // @[Top.scala 174:13]
  assign n152_I1_4 = n150_O_4; // @[Top.scala 174:13]
  assign n152_I1_5 = n150_O_5; // @[Top.scala 174:13]
  assign n152_I1_6 = n150_O_6; // @[Top.scala 174:13]
  assign n152_I1_7 = n150_O_7; // @[Top.scala 174:13]
  assign n152_I1_8 = n150_O_8; // @[Top.scala 174:13]
  assign n152_I1_9 = n150_O_9; // @[Top.scala 174:13]
  assign n152_I1_10 = n150_O_10; // @[Top.scala 174:13]
  assign n152_I1_11 = n150_O_11; // @[Top.scala 174:13]
  assign n152_I1_12 = n150_O_12; // @[Top.scala 174:13]
  assign n152_I1_13 = n150_O_13; // @[Top.scala 174:13]
  assign n152_I1_14 = n150_O_14; // @[Top.scala 174:13]
  assign n152_I1_15 = n150_O_15; // @[Top.scala 174:13]
  assign n161_valid_up = n152_valid_down; // @[Top.scala 178:19]
  assign n161_I_0_0 = n152_O_0_0; // @[Top.scala 177:12]
  assign n161_I_0_1 = n152_O_0_1; // @[Top.scala 177:12]
  assign n161_I_1_0 = n152_O_1_0; // @[Top.scala 177:12]
  assign n161_I_1_1 = n152_O_1_1; // @[Top.scala 177:12]
  assign n161_I_2_0 = n152_O_2_0; // @[Top.scala 177:12]
  assign n161_I_2_1 = n152_O_2_1; // @[Top.scala 177:12]
  assign n161_I_3_0 = n152_O_3_0; // @[Top.scala 177:12]
  assign n161_I_3_1 = n152_O_3_1; // @[Top.scala 177:12]
  assign n161_I_4_0 = n152_O_4_0; // @[Top.scala 177:12]
  assign n161_I_4_1 = n152_O_4_1; // @[Top.scala 177:12]
  assign n161_I_5_0 = n152_O_5_0; // @[Top.scala 177:12]
  assign n161_I_5_1 = n152_O_5_1; // @[Top.scala 177:12]
  assign n161_I_6_0 = n152_O_6_0; // @[Top.scala 177:12]
  assign n161_I_6_1 = n152_O_6_1; // @[Top.scala 177:12]
  assign n161_I_7_0 = n152_O_7_0; // @[Top.scala 177:12]
  assign n161_I_7_1 = n152_O_7_1; // @[Top.scala 177:12]
  assign n161_I_8_0 = n152_O_8_0; // @[Top.scala 177:12]
  assign n161_I_8_1 = n152_O_8_1; // @[Top.scala 177:12]
  assign n161_I_9_0 = n152_O_9_0; // @[Top.scala 177:12]
  assign n161_I_9_1 = n152_O_9_1; // @[Top.scala 177:12]
  assign n161_I_10_0 = n152_O_10_0; // @[Top.scala 177:12]
  assign n161_I_10_1 = n152_O_10_1; // @[Top.scala 177:12]
  assign n161_I_11_0 = n152_O_11_0; // @[Top.scala 177:12]
  assign n161_I_11_1 = n152_O_11_1; // @[Top.scala 177:12]
  assign n161_I_12_0 = n152_O_12_0; // @[Top.scala 177:12]
  assign n161_I_12_1 = n152_O_12_1; // @[Top.scala 177:12]
  assign n161_I_13_0 = n152_O_13_0; // @[Top.scala 177:12]
  assign n161_I_13_1 = n152_O_13_1; // @[Top.scala 177:12]
  assign n161_I_14_0 = n152_O_14_0; // @[Top.scala 177:12]
  assign n161_I_14_1 = n152_O_14_1; // @[Top.scala 177:12]
  assign n161_I_15_0 = n152_O_15_0; // @[Top.scala 177:12]
  assign n161_I_15_1 = n152_O_15_1; // @[Top.scala 177:12]
  assign n168_valid_up = n161_valid_down; // @[Top.scala 181:19]
  assign n168_I_0_0_0 = n161_O_0_0_0; // @[Top.scala 180:12]
  assign n168_I_0_0_1 = n161_O_0_0_1; // @[Top.scala 180:12]
  assign n168_I_1_0_0 = n161_O_1_0_0; // @[Top.scala 180:12]
  assign n168_I_1_0_1 = n161_O_1_0_1; // @[Top.scala 180:12]
  assign n168_I_2_0_0 = n161_O_2_0_0; // @[Top.scala 180:12]
  assign n168_I_2_0_1 = n161_O_2_0_1; // @[Top.scala 180:12]
  assign n168_I_3_0_0 = n161_O_3_0_0; // @[Top.scala 180:12]
  assign n168_I_3_0_1 = n161_O_3_0_1; // @[Top.scala 180:12]
  assign n168_I_4_0_0 = n161_O_4_0_0; // @[Top.scala 180:12]
  assign n168_I_4_0_1 = n161_O_4_0_1; // @[Top.scala 180:12]
  assign n168_I_5_0_0 = n161_O_5_0_0; // @[Top.scala 180:12]
  assign n168_I_5_0_1 = n161_O_5_0_1; // @[Top.scala 180:12]
  assign n168_I_6_0_0 = n161_O_6_0_0; // @[Top.scala 180:12]
  assign n168_I_6_0_1 = n161_O_6_0_1; // @[Top.scala 180:12]
  assign n168_I_7_0_0 = n161_O_7_0_0; // @[Top.scala 180:12]
  assign n168_I_7_0_1 = n161_O_7_0_1; // @[Top.scala 180:12]
  assign n168_I_8_0_0 = n161_O_8_0_0; // @[Top.scala 180:12]
  assign n168_I_8_0_1 = n161_O_8_0_1; // @[Top.scala 180:12]
  assign n168_I_9_0_0 = n161_O_9_0_0; // @[Top.scala 180:12]
  assign n168_I_9_0_1 = n161_O_9_0_1; // @[Top.scala 180:12]
  assign n168_I_10_0_0 = n161_O_10_0_0; // @[Top.scala 180:12]
  assign n168_I_10_0_1 = n161_O_10_0_1; // @[Top.scala 180:12]
  assign n168_I_11_0_0 = n161_O_11_0_0; // @[Top.scala 180:12]
  assign n168_I_11_0_1 = n161_O_11_0_1; // @[Top.scala 180:12]
  assign n168_I_12_0_0 = n161_O_12_0_0; // @[Top.scala 180:12]
  assign n168_I_12_0_1 = n161_O_12_0_1; // @[Top.scala 180:12]
  assign n168_I_13_0_0 = n161_O_13_0_0; // @[Top.scala 180:12]
  assign n168_I_13_0_1 = n161_O_13_0_1; // @[Top.scala 180:12]
  assign n168_I_14_0_0 = n161_O_14_0_0; // @[Top.scala 180:12]
  assign n168_I_14_0_1 = n161_O_14_0_1; // @[Top.scala 180:12]
  assign n168_I_15_0_0 = n161_O_15_0_0; // @[Top.scala 180:12]
  assign n168_I_15_0_1 = n161_O_15_0_1; // @[Top.scala 180:12]
  assign n169_clock = clock;
  assign n169_valid_up = n149_valid_down; // @[Top.scala 184:19]
  assign n169_I_0 = n149_O_0; // @[Top.scala 183:12]
  assign n169_I_1 = n149_O_1; // @[Top.scala 183:12]
  assign n169_I_2 = n149_O_2; // @[Top.scala 183:12]
  assign n169_I_3 = n149_O_3; // @[Top.scala 183:12]
  assign n169_I_4 = n149_O_4; // @[Top.scala 183:12]
  assign n169_I_5 = n149_O_5; // @[Top.scala 183:12]
  assign n169_I_6 = n149_O_6; // @[Top.scala 183:12]
  assign n169_I_7 = n149_O_7; // @[Top.scala 183:12]
  assign n169_I_8 = n149_O_8; // @[Top.scala 183:12]
  assign n169_I_9 = n149_O_9; // @[Top.scala 183:12]
  assign n169_I_10 = n149_O_10; // @[Top.scala 183:12]
  assign n169_I_11 = n149_O_11; // @[Top.scala 183:12]
  assign n169_I_12 = n149_O_12; // @[Top.scala 183:12]
  assign n169_I_13 = n149_O_13; // @[Top.scala 183:12]
  assign n169_I_14 = n149_O_14; // @[Top.scala 183:12]
  assign n169_I_15 = n149_O_15; // @[Top.scala 183:12]
  assign n170_valid_up = n169_valid_down & n149_valid_down; // @[Top.scala 188:19]
  assign n170_I0_0 = n169_O_0; // @[Top.scala 186:13]
  assign n170_I0_1 = n169_O_1; // @[Top.scala 186:13]
  assign n170_I0_2 = n169_O_2; // @[Top.scala 186:13]
  assign n170_I0_3 = n169_O_3; // @[Top.scala 186:13]
  assign n170_I0_4 = n169_O_4; // @[Top.scala 186:13]
  assign n170_I0_5 = n169_O_5; // @[Top.scala 186:13]
  assign n170_I0_6 = n169_O_6; // @[Top.scala 186:13]
  assign n170_I0_7 = n169_O_7; // @[Top.scala 186:13]
  assign n170_I0_8 = n169_O_8; // @[Top.scala 186:13]
  assign n170_I0_9 = n169_O_9; // @[Top.scala 186:13]
  assign n170_I0_10 = n169_O_10; // @[Top.scala 186:13]
  assign n170_I0_11 = n169_O_11; // @[Top.scala 186:13]
  assign n170_I0_12 = n169_O_12; // @[Top.scala 186:13]
  assign n170_I0_13 = n169_O_13; // @[Top.scala 186:13]
  assign n170_I0_14 = n169_O_14; // @[Top.scala 186:13]
  assign n170_I0_15 = n169_O_15; // @[Top.scala 186:13]
  assign n170_I1_0 = n149_O_0; // @[Top.scala 187:13]
  assign n170_I1_1 = n149_O_1; // @[Top.scala 187:13]
  assign n170_I1_2 = n149_O_2; // @[Top.scala 187:13]
  assign n170_I1_3 = n149_O_3; // @[Top.scala 187:13]
  assign n170_I1_4 = n149_O_4; // @[Top.scala 187:13]
  assign n170_I1_5 = n149_O_5; // @[Top.scala 187:13]
  assign n170_I1_6 = n149_O_6; // @[Top.scala 187:13]
  assign n170_I1_7 = n149_O_7; // @[Top.scala 187:13]
  assign n170_I1_8 = n149_O_8; // @[Top.scala 187:13]
  assign n170_I1_9 = n149_O_9; // @[Top.scala 187:13]
  assign n170_I1_10 = n149_O_10; // @[Top.scala 187:13]
  assign n170_I1_11 = n149_O_11; // @[Top.scala 187:13]
  assign n170_I1_12 = n149_O_12; // @[Top.scala 187:13]
  assign n170_I1_13 = n149_O_13; // @[Top.scala 187:13]
  assign n170_I1_14 = n149_O_14; // @[Top.scala 187:13]
  assign n170_I1_15 = n149_O_15; // @[Top.scala 187:13]
  assign n179_valid_up = n170_valid_down; // @[Top.scala 191:19]
  assign n179_I_0_0 = n170_O_0_0; // @[Top.scala 190:12]
  assign n179_I_0_1 = n170_O_0_1; // @[Top.scala 190:12]
  assign n179_I_1_0 = n170_O_1_0; // @[Top.scala 190:12]
  assign n179_I_1_1 = n170_O_1_1; // @[Top.scala 190:12]
  assign n179_I_2_0 = n170_O_2_0; // @[Top.scala 190:12]
  assign n179_I_2_1 = n170_O_2_1; // @[Top.scala 190:12]
  assign n179_I_3_0 = n170_O_3_0; // @[Top.scala 190:12]
  assign n179_I_3_1 = n170_O_3_1; // @[Top.scala 190:12]
  assign n179_I_4_0 = n170_O_4_0; // @[Top.scala 190:12]
  assign n179_I_4_1 = n170_O_4_1; // @[Top.scala 190:12]
  assign n179_I_5_0 = n170_O_5_0; // @[Top.scala 190:12]
  assign n179_I_5_1 = n170_O_5_1; // @[Top.scala 190:12]
  assign n179_I_6_0 = n170_O_6_0; // @[Top.scala 190:12]
  assign n179_I_6_1 = n170_O_6_1; // @[Top.scala 190:12]
  assign n179_I_7_0 = n170_O_7_0; // @[Top.scala 190:12]
  assign n179_I_7_1 = n170_O_7_1; // @[Top.scala 190:12]
  assign n179_I_8_0 = n170_O_8_0; // @[Top.scala 190:12]
  assign n179_I_8_1 = n170_O_8_1; // @[Top.scala 190:12]
  assign n179_I_9_0 = n170_O_9_0; // @[Top.scala 190:12]
  assign n179_I_9_1 = n170_O_9_1; // @[Top.scala 190:12]
  assign n179_I_10_0 = n170_O_10_0; // @[Top.scala 190:12]
  assign n179_I_10_1 = n170_O_10_1; // @[Top.scala 190:12]
  assign n179_I_11_0 = n170_O_11_0; // @[Top.scala 190:12]
  assign n179_I_11_1 = n170_O_11_1; // @[Top.scala 190:12]
  assign n179_I_12_0 = n170_O_12_0; // @[Top.scala 190:12]
  assign n179_I_12_1 = n170_O_12_1; // @[Top.scala 190:12]
  assign n179_I_13_0 = n170_O_13_0; // @[Top.scala 190:12]
  assign n179_I_13_1 = n170_O_13_1; // @[Top.scala 190:12]
  assign n179_I_14_0 = n170_O_14_0; // @[Top.scala 190:12]
  assign n179_I_14_1 = n170_O_14_1; // @[Top.scala 190:12]
  assign n179_I_15_0 = n170_O_15_0; // @[Top.scala 190:12]
  assign n179_I_15_1 = n170_O_15_1; // @[Top.scala 190:12]
  assign n186_valid_up = n179_valid_down; // @[Top.scala 194:19]
  assign n186_I_0_0_0 = n179_O_0_0_0; // @[Top.scala 193:12]
  assign n186_I_0_0_1 = n179_O_0_0_1; // @[Top.scala 193:12]
  assign n186_I_1_0_0 = n179_O_1_0_0; // @[Top.scala 193:12]
  assign n186_I_1_0_1 = n179_O_1_0_1; // @[Top.scala 193:12]
  assign n186_I_2_0_0 = n179_O_2_0_0; // @[Top.scala 193:12]
  assign n186_I_2_0_1 = n179_O_2_0_1; // @[Top.scala 193:12]
  assign n186_I_3_0_0 = n179_O_3_0_0; // @[Top.scala 193:12]
  assign n186_I_3_0_1 = n179_O_3_0_1; // @[Top.scala 193:12]
  assign n186_I_4_0_0 = n179_O_4_0_0; // @[Top.scala 193:12]
  assign n186_I_4_0_1 = n179_O_4_0_1; // @[Top.scala 193:12]
  assign n186_I_5_0_0 = n179_O_5_0_0; // @[Top.scala 193:12]
  assign n186_I_5_0_1 = n179_O_5_0_1; // @[Top.scala 193:12]
  assign n186_I_6_0_0 = n179_O_6_0_0; // @[Top.scala 193:12]
  assign n186_I_6_0_1 = n179_O_6_0_1; // @[Top.scala 193:12]
  assign n186_I_7_0_0 = n179_O_7_0_0; // @[Top.scala 193:12]
  assign n186_I_7_0_1 = n179_O_7_0_1; // @[Top.scala 193:12]
  assign n186_I_8_0_0 = n179_O_8_0_0; // @[Top.scala 193:12]
  assign n186_I_8_0_1 = n179_O_8_0_1; // @[Top.scala 193:12]
  assign n186_I_9_0_0 = n179_O_9_0_0; // @[Top.scala 193:12]
  assign n186_I_9_0_1 = n179_O_9_0_1; // @[Top.scala 193:12]
  assign n186_I_10_0_0 = n179_O_10_0_0; // @[Top.scala 193:12]
  assign n186_I_10_0_1 = n179_O_10_0_1; // @[Top.scala 193:12]
  assign n186_I_11_0_0 = n179_O_11_0_0; // @[Top.scala 193:12]
  assign n186_I_11_0_1 = n179_O_11_0_1; // @[Top.scala 193:12]
  assign n186_I_12_0_0 = n179_O_12_0_0; // @[Top.scala 193:12]
  assign n186_I_12_0_1 = n179_O_12_0_1; // @[Top.scala 193:12]
  assign n186_I_13_0_0 = n179_O_13_0_0; // @[Top.scala 193:12]
  assign n186_I_13_0_1 = n179_O_13_0_1; // @[Top.scala 193:12]
  assign n186_I_14_0_0 = n179_O_14_0_0; // @[Top.scala 193:12]
  assign n186_I_14_0_1 = n179_O_14_0_1; // @[Top.scala 193:12]
  assign n186_I_15_0_0 = n179_O_15_0_0; // @[Top.scala 193:12]
  assign n186_I_15_0_1 = n179_O_15_0_1; // @[Top.scala 193:12]
  assign n187_valid_up = n168_valid_down & n186_valid_down; // @[Top.scala 198:19]
  assign n187_I0_0_0 = n168_O_0_0; // @[Top.scala 196:13]
  assign n187_I0_0_1 = n168_O_0_1; // @[Top.scala 196:13]
  assign n187_I0_1_0 = n168_O_1_0; // @[Top.scala 196:13]
  assign n187_I0_1_1 = n168_O_1_1; // @[Top.scala 196:13]
  assign n187_I0_2_0 = n168_O_2_0; // @[Top.scala 196:13]
  assign n187_I0_2_1 = n168_O_2_1; // @[Top.scala 196:13]
  assign n187_I0_3_0 = n168_O_3_0; // @[Top.scala 196:13]
  assign n187_I0_3_1 = n168_O_3_1; // @[Top.scala 196:13]
  assign n187_I0_4_0 = n168_O_4_0; // @[Top.scala 196:13]
  assign n187_I0_4_1 = n168_O_4_1; // @[Top.scala 196:13]
  assign n187_I0_5_0 = n168_O_5_0; // @[Top.scala 196:13]
  assign n187_I0_5_1 = n168_O_5_1; // @[Top.scala 196:13]
  assign n187_I0_6_0 = n168_O_6_0; // @[Top.scala 196:13]
  assign n187_I0_6_1 = n168_O_6_1; // @[Top.scala 196:13]
  assign n187_I0_7_0 = n168_O_7_0; // @[Top.scala 196:13]
  assign n187_I0_7_1 = n168_O_7_1; // @[Top.scala 196:13]
  assign n187_I0_8_0 = n168_O_8_0; // @[Top.scala 196:13]
  assign n187_I0_8_1 = n168_O_8_1; // @[Top.scala 196:13]
  assign n187_I0_9_0 = n168_O_9_0; // @[Top.scala 196:13]
  assign n187_I0_9_1 = n168_O_9_1; // @[Top.scala 196:13]
  assign n187_I0_10_0 = n168_O_10_0; // @[Top.scala 196:13]
  assign n187_I0_10_1 = n168_O_10_1; // @[Top.scala 196:13]
  assign n187_I0_11_0 = n168_O_11_0; // @[Top.scala 196:13]
  assign n187_I0_11_1 = n168_O_11_1; // @[Top.scala 196:13]
  assign n187_I0_12_0 = n168_O_12_0; // @[Top.scala 196:13]
  assign n187_I0_12_1 = n168_O_12_1; // @[Top.scala 196:13]
  assign n187_I0_13_0 = n168_O_13_0; // @[Top.scala 196:13]
  assign n187_I0_13_1 = n168_O_13_1; // @[Top.scala 196:13]
  assign n187_I0_14_0 = n168_O_14_0; // @[Top.scala 196:13]
  assign n187_I0_14_1 = n168_O_14_1; // @[Top.scala 196:13]
  assign n187_I0_15_0 = n168_O_15_0; // @[Top.scala 196:13]
  assign n187_I0_15_1 = n168_O_15_1; // @[Top.scala 196:13]
  assign n187_I1_0_0 = n186_O_0_0; // @[Top.scala 197:13]
  assign n187_I1_0_1 = n186_O_0_1; // @[Top.scala 197:13]
  assign n187_I1_1_0 = n186_O_1_0; // @[Top.scala 197:13]
  assign n187_I1_1_1 = n186_O_1_1; // @[Top.scala 197:13]
  assign n187_I1_2_0 = n186_O_2_0; // @[Top.scala 197:13]
  assign n187_I1_2_1 = n186_O_2_1; // @[Top.scala 197:13]
  assign n187_I1_3_0 = n186_O_3_0; // @[Top.scala 197:13]
  assign n187_I1_3_1 = n186_O_3_1; // @[Top.scala 197:13]
  assign n187_I1_4_0 = n186_O_4_0; // @[Top.scala 197:13]
  assign n187_I1_4_1 = n186_O_4_1; // @[Top.scala 197:13]
  assign n187_I1_5_0 = n186_O_5_0; // @[Top.scala 197:13]
  assign n187_I1_5_1 = n186_O_5_1; // @[Top.scala 197:13]
  assign n187_I1_6_0 = n186_O_6_0; // @[Top.scala 197:13]
  assign n187_I1_6_1 = n186_O_6_1; // @[Top.scala 197:13]
  assign n187_I1_7_0 = n186_O_7_0; // @[Top.scala 197:13]
  assign n187_I1_7_1 = n186_O_7_1; // @[Top.scala 197:13]
  assign n187_I1_8_0 = n186_O_8_0; // @[Top.scala 197:13]
  assign n187_I1_8_1 = n186_O_8_1; // @[Top.scala 197:13]
  assign n187_I1_9_0 = n186_O_9_0; // @[Top.scala 197:13]
  assign n187_I1_9_1 = n186_O_9_1; // @[Top.scala 197:13]
  assign n187_I1_10_0 = n186_O_10_0; // @[Top.scala 197:13]
  assign n187_I1_10_1 = n186_O_10_1; // @[Top.scala 197:13]
  assign n187_I1_11_0 = n186_O_11_0; // @[Top.scala 197:13]
  assign n187_I1_11_1 = n186_O_11_1; // @[Top.scala 197:13]
  assign n187_I1_12_0 = n186_O_12_0; // @[Top.scala 197:13]
  assign n187_I1_12_1 = n186_O_12_1; // @[Top.scala 197:13]
  assign n187_I1_13_0 = n186_O_13_0; // @[Top.scala 197:13]
  assign n187_I1_13_1 = n186_O_13_1; // @[Top.scala 197:13]
  assign n187_I1_14_0 = n186_O_14_0; // @[Top.scala 197:13]
  assign n187_I1_14_1 = n186_O_14_1; // @[Top.scala 197:13]
  assign n187_I1_15_0 = n186_O_15_0; // @[Top.scala 197:13]
  assign n187_I1_15_1 = n186_O_15_1; // @[Top.scala 197:13]
  assign n196_valid_up = n187_valid_down; // @[Top.scala 201:19]
  assign n196_I_0_0_0 = n187_O_0_0_0; // @[Top.scala 200:12]
  assign n196_I_0_0_1 = n187_O_0_0_1; // @[Top.scala 200:12]
  assign n196_I_0_1_0 = n187_O_0_1_0; // @[Top.scala 200:12]
  assign n196_I_0_1_1 = n187_O_0_1_1; // @[Top.scala 200:12]
  assign n196_I_1_0_0 = n187_O_1_0_0; // @[Top.scala 200:12]
  assign n196_I_1_0_1 = n187_O_1_0_1; // @[Top.scala 200:12]
  assign n196_I_1_1_0 = n187_O_1_1_0; // @[Top.scala 200:12]
  assign n196_I_1_1_1 = n187_O_1_1_1; // @[Top.scala 200:12]
  assign n196_I_2_0_0 = n187_O_2_0_0; // @[Top.scala 200:12]
  assign n196_I_2_0_1 = n187_O_2_0_1; // @[Top.scala 200:12]
  assign n196_I_2_1_0 = n187_O_2_1_0; // @[Top.scala 200:12]
  assign n196_I_2_1_1 = n187_O_2_1_1; // @[Top.scala 200:12]
  assign n196_I_3_0_0 = n187_O_3_0_0; // @[Top.scala 200:12]
  assign n196_I_3_0_1 = n187_O_3_0_1; // @[Top.scala 200:12]
  assign n196_I_3_1_0 = n187_O_3_1_0; // @[Top.scala 200:12]
  assign n196_I_3_1_1 = n187_O_3_1_1; // @[Top.scala 200:12]
  assign n196_I_4_0_0 = n187_O_4_0_0; // @[Top.scala 200:12]
  assign n196_I_4_0_1 = n187_O_4_0_1; // @[Top.scala 200:12]
  assign n196_I_4_1_0 = n187_O_4_1_0; // @[Top.scala 200:12]
  assign n196_I_4_1_1 = n187_O_4_1_1; // @[Top.scala 200:12]
  assign n196_I_5_0_0 = n187_O_5_0_0; // @[Top.scala 200:12]
  assign n196_I_5_0_1 = n187_O_5_0_1; // @[Top.scala 200:12]
  assign n196_I_5_1_0 = n187_O_5_1_0; // @[Top.scala 200:12]
  assign n196_I_5_1_1 = n187_O_5_1_1; // @[Top.scala 200:12]
  assign n196_I_6_0_0 = n187_O_6_0_0; // @[Top.scala 200:12]
  assign n196_I_6_0_1 = n187_O_6_0_1; // @[Top.scala 200:12]
  assign n196_I_6_1_0 = n187_O_6_1_0; // @[Top.scala 200:12]
  assign n196_I_6_1_1 = n187_O_6_1_1; // @[Top.scala 200:12]
  assign n196_I_7_0_0 = n187_O_7_0_0; // @[Top.scala 200:12]
  assign n196_I_7_0_1 = n187_O_7_0_1; // @[Top.scala 200:12]
  assign n196_I_7_1_0 = n187_O_7_1_0; // @[Top.scala 200:12]
  assign n196_I_7_1_1 = n187_O_7_1_1; // @[Top.scala 200:12]
  assign n196_I_8_0_0 = n187_O_8_0_0; // @[Top.scala 200:12]
  assign n196_I_8_0_1 = n187_O_8_0_1; // @[Top.scala 200:12]
  assign n196_I_8_1_0 = n187_O_8_1_0; // @[Top.scala 200:12]
  assign n196_I_8_1_1 = n187_O_8_1_1; // @[Top.scala 200:12]
  assign n196_I_9_0_0 = n187_O_9_0_0; // @[Top.scala 200:12]
  assign n196_I_9_0_1 = n187_O_9_0_1; // @[Top.scala 200:12]
  assign n196_I_9_1_0 = n187_O_9_1_0; // @[Top.scala 200:12]
  assign n196_I_9_1_1 = n187_O_9_1_1; // @[Top.scala 200:12]
  assign n196_I_10_0_0 = n187_O_10_0_0; // @[Top.scala 200:12]
  assign n196_I_10_0_1 = n187_O_10_0_1; // @[Top.scala 200:12]
  assign n196_I_10_1_0 = n187_O_10_1_0; // @[Top.scala 200:12]
  assign n196_I_10_1_1 = n187_O_10_1_1; // @[Top.scala 200:12]
  assign n196_I_11_0_0 = n187_O_11_0_0; // @[Top.scala 200:12]
  assign n196_I_11_0_1 = n187_O_11_0_1; // @[Top.scala 200:12]
  assign n196_I_11_1_0 = n187_O_11_1_0; // @[Top.scala 200:12]
  assign n196_I_11_1_1 = n187_O_11_1_1; // @[Top.scala 200:12]
  assign n196_I_12_0_0 = n187_O_12_0_0; // @[Top.scala 200:12]
  assign n196_I_12_0_1 = n187_O_12_0_1; // @[Top.scala 200:12]
  assign n196_I_12_1_0 = n187_O_12_1_0; // @[Top.scala 200:12]
  assign n196_I_12_1_1 = n187_O_12_1_1; // @[Top.scala 200:12]
  assign n196_I_13_0_0 = n187_O_13_0_0; // @[Top.scala 200:12]
  assign n196_I_13_0_1 = n187_O_13_0_1; // @[Top.scala 200:12]
  assign n196_I_13_1_0 = n187_O_13_1_0; // @[Top.scala 200:12]
  assign n196_I_13_1_1 = n187_O_13_1_1; // @[Top.scala 200:12]
  assign n196_I_14_0_0 = n187_O_14_0_0; // @[Top.scala 200:12]
  assign n196_I_14_0_1 = n187_O_14_0_1; // @[Top.scala 200:12]
  assign n196_I_14_1_0 = n187_O_14_1_0; // @[Top.scala 200:12]
  assign n196_I_14_1_1 = n187_O_14_1_1; // @[Top.scala 200:12]
  assign n196_I_15_0_0 = n187_O_15_0_0; // @[Top.scala 200:12]
  assign n196_I_15_0_1 = n187_O_15_0_1; // @[Top.scala 200:12]
  assign n196_I_15_1_0 = n187_O_15_1_0; // @[Top.scala 200:12]
  assign n196_I_15_1_1 = n187_O_15_1_1; // @[Top.scala 200:12]
  assign n203_valid_up = n196_valid_down; // @[Top.scala 204:19]
  assign n203_I_0_0_0_0 = n196_O_0_0_0_0; // @[Top.scala 203:12]
  assign n203_I_0_0_0_1 = n196_O_0_0_0_1; // @[Top.scala 203:12]
  assign n203_I_0_0_1_0 = n196_O_0_0_1_0; // @[Top.scala 203:12]
  assign n203_I_0_0_1_1 = n196_O_0_0_1_1; // @[Top.scala 203:12]
  assign n203_I_1_0_0_0 = n196_O_1_0_0_0; // @[Top.scala 203:12]
  assign n203_I_1_0_0_1 = n196_O_1_0_0_1; // @[Top.scala 203:12]
  assign n203_I_1_0_1_0 = n196_O_1_0_1_0; // @[Top.scala 203:12]
  assign n203_I_1_0_1_1 = n196_O_1_0_1_1; // @[Top.scala 203:12]
  assign n203_I_2_0_0_0 = n196_O_2_0_0_0; // @[Top.scala 203:12]
  assign n203_I_2_0_0_1 = n196_O_2_0_0_1; // @[Top.scala 203:12]
  assign n203_I_2_0_1_0 = n196_O_2_0_1_0; // @[Top.scala 203:12]
  assign n203_I_2_0_1_1 = n196_O_2_0_1_1; // @[Top.scala 203:12]
  assign n203_I_3_0_0_0 = n196_O_3_0_0_0; // @[Top.scala 203:12]
  assign n203_I_3_0_0_1 = n196_O_3_0_0_1; // @[Top.scala 203:12]
  assign n203_I_3_0_1_0 = n196_O_3_0_1_0; // @[Top.scala 203:12]
  assign n203_I_3_0_1_1 = n196_O_3_0_1_1; // @[Top.scala 203:12]
  assign n203_I_4_0_0_0 = n196_O_4_0_0_0; // @[Top.scala 203:12]
  assign n203_I_4_0_0_1 = n196_O_4_0_0_1; // @[Top.scala 203:12]
  assign n203_I_4_0_1_0 = n196_O_4_0_1_0; // @[Top.scala 203:12]
  assign n203_I_4_0_1_1 = n196_O_4_0_1_1; // @[Top.scala 203:12]
  assign n203_I_5_0_0_0 = n196_O_5_0_0_0; // @[Top.scala 203:12]
  assign n203_I_5_0_0_1 = n196_O_5_0_0_1; // @[Top.scala 203:12]
  assign n203_I_5_0_1_0 = n196_O_5_0_1_0; // @[Top.scala 203:12]
  assign n203_I_5_0_1_1 = n196_O_5_0_1_1; // @[Top.scala 203:12]
  assign n203_I_6_0_0_0 = n196_O_6_0_0_0; // @[Top.scala 203:12]
  assign n203_I_6_0_0_1 = n196_O_6_0_0_1; // @[Top.scala 203:12]
  assign n203_I_6_0_1_0 = n196_O_6_0_1_0; // @[Top.scala 203:12]
  assign n203_I_6_0_1_1 = n196_O_6_0_1_1; // @[Top.scala 203:12]
  assign n203_I_7_0_0_0 = n196_O_7_0_0_0; // @[Top.scala 203:12]
  assign n203_I_7_0_0_1 = n196_O_7_0_0_1; // @[Top.scala 203:12]
  assign n203_I_7_0_1_0 = n196_O_7_0_1_0; // @[Top.scala 203:12]
  assign n203_I_7_0_1_1 = n196_O_7_0_1_1; // @[Top.scala 203:12]
  assign n203_I_8_0_0_0 = n196_O_8_0_0_0; // @[Top.scala 203:12]
  assign n203_I_8_0_0_1 = n196_O_8_0_0_1; // @[Top.scala 203:12]
  assign n203_I_8_0_1_0 = n196_O_8_0_1_0; // @[Top.scala 203:12]
  assign n203_I_8_0_1_1 = n196_O_8_0_1_1; // @[Top.scala 203:12]
  assign n203_I_9_0_0_0 = n196_O_9_0_0_0; // @[Top.scala 203:12]
  assign n203_I_9_0_0_1 = n196_O_9_0_0_1; // @[Top.scala 203:12]
  assign n203_I_9_0_1_0 = n196_O_9_0_1_0; // @[Top.scala 203:12]
  assign n203_I_9_0_1_1 = n196_O_9_0_1_1; // @[Top.scala 203:12]
  assign n203_I_10_0_0_0 = n196_O_10_0_0_0; // @[Top.scala 203:12]
  assign n203_I_10_0_0_1 = n196_O_10_0_0_1; // @[Top.scala 203:12]
  assign n203_I_10_0_1_0 = n196_O_10_0_1_0; // @[Top.scala 203:12]
  assign n203_I_10_0_1_1 = n196_O_10_0_1_1; // @[Top.scala 203:12]
  assign n203_I_11_0_0_0 = n196_O_11_0_0_0; // @[Top.scala 203:12]
  assign n203_I_11_0_0_1 = n196_O_11_0_0_1; // @[Top.scala 203:12]
  assign n203_I_11_0_1_0 = n196_O_11_0_1_0; // @[Top.scala 203:12]
  assign n203_I_11_0_1_1 = n196_O_11_0_1_1; // @[Top.scala 203:12]
  assign n203_I_12_0_0_0 = n196_O_12_0_0_0; // @[Top.scala 203:12]
  assign n203_I_12_0_0_1 = n196_O_12_0_0_1; // @[Top.scala 203:12]
  assign n203_I_12_0_1_0 = n196_O_12_0_1_0; // @[Top.scala 203:12]
  assign n203_I_12_0_1_1 = n196_O_12_0_1_1; // @[Top.scala 203:12]
  assign n203_I_13_0_0_0 = n196_O_13_0_0_0; // @[Top.scala 203:12]
  assign n203_I_13_0_0_1 = n196_O_13_0_0_1; // @[Top.scala 203:12]
  assign n203_I_13_0_1_0 = n196_O_13_0_1_0; // @[Top.scala 203:12]
  assign n203_I_13_0_1_1 = n196_O_13_0_1_1; // @[Top.scala 203:12]
  assign n203_I_14_0_0_0 = n196_O_14_0_0_0; // @[Top.scala 203:12]
  assign n203_I_14_0_0_1 = n196_O_14_0_0_1; // @[Top.scala 203:12]
  assign n203_I_14_0_1_0 = n196_O_14_0_1_0; // @[Top.scala 203:12]
  assign n203_I_14_0_1_1 = n196_O_14_0_1_1; // @[Top.scala 203:12]
  assign n203_I_15_0_0_0 = n196_O_15_0_0_0; // @[Top.scala 203:12]
  assign n203_I_15_0_0_1 = n196_O_15_0_0_1; // @[Top.scala 203:12]
  assign n203_I_15_0_1_0 = n196_O_15_0_1_0; // @[Top.scala 203:12]
  assign n203_I_15_0_1_1 = n196_O_15_0_1_1; // @[Top.scala 203:12]
  assign n245_clock = clock;
  assign n245_reset = reset;
  assign n245_valid_up = n203_valid_down; // @[Top.scala 207:19]
  assign n245_I_0_0_0 = n203_O_0_0_0; // @[Top.scala 206:12]
  assign n245_I_0_0_1 = n203_O_0_0_1; // @[Top.scala 206:12]
  assign n245_I_0_1_0 = n203_O_0_1_0; // @[Top.scala 206:12]
  assign n245_I_0_1_1 = n203_O_0_1_1; // @[Top.scala 206:12]
  assign n245_I_1_0_0 = n203_O_1_0_0; // @[Top.scala 206:12]
  assign n245_I_1_0_1 = n203_O_1_0_1; // @[Top.scala 206:12]
  assign n245_I_1_1_0 = n203_O_1_1_0; // @[Top.scala 206:12]
  assign n245_I_1_1_1 = n203_O_1_1_1; // @[Top.scala 206:12]
  assign n245_I_2_0_0 = n203_O_2_0_0; // @[Top.scala 206:12]
  assign n245_I_2_0_1 = n203_O_2_0_1; // @[Top.scala 206:12]
  assign n245_I_2_1_0 = n203_O_2_1_0; // @[Top.scala 206:12]
  assign n245_I_2_1_1 = n203_O_2_1_1; // @[Top.scala 206:12]
  assign n245_I_3_0_0 = n203_O_3_0_0; // @[Top.scala 206:12]
  assign n245_I_3_0_1 = n203_O_3_0_1; // @[Top.scala 206:12]
  assign n245_I_3_1_0 = n203_O_3_1_0; // @[Top.scala 206:12]
  assign n245_I_3_1_1 = n203_O_3_1_1; // @[Top.scala 206:12]
  assign n245_I_4_0_0 = n203_O_4_0_0; // @[Top.scala 206:12]
  assign n245_I_4_0_1 = n203_O_4_0_1; // @[Top.scala 206:12]
  assign n245_I_4_1_0 = n203_O_4_1_0; // @[Top.scala 206:12]
  assign n245_I_4_1_1 = n203_O_4_1_1; // @[Top.scala 206:12]
  assign n245_I_5_0_0 = n203_O_5_0_0; // @[Top.scala 206:12]
  assign n245_I_5_0_1 = n203_O_5_0_1; // @[Top.scala 206:12]
  assign n245_I_5_1_0 = n203_O_5_1_0; // @[Top.scala 206:12]
  assign n245_I_5_1_1 = n203_O_5_1_1; // @[Top.scala 206:12]
  assign n245_I_6_0_0 = n203_O_6_0_0; // @[Top.scala 206:12]
  assign n245_I_6_0_1 = n203_O_6_0_1; // @[Top.scala 206:12]
  assign n245_I_6_1_0 = n203_O_6_1_0; // @[Top.scala 206:12]
  assign n245_I_6_1_1 = n203_O_6_1_1; // @[Top.scala 206:12]
  assign n245_I_7_0_0 = n203_O_7_0_0; // @[Top.scala 206:12]
  assign n245_I_7_0_1 = n203_O_7_0_1; // @[Top.scala 206:12]
  assign n245_I_7_1_0 = n203_O_7_1_0; // @[Top.scala 206:12]
  assign n245_I_7_1_1 = n203_O_7_1_1; // @[Top.scala 206:12]
  assign n245_I_8_0_0 = n203_O_8_0_0; // @[Top.scala 206:12]
  assign n245_I_8_0_1 = n203_O_8_0_1; // @[Top.scala 206:12]
  assign n245_I_8_1_0 = n203_O_8_1_0; // @[Top.scala 206:12]
  assign n245_I_8_1_1 = n203_O_8_1_1; // @[Top.scala 206:12]
  assign n245_I_9_0_0 = n203_O_9_0_0; // @[Top.scala 206:12]
  assign n245_I_9_0_1 = n203_O_9_0_1; // @[Top.scala 206:12]
  assign n245_I_9_1_0 = n203_O_9_1_0; // @[Top.scala 206:12]
  assign n245_I_9_1_1 = n203_O_9_1_1; // @[Top.scala 206:12]
  assign n245_I_10_0_0 = n203_O_10_0_0; // @[Top.scala 206:12]
  assign n245_I_10_0_1 = n203_O_10_0_1; // @[Top.scala 206:12]
  assign n245_I_10_1_0 = n203_O_10_1_0; // @[Top.scala 206:12]
  assign n245_I_10_1_1 = n203_O_10_1_1; // @[Top.scala 206:12]
  assign n245_I_11_0_0 = n203_O_11_0_0; // @[Top.scala 206:12]
  assign n245_I_11_0_1 = n203_O_11_0_1; // @[Top.scala 206:12]
  assign n245_I_11_1_0 = n203_O_11_1_0; // @[Top.scala 206:12]
  assign n245_I_11_1_1 = n203_O_11_1_1; // @[Top.scala 206:12]
  assign n245_I_12_0_0 = n203_O_12_0_0; // @[Top.scala 206:12]
  assign n245_I_12_0_1 = n203_O_12_0_1; // @[Top.scala 206:12]
  assign n245_I_12_1_0 = n203_O_12_1_0; // @[Top.scala 206:12]
  assign n245_I_12_1_1 = n203_O_12_1_1; // @[Top.scala 206:12]
  assign n245_I_13_0_0 = n203_O_13_0_0; // @[Top.scala 206:12]
  assign n245_I_13_0_1 = n203_O_13_0_1; // @[Top.scala 206:12]
  assign n245_I_13_1_0 = n203_O_13_1_0; // @[Top.scala 206:12]
  assign n245_I_13_1_1 = n203_O_13_1_1; // @[Top.scala 206:12]
  assign n245_I_14_0_0 = n203_O_14_0_0; // @[Top.scala 206:12]
  assign n245_I_14_0_1 = n203_O_14_0_1; // @[Top.scala 206:12]
  assign n245_I_14_1_0 = n203_O_14_1_0; // @[Top.scala 206:12]
  assign n245_I_14_1_1 = n203_O_14_1_1; // @[Top.scala 206:12]
  assign n245_I_15_0_0 = n203_O_15_0_0; // @[Top.scala 206:12]
  assign n245_I_15_0_1 = n203_O_15_0_1; // @[Top.scala 206:12]
  assign n245_I_15_1_0 = n203_O_15_1_0; // @[Top.scala 206:12]
  assign n245_I_15_1_1 = n203_O_15_1_1; // @[Top.scala 206:12]
  assign n246_valid_up = n245_valid_down; // @[Top.scala 210:19]
  assign n246_I_0_0_0 = n245_O_0_0_0; // @[Top.scala 209:12]
  assign n246_I_1_0_0 = n245_O_1_0_0; // @[Top.scala 209:12]
  assign n246_I_2_0_0 = n245_O_2_0_0; // @[Top.scala 209:12]
  assign n246_I_3_0_0 = n245_O_3_0_0; // @[Top.scala 209:12]
  assign n246_I_4_0_0 = n245_O_4_0_0; // @[Top.scala 209:12]
  assign n246_I_5_0_0 = n245_O_5_0_0; // @[Top.scala 209:12]
  assign n246_I_6_0_0 = n245_O_6_0_0; // @[Top.scala 209:12]
  assign n246_I_7_0_0 = n245_O_7_0_0; // @[Top.scala 209:12]
  assign n246_I_8_0_0 = n245_O_8_0_0; // @[Top.scala 209:12]
  assign n246_I_9_0_0 = n245_O_9_0_0; // @[Top.scala 209:12]
  assign n246_I_10_0_0 = n245_O_10_0_0; // @[Top.scala 209:12]
  assign n246_I_11_0_0 = n245_O_11_0_0; // @[Top.scala 209:12]
  assign n246_I_12_0_0 = n245_O_12_0_0; // @[Top.scala 209:12]
  assign n246_I_13_0_0 = n245_O_13_0_0; // @[Top.scala 209:12]
  assign n246_I_14_0_0 = n245_O_14_0_0; // @[Top.scala 209:12]
  assign n246_I_15_0_0 = n245_O_15_0_0; // @[Top.scala 209:12]
  assign n247_valid_up = n246_valid_down; // @[Top.scala 213:19]
  assign n247_I_0_0 = n246_O_0_0; // @[Top.scala 212:12]
  assign n247_I_1_0 = n246_O_1_0; // @[Top.scala 212:12]
  assign n247_I_2_0 = n246_O_2_0; // @[Top.scala 212:12]
  assign n247_I_3_0 = n246_O_3_0; // @[Top.scala 212:12]
  assign n247_I_4_0 = n246_O_4_0; // @[Top.scala 212:12]
  assign n247_I_5_0 = n246_O_5_0; // @[Top.scala 212:12]
  assign n247_I_6_0 = n246_O_6_0; // @[Top.scala 212:12]
  assign n247_I_7_0 = n246_O_7_0; // @[Top.scala 212:12]
  assign n247_I_8_0 = n246_O_8_0; // @[Top.scala 212:12]
  assign n247_I_9_0 = n246_O_9_0; // @[Top.scala 212:12]
  assign n247_I_10_0 = n246_O_10_0; // @[Top.scala 212:12]
  assign n247_I_11_0 = n246_O_11_0; // @[Top.scala 212:12]
  assign n247_I_12_0 = n246_O_12_0; // @[Top.scala 212:12]
  assign n247_I_13_0 = n246_O_13_0; // @[Top.scala 212:12]
  assign n247_I_14_0 = n246_O_14_0; // @[Top.scala 212:12]
  assign n247_I_15_0 = n246_O_15_0; // @[Top.scala 212:12]
  assign n248_clock = clock;
  assign n248_reset = reset;
  assign n248_valid_up = n247_valid_down; // @[Top.scala 216:19]
  assign n248_I_0 = n247_O_0; // @[Top.scala 215:12]
  assign n248_I_1 = n247_O_1; // @[Top.scala 215:12]
  assign n248_I_2 = n247_O_2; // @[Top.scala 215:12]
  assign n248_I_3 = n247_O_3; // @[Top.scala 215:12]
  assign n248_I_4 = n247_O_4; // @[Top.scala 215:12]
  assign n248_I_5 = n247_O_5; // @[Top.scala 215:12]
  assign n248_I_6 = n247_O_6; // @[Top.scala 215:12]
  assign n248_I_7 = n247_O_7; // @[Top.scala 215:12]
  assign n248_I_8 = n247_O_8; // @[Top.scala 215:12]
  assign n248_I_9 = n247_O_9; // @[Top.scala 215:12]
  assign n248_I_10 = n247_O_10; // @[Top.scala 215:12]
  assign n248_I_11 = n247_O_11; // @[Top.scala 215:12]
  assign n248_I_12 = n247_O_12; // @[Top.scala 215:12]
  assign n248_I_13 = n247_O_13; // @[Top.scala 215:12]
  assign n248_I_14 = n247_O_14; // @[Top.scala 215:12]
  assign n248_I_15 = n247_O_15; // @[Top.scala 215:12]
  assign n249_clock = clock;
  assign n249_reset = reset;
  assign n249_valid_up = n248_valid_down; // @[Top.scala 219:19]
  assign n249_I_0 = n248_O_0; // @[Top.scala 218:12]
  assign n249_I_1 = n248_O_1; // @[Top.scala 218:12]
  assign n249_I_2 = n248_O_2; // @[Top.scala 218:12]
  assign n249_I_3 = n248_O_3; // @[Top.scala 218:12]
  assign n249_I_4 = n248_O_4; // @[Top.scala 218:12]
  assign n249_I_5 = n248_O_5; // @[Top.scala 218:12]
  assign n249_I_6 = n248_O_6; // @[Top.scala 218:12]
  assign n249_I_7 = n248_O_7; // @[Top.scala 218:12]
  assign n249_I_8 = n248_O_8; // @[Top.scala 218:12]
  assign n249_I_9 = n248_O_9; // @[Top.scala 218:12]
  assign n249_I_10 = n248_O_10; // @[Top.scala 218:12]
  assign n249_I_11 = n248_O_11; // @[Top.scala 218:12]
  assign n249_I_12 = n248_O_12; // @[Top.scala 218:12]
  assign n249_I_13 = n248_O_13; // @[Top.scala 218:12]
  assign n249_I_14 = n248_O_14; // @[Top.scala 218:12]
  assign n249_I_15 = n248_O_15; // @[Top.scala 218:12]
  assign n250_clock = clock;
  assign n250_reset = reset;
  assign n250_valid_up = n249_valid_down; // @[Top.scala 222:19]
  assign n250_I_0 = n249_O_0; // @[Top.scala 221:12]
  assign n250_I_1 = n249_O_1; // @[Top.scala 221:12]
  assign n250_I_2 = n249_O_2; // @[Top.scala 221:12]
  assign n250_I_3 = n249_O_3; // @[Top.scala 221:12]
  assign n250_I_4 = n249_O_4; // @[Top.scala 221:12]
  assign n250_I_5 = n249_O_5; // @[Top.scala 221:12]
  assign n250_I_6 = n249_O_6; // @[Top.scala 221:12]
  assign n250_I_7 = n249_O_7; // @[Top.scala 221:12]
  assign n250_I_8 = n249_O_8; // @[Top.scala 221:12]
  assign n250_I_9 = n249_O_9; // @[Top.scala 221:12]
  assign n250_I_10 = n249_O_10; // @[Top.scala 221:12]
  assign n250_I_11 = n249_O_11; // @[Top.scala 221:12]
  assign n250_I_12 = n249_O_12; // @[Top.scala 221:12]
  assign n250_I_13 = n249_O_13; // @[Top.scala 221:12]
  assign n250_I_14 = n249_O_14; // @[Top.scala 221:12]
  assign n250_I_15 = n249_O_15; // @[Top.scala 221:12]
endmodule
