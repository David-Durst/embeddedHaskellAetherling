// Latency = 4
module Top(
  input        clock,
  input        reset,
  input        valid_up,
  output       valid_down,
  input  [31:0] I_0,
  input  [31:0] I_1,
  output [31:0] O_0,
  output [31:0] O_1
);
  wire dontcare;
  wire [31:0] io_output_counts_1;
  wire [31:0] io_output_counts_0;

  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1 sampler_box ( // @[m_x55_ctr_0.scala 26:17:@1721.4]
    .clock(clock), // @[:@1296.4]
    .reset(reset), // @[:@1297.4]
    .io_in_x221_TREADY(dontcare), // @[:@1298.4]
    .io_in_x221_TDATA({I_0,I_1}), // @[:@1298.4]
    .io_in_x221_TID(8'h0),
    .io_in_x221_TDEST(8'h0),
    .io_in_x222_TVALID(valid_down), // @[:@1298.4]
    .io_in_x222_TDATA({O_0,O_1}), // @[:@1298.4]
    .io_in_x222_TREADY(1'b1), // @[:@1298.4]
    .io_sigsIn_datapathEn(valid_up), // @[:@1298.4]
    .io_sigsIn_backpressure(1'b1), // @[:@20563.4]
    .io_sigsIn_break(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_1(io_output_counts_1), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_counts_0(io_output_counts_0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_0(1'b0), // @[:@20563.4]
    .io_sigsIn_cchainOutputs_0_oobs_1(1'b0), // @[:@20563.4]
    .io_rr('b1) // @[:@1298.4]
  );

  wire dontcare2;

  wire io_output_oobs_0;
  wire io_output_oobs_1;
  x229_ctrchain cchain ( // @[:@2879.2]
    .clock(clock), // @[:@2880.4]
    .reset(reset), // @[:@2881.4]
    .io_input_reset(1'b0), // @[:@2882.4]
    .io_input_enable(valid_up), // @[:@2882.4]
    .io_output_counts_1(io_output_counts_1), // @[:@2882.4]
    .io_output_counts_0(io_output_counts_0), // @[:@2882.4]
    .io_output_oobs_0(io_output_oobs_0), // @[:@2882.4]
    .io_output_oobs_1(io_output_oobs_1), // @[:@2882.4]
    .io_output_done(dontcare2) // @[:@2882.4]
  );

endmodule


module RetimeShiftRegister
#(
    parameter WIDTH = 1,
    parameter STAGES = 1)
(
    input clock,
    input reset,
    input flow,
    input [WIDTH-1:0] init,
    input [WIDTH-1:0] in,
    output reg [WIDTH-1:0] out
);
  integer i;
  reg [WIDTH-1:0] sr[STAGES:0]; // Create 'STAGES' number of register, each 'WIDTH' bits wide

   /* synopsys dc_tcl_script_begin
    set_ungroup [current_design] true
    set_flatten true -effort high -phase true -design [current_design]
    set_dont_retime [current_design] false
    set_optimize_registers true -design [current_design]
    */
  always @(posedge clock) begin
    if (reset) begin
      for(i=0; i<STAGES; i=i+1) begin
        sr[i] <= init;
      end
    end else begin
      if (flow) begin 
        sr[0] <= in;
        for(i=1; i<STAGES; i=i+1) begin
          sr[i] <= sr[i-1];
        end
      end
    end
  end

  always @(*) begin
    out = sr[STAGES-1];
  end
endmodule


// End boilerplate
module FF( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output [31:0] io_rPort_0_output_0, // @[:@6.4]
  input  [31:0] io_wPort_0_data_0, // @[:@6.4]
  input         io_wPort_0_reset // @[:@6.4]
);
  reg [31:0] ff; // @[MemPrimitives.scala 321:19:@21.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_69; // @[MemPrimitives.scala 325:12:@24.4]
  assign _T_69 = io_wPort_0_reset ? 32'h0 : io_wPort_0_data_0; // @[MemPrimitives.scala 325:12:@24.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@26.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 32'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 32'h0;
      end else begin
        ff <= io_wPort_0_data_0;
      end
    end
  end
endmodule
module SRFF( // @[:@28.2]
  input   clock, // @[:@29.4]
  input   reset, // @[:@30.4]
  input   io_input_set, // @[:@31.4]
  input   io_input_reset, // @[:@31.4]
  input   io_input_asyn_reset, // @[:@31.4]
  output  io_output // @[:@31.4]
);
  reg  _T_15; // @[SRFF.scala 20:21:@33.4]
  reg [31:0] _RAND_0;
  wire  _T_19; // @[SRFF.scala 21:74:@34.4]
  wire  _T_20; // @[SRFF.scala 21:48:@35.4]
  wire  _T_21; // @[SRFF.scala 21:14:@36.4]
  assign _T_19 = io_input_reset ? 1'h0 : _T_15; // @[SRFF.scala 21:74:@34.4]
  assign _T_20 = io_input_set ? 1'h1 : _T_19; // @[SRFF.scala 21:48:@35.4]
  assign _T_21 = io_input_asyn_reset ? 1'h0 : _T_20; // @[SRFF.scala 21:14:@36.4]
  assign io_output = io_input_asyn_reset ? 1'h0 : _T_15; // @[SRFF.scala 22:15:@39.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_15 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_15 <= 1'h0;
    end else begin
      if (io_input_asyn_reset) begin
        _T_15 <= 1'h0;
      end else begin
        if (io_input_set) begin
          _T_15 <= 1'h1;
        end else begin
          if (io_input_reset) begin
            _T_15 <= 1'h0;
          end
        end
      end
    end
  end
endmodule
module SingleCounter( // @[:@41.2]
  input   clock, // @[:@42.4]
  input   reset, // @[:@43.4]
  input   io_input_reset, // @[:@44.4]
  output  io_output_done // @[:@44.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@57.4]
  wire [31:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@57.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@57.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@73.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@73.4]
  wire [31:0] _T_48; // @[Counter.scala 287:52:@101.4]
  wire [32:0] _T_50; // @[Counter.scala 291:33:@102.4]
  wire [31:0] _T_51; // @[Counter.scala 291:33:@103.4]
  wire [31:0] _T_52; // @[Counter.scala 291:33:@104.4]
  wire  _T_57; // @[Counter.scala 293:18:@106.4]
  wire [31:0] _T_68; // @[Counter.scala 299:115:@114.4]
  wire [31:0] _T_71; // @[Counter.scala 299:152:@117.4]
  wire [31:0] _T_72; // @[Counter.scala 299:74:@118.4]
  FF bases_0 ( // @[Counter.scala 261:53:@57.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@73.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@101.4]
  assign _T_50 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@102.4]
  assign _T_51 = $signed(_T_48) + $signed(32'sh1); // @[Counter.scala 291:33:@103.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@104.4]
  assign _T_57 = $signed(_T_52) >= $signed(32'sh1e); // @[Counter.scala 293:18:@106.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@114.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@117.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@118.4]
  assign io_output_done = $signed(_T_52) >= $signed(32'sh1e); // @[Counter.scala 333:20:@127.4]
  assign bases_0_clock = clock; // @[:@58.4]
  assign bases_0_reset = reset; // @[:@59.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 32'h0 : _T_72; // @[Counter.scala 299:31:@120.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@99.4]
  assign SRFF_clock = clock; // @[:@74.4]
  assign SRFF_reset = reset; // @[:@75.4]
  assign SRFF_io_input_set = io_input_reset == 1'h0; // @[Counter.scala 264:23:@78.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@80.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@81.4]
endmodule
module RetimeWrapper( // @[:@144.2]
  input   clock, // @[:@145.4]
  input   reset, // @[:@146.4]
  input   io_flow, // @[:@147.4]
  input   io_in, // @[:@147.4]
  output  io_out // @[:@147.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@149.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@149.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@149.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@162.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@161.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@160.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@159.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@158.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@156.4]
endmodule
module RootController_sm( // @[:@312.2]
  input   clock, // @[:@313.4]
  input   reset, // @[:@314.4]
  input   io_enable, // @[:@315.4]
  output  io_done, // @[:@315.4]
  input   io_rst, // @[:@315.4]
  input   io_ctrDone, // @[:@315.4]
  output  io_ctrInc, // @[:@315.4]
  input   io_parentAck, // @[:@315.4]
  input   io_doneIn_0, // @[:@315.4]
  output  io_enableOut_0, // @[:@315.4]
  output  io_childAck_0 // @[:@315.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@318.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@318.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@321.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@321.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@338.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@338.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@357.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@416.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@433.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@433.4]
  wire  finished; // @[Controllers.scala 81:26:@324.4]
  wire  _T_81; // @[Controllers.scala 86:43:@328.4]
  wire  synchronize; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  wire  _T_93; // @[Controllers.scala 92:52:@342.4]
  wire  _T_122; // @[Controllers.scala 128:33:@371.4]
  wire  _T_124; // @[Controllers.scala 128:54:@372.4]
  wire  _T_125; // @[Controllers.scala 128:52:@373.4]
  wire  _T_126; // @[Controllers.scala 128:66:@374.4]
  wire  _T_128; // @[Controllers.scala 128:98:@376.4]
  wire  _T_129; // @[Controllers.scala 128:96:@377.4]
  wire  _T_131; // @[Controllers.scala 128:123:@378.4]
  wire  _T_133; // @[Controllers.scala 129:48:@381.4]
  wire  _T_134; // @[Controllers.scala 129:57:@382.4]
  wire  _T_138; // @[Controllers.scala 130:52:@386.4]
  wire  _T_139; // @[Controllers.scala 130:50:@387.4]
  wire  _T_147; // @[Controllers.scala 130:129:@393.4]
  wire  _T_150; // @[Controllers.scala 131:45:@396.4]
  wire  _T_154; // @[Controllers.scala 213:68:@402.4]
  wire  _T_156; // @[Controllers.scala 213:90:@404.4]
  wire  _T_158; // @[Controllers.scala 213:132:@406.4]
  wire  _T_159; // @[Controllers.scala 213:130:@407.4]
  wire  _T_160; // @[Controllers.scala 213:156:@408.4]
  reg  _T_166; // @[package.scala 48:56:@412.4]
  reg [31:0] _RAND_0;
  wire  _T_167; // @[package.scala 100:41:@414.4]
  reg  _T_180; // @[package.scala 48:56:@430.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@318.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@321.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@338.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@357.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@416.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@433.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  assign finished = done_0_io_output | io_done; // @[Controllers.scala 81:26:@324.4]
  assign _T_81 = io_rst | done_0_io_output; // @[Controllers.scala 86:43:@328.4]
  assign synchronize = RetimeWrapper_io_out; // @[package.scala 96:25:@362.4 package.scala 96:25:@363.4]
  assign _T_93 = synchronize | io_rst; // @[Controllers.scala 92:52:@342.4]
  assign _T_122 = done_0_io_output == 1'h0; // @[Controllers.scala 128:33:@371.4]
  assign _T_124 = io_ctrDone == 1'h0; // @[Controllers.scala 128:54:@372.4]
  assign _T_125 = _T_122 & _T_124; // @[Controllers.scala 128:52:@373.4]
  assign _T_126 = _T_125 & io_enable; // @[Controllers.scala 128:66:@374.4]
  assign _T_128 = ~ iterDone_0_io_output; // @[Controllers.scala 128:98:@376.4]
  assign _T_129 = _T_126 & _T_128; // @[Controllers.scala 128:96:@377.4]
  assign _T_131 = io_doneIn_0 == 1'h0; // @[Controllers.scala 128:123:@378.4]
  assign _T_133 = io_doneIn_0 | io_rst; // @[Controllers.scala 129:48:@381.4]
  assign _T_134 = _T_133 | io_parentAck; // @[Controllers.scala 129:57:@382.4]
  assign _T_138 = synchronize == 1'h0; // @[Controllers.scala 130:52:@386.4]
  assign _T_139 = io_doneIn_0 & _T_138; // @[Controllers.scala 130:50:@387.4]
  assign _T_147 = finished == 1'h0; // @[Controllers.scala 130:129:@393.4]
  assign _T_150 = io_rst == 1'h0; // @[Controllers.scala 131:45:@396.4]
  assign _T_154 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@402.4]
  assign _T_156 = _T_154 & _T_128; // @[Controllers.scala 213:90:@404.4]
  assign _T_158 = ~ done_0_io_output; // @[Controllers.scala 213:132:@406.4]
  assign _T_159 = _T_156 & _T_158; // @[Controllers.scala 213:130:@407.4]
  assign _T_160 = ~ io_ctrDone; // @[Controllers.scala 213:156:@408.4]
  assign _T_167 = done_0_io_output & _T_166; // @[package.scala 100:41:@414.4]
  assign io_done = RetimeWrapper_2_io_out; // @[Controllers.scala 245:13:@440.4]
  assign io_ctrInc = io_doneIn_0; // @[Controllers.scala 122:17:@356.4]
  assign io_enableOut_0 = _T_159 & _T_160; // @[Controllers.scala 213:55:@410.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@401.4]
  assign active_0_clock = clock; // @[:@319.4]
  assign active_0_reset = reset; // @[:@320.4]
  assign active_0_io_input_set = _T_129 & _T_131; // @[Controllers.scala 128:30:@380.4]
  assign active_0_io_input_reset = _T_134 | done_0_io_output; // @[Controllers.scala 129:32:@385.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@326.4]
  assign done_0_clock = clock; // @[:@322.4]
  assign done_0_reset = reset; // @[:@323.4]
  assign done_0_io_input_set = io_ctrDone & _T_150; // @[Controllers.scala 131:28:@399.4]
  assign done_0_io_input_reset = _T_81 | io_parentAck; // @[Controllers.scala 86:33:@336.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@327.4]
  assign iterDone_0_clock = clock; // @[:@339.4]
  assign iterDone_0_reset = reset; // @[:@340.4]
  assign iterDone_0_io_input_set = _T_139 & _T_147; // @[Controllers.scala 130:32:@395.4]
  assign iterDone_0_io_input_reset = _T_93 | io_parentAck; // @[Controllers.scala 92:37:@350.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@341.4]
  assign RetimeWrapper_clock = clock; // @[:@358.4]
  assign RetimeWrapper_reset = reset; // @[:@359.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@361.4]
  assign RetimeWrapper_io_in = io_doneIn_0; // @[package.scala 94:16:@360.4]
  assign RetimeWrapper_1_clock = clock; // @[:@417.4]
  assign RetimeWrapper_1_reset = reset; // @[:@418.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@420.4]
  assign RetimeWrapper_1_io_in = _T_167 | io_parentAck; // @[package.scala 94:16:@419.4]
  assign RetimeWrapper_2_clock = clock; // @[:@434.4]
  assign RetimeWrapper_2_reset = reset; // @[:@435.4]
  assign RetimeWrapper_2_io_flow = io_enable; // @[package.scala 95:18:@437.4]
  assign RetimeWrapper_2_io_in = done_0_io_output & _T_180; // @[package.scala 94:16:@436.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_166 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_180 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_166 <= 1'h0;
    end else begin
      _T_166 <= _T_122;
    end
    if (reset) begin
      _T_180 <= 1'h0;
    end else begin
      _T_180 <= _T_122;
    end
  end
endmodule
module SRAM( // @[:@507.2]
  input         clock, // @[:@508.4]
  input  [20:0] io_raddr, // @[:@510.4]
  output [31:0] io_rdata, // @[:@510.4]
  input         io_backpressure // @[:@510.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@512.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@512.4]
  wire [20:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@512.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@512.4]
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(2073600), .AWIDTH(21)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@512.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign io_rdata = SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@539.4]
  assign SRAMVerilogAWS_wdata = 32'h0; // @[SRAM.scala 175:20:@526.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@527.4]
  assign SRAMVerilogAWS_wen = 1'h0; // @[SRAM.scala 173:18:@524.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@529.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@528.4]
  assign SRAMVerilogAWS_waddr = 21'h0; // @[SRAM.scala 174:20:@525.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@523.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@522.4]
endmodule
module RetimeWrapper_5( // @[:@553.2]
  input         clock, // @[:@554.4]
  input         reset, // @[:@555.4]
  input         io_flow, // @[:@556.4]
  input  [20:0] io_in, // @[:@556.4]
  output [20:0] io_out // @[:@556.4]
);
  wire [20:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire [20:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@558.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@558.4]
  RetimeShiftRegister #(.WIDTH(21), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@558.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@571.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@570.4]
  assign sr_init = 21'h0; // @[RetimeShiftRegister.scala 19:16:@569.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@568.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@567.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@565.4]
endmodule
module Mem1D( // @[:@573.2]
  input         clock, // @[:@574.4]
  input         reset, // @[:@575.4]
  input  [20:0] io_r_ofs_0, // @[:@576.4]
  input         io_r_backpressure, // @[:@576.4]
  output [31:0] io_output // @[:@576.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@580.4]
  wire [20:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@580.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@580.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@580.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@583.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_in; // @[package.scala 93:22:@583.4]
  wire [20:0] RetimeWrapper_io_out; // @[package.scala 93:22:@583.4]
  SRAM SRAM ( // @[MemPrimitives.scala 715:21:@580.4]
    .clock(SRAM_clock),
    .io_raddr(SRAM_io_raddr),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_5 RetimeWrapper ( // @[package.scala 93:22:@583.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@596.4]
  assign SRAM_clock = clock; // @[:@581.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@590.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@595.4]
  assign RetimeWrapper_clock = clock; // @[:@584.4]
  assign RetimeWrapper_reset = reset; // @[:@585.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@587.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@586.4]
endmodule
module StickySelects( // @[:@598.2]
  input   io_ins_0, // @[:@601.4]
  output  io_outs_0 // @[:@601.4]
);
  assign io_outs_0 = io_ins_0; // @[StickySelects.scala 34:26:@603.4]
endmodule
module RetimeWrapper_6( // @[:@617.2]
  input   clock, // @[:@618.4]
  input   reset, // @[:@619.4]
  input   io_flow, // @[:@620.4]
  input   io_in, // @[:@620.4]
  output  io_out // @[:@620.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@622.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@622.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@622.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@635.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@634.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@633.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@632.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@631.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@629.4]
endmodule
module x223_outbuf_0( // @[:@637.2]
  input         clock, // @[:@638.4]
  input         reset, // @[:@639.4]
  input  [20:0] io_rPort_0_ofs_0, // @[:@640.4]
  input         io_rPort_0_en_0, // @[:@640.4]
  input         io_rPort_0_backpressure, // @[:@640.4]
  output [31:0] io_rPort_0_output_0 // @[:@640.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@655.4]
  wire [20:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@655.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@655.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@655.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@681.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@695.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@695.4]
  wire  _T_76; // @[MemPrimitives.scala 126:35:@685.4]
  wire [22:0] _T_78; // @[Cat.scala 30:58:@687.4]
  Mem1D Mem1D ( // @[MemPrimitives.scala 64:21:@655.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_output(Mem1D_io_output)
  );
  StickySelects StickySelects ( // @[MemPrimitives.scala 124:33:@681.4]
    .io_ins_0(StickySelects_io_ins_0),
    .io_outs_0(StickySelects_io_outs_0)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@695.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_76 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@685.4]
  assign _T_78 = {_T_76,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@687.4]
  assign io_rPort_0_output_0 = Mem1D_io_output; // @[MemPrimitives.scala 152:13:@702.4]
  assign Mem1D_clock = clock; // @[:@656.4]
  assign Mem1D_reset = reset; // @[:@657.4]
  assign Mem1D_io_r_ofs_0 = _T_78[20:0]; // @[MemPrimitives.scala 131:28:@691.4]
  assign Mem1D_io_r_backpressure = _T_78[21]; // @[MemPrimitives.scala 132:32:@692.4]
  assign StickySelects_io_ins_0 = io_rPort_0_en_0; // @[MemPrimitives.scala 125:64:@684.4]
  assign RetimeWrapper_clock = clock; // @[:@696.4]
  assign RetimeWrapper_reset = reset; // @[:@697.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@699.4]
  assign RetimeWrapper_io_in = io_rPort_0_en_0; // @[package.scala 94:16:@698.4]
endmodule
module x478_sm( // @[:@846.2]
  input   clock, // @[:@847.4]
  input   reset, // @[:@848.4]
  input   io_enable, // @[:@849.4]
  output  io_done, // @[:@849.4]
  input   io_ctrDone, // @[:@849.4]
  output  io_ctrInc, // @[:@849.4]
  input   io_parentAck, // @[:@849.4]
  input   io_doneIn_0, // @[:@849.4]
  input   io_doneIn_1, // @[:@849.4]
  output  io_enableOut_0, // @[:@849.4]
  output  io_enableOut_1, // @[:@849.4]
  output  io_childAck_0, // @[:@849.4]
  output  io_childAck_1 // @[:@849.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@852.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@852.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@855.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@855.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@858.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@858.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@861.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@861.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@890.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@893.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@893.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@994.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1011.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1011.4]
  wire  allDone; // @[Controllers.scala 80:47:@864.4]
  wire  synchronize; // @[Controllers.scala 146:56:@918.4]
  wire  _T_127; // @[Controllers.scala 150:35:@920.4]
  wire  _T_129; // @[Controllers.scala 150:60:@921.4]
  wire  _T_130; // @[Controllers.scala 150:58:@922.4]
  wire  _T_132; // @[Controllers.scala 150:76:@923.4]
  wire  _T_133; // @[Controllers.scala 150:74:@924.4]
  wire  _T_135; // @[Controllers.scala 150:97:@925.4]
  wire  _T_136; // @[Controllers.scala 150:95:@926.4]
  wire  _T_152; // @[Controllers.scala 150:35:@944.4]
  wire  _T_154; // @[Controllers.scala 150:60:@945.4]
  wire  _T_155; // @[Controllers.scala 150:58:@946.4]
  wire  _T_157; // @[Controllers.scala 150:76:@947.4]
  wire  _T_158; // @[Controllers.scala 150:74:@948.4]
  wire  _T_161; // @[Controllers.scala 150:95:@950.4]
  wire  _T_179; // @[Controllers.scala 213:68:@972.4]
  wire  _T_181; // @[Controllers.scala 213:90:@974.4]
  wire  _T_183; // @[Controllers.scala 213:132:@976.4]
  wire  _T_184; // @[Controllers.scala 213:130:@977.4]
  wire  _T_185; // @[Controllers.scala 213:156:@978.4]
  wire  _T_187; // @[Controllers.scala 213:68:@981.4]
  wire  _T_189; // @[Controllers.scala 213:90:@983.4]
  wire  _T_196; // @[package.scala 100:49:@989.4]
  reg  _T_199; // @[package.scala 48:56:@990.4]
  reg [31:0] _RAND_0;
  wire  _T_200; // @[package.scala 100:41:@992.4]
  reg  _T_213; // @[package.scala 48:56:@1008.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@852.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@855.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@858.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@861.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@890.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@893.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@994.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1011.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@864.4]
  assign synchronize = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 146:56:@918.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 150:35:@920.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 150:60:@921.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 150:58:@922.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 150:76:@923.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 150:74:@924.4]
  assign _T_135 = io_ctrDone == 1'h0; // @[Controllers.scala 150:97:@925.4]
  assign _T_136 = _T_133 & _T_135; // @[Controllers.scala 150:95:@926.4]
  assign _T_152 = ~ iterDone_1_io_output; // @[Controllers.scala 150:35:@944.4]
  assign _T_154 = io_doneIn_1 == 1'h0; // @[Controllers.scala 150:60:@945.4]
  assign _T_155 = _T_152 & _T_154; // @[Controllers.scala 150:58:@946.4]
  assign _T_157 = done_1_io_output == 1'h0; // @[Controllers.scala 150:76:@947.4]
  assign _T_158 = _T_155 & _T_157; // @[Controllers.scala 150:74:@948.4]
  assign _T_161 = _T_158 & _T_135; // @[Controllers.scala 150:95:@950.4]
  assign _T_179 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@972.4]
  assign _T_181 = _T_179 & _T_127; // @[Controllers.scala 213:90:@974.4]
  assign _T_183 = ~ allDone; // @[Controllers.scala 213:132:@976.4]
  assign _T_184 = _T_181 & _T_183; // @[Controllers.scala 213:130:@977.4]
  assign _T_185 = ~ io_ctrDone; // @[Controllers.scala 213:156:@978.4]
  assign _T_187 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@981.4]
  assign _T_189 = _T_187 & _T_152; // @[Controllers.scala 213:90:@983.4]
  assign _T_196 = allDone == 1'h0; // @[package.scala 100:49:@989.4]
  assign _T_200 = allDone & _T_199; // @[package.scala 100:41:@992.4]
  assign io_done = RetimeWrapper_1_io_out; // @[Controllers.scala 245:13:@1018.4]
  assign io_ctrInc = iterDone_0_io_output & iterDone_1_io_output; // @[Controllers.scala 143:17:@917.4]
  assign io_enableOut_0 = _T_184 & _T_185; // @[Controllers.scala 213:55:@980.4]
  assign io_enableOut_1 = _T_189 & _T_183; // @[Controllers.scala 213:55:@988.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@969.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@971.4]
  assign active_0_clock = clock; // @[:@853.4]
  assign active_0_reset = reset; // @[:@854.4]
  assign active_0_io_input_set = _T_136 & io_enable; // @[Controllers.scala 150:32:@929.4]
  assign active_0_io_input_reset = io_doneIn_0 | io_parentAck; // @[Controllers.scala 151:34:@933.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@867.4]
  assign active_1_clock = clock; // @[:@856.4]
  assign active_1_reset = reset; // @[:@857.4]
  assign active_1_io_input_set = _T_161 & io_enable; // @[Controllers.scala 150:32:@953.4]
  assign active_1_io_input_reset = io_doneIn_1 | io_parentAck; // @[Controllers.scala 151:34:@957.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@868.4]
  assign done_0_clock = clock; // @[:@859.4]
  assign done_0_reset = reset; // @[:@860.4]
  assign done_0_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@943.4]
  assign done_0_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@879.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@869.4]
  assign done_1_clock = clock; // @[:@862.4]
  assign done_1_reset = reset; // @[:@863.4]
  assign done_1_io_input_set = io_ctrDone; // @[Controllers.scala 153:30:@967.4]
  assign done_1_io_input_reset = allDone | io_parentAck; // @[Controllers.scala 86:33:@888.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@870.4]
  assign iterDone_0_clock = clock; // @[:@891.4]
  assign iterDone_0_reset = reset; // @[:@892.4]
  assign iterDone_0_io_input_set = io_doneIn_0; // @[Controllers.scala 152:34:@939.4]
  assign iterDone_0_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@896.4]
  assign iterDone_1_clock = clock; // @[:@894.4]
  assign iterDone_1_reset = reset; // @[:@895.4]
  assign iterDone_1_io_input_set = io_doneIn_1; // @[Controllers.scala 152:34:@963.4]
  assign iterDone_1_io_input_reset = synchronize | io_parentAck; // @[Controllers.scala 92:37:@915.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@897.4]
  assign RetimeWrapper_clock = clock; // @[:@995.4]
  assign RetimeWrapper_reset = reset; // @[:@996.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@998.4]
  assign RetimeWrapper_io_in = _T_200 | io_parentAck; // @[package.scala 94:16:@997.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1012.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1013.4]
  assign RetimeWrapper_1_io_flow = io_enable; // @[package.scala 95:18:@1015.4]
  assign RetimeWrapper_1_io_in = allDone & _T_213; // @[package.scala 94:16:@1014.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_199 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_213 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_199 <= 1'h0;
    end else begin
      _T_199 <= _T_196;
    end
    if (reset) begin
      _T_213 <= 1'h0;
    end else begin
      _T_213 <= _T_196;
    end
  end
endmodule
module x403_outr_UnitPipe_sm( // @[:@1435.2]
  input   clock, // @[:@1436.4]
  input   reset, // @[:@1437.4]
  input   io_enable, // @[:@1438.4]
  output  io_done, // @[:@1438.4]
  input   io_parentAck, // @[:@1438.4]
  input   io_doneIn_0, // @[:@1438.4]
  input   io_doneIn_1, // @[:@1438.4]
  output  io_enableOut_0, // @[:@1438.4]
  output  io_enableOut_1, // @[:@1438.4]
  output  io_childAck_0, // @[:@1438.4]
  output  io_childAck_1, // @[:@1438.4]
  input   io_ctrCopyDone_0, // @[:@1438.4]
  input   io_ctrCopyDone_1 // @[:@1438.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@1441.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@1441.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@1444.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@1444.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@1447.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@1447.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@1450.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@1450.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@1479.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@1482.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@1482.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@1523.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@1537.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@1555.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@1592.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@1606.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@1624.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@1671.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@1688.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@1688.4]
  wire  allDone; // @[Controllers.scala 80:47:@1453.4]
  wire  _T_127; // @[Controllers.scala 165:35:@1507.4]
  wire  _T_129; // @[Controllers.scala 165:60:@1508.4]
  wire  _T_130; // @[Controllers.scala 165:58:@1509.4]
  wire  _T_132; // @[Controllers.scala 165:76:@1510.4]
  wire  _T_133; // @[Controllers.scala 165:74:@1511.4]
  wire  _T_137; // @[Controllers.scala 165:109:@1514.4]
  wire  _T_140; // @[Controllers.scala 165:141:@1516.4]
  wire  _T_148; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  wire  _T_152; // @[Controllers.scala 167:54:@1531.4]
  wire  _T_153; // @[Controllers.scala 167:52:@1532.4]
  wire  _T_160; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  wire  _T_178; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  wire  _T_182; // @[Controllers.scala 169:67:@1563.4]
  wire  _T_183; // @[Controllers.scala 169:86:@1564.4]
  wire  _T_195; // @[Controllers.scala 165:35:@1576.4]
  wire  _T_197; // @[Controllers.scala 165:60:@1577.4]
  wire  _T_198; // @[Controllers.scala 165:58:@1578.4]
  wire  _T_200; // @[Controllers.scala 165:76:@1579.4]
  wire  _T_201; // @[Controllers.scala 165:74:@1580.4]
  wire  _T_205; // @[Controllers.scala 165:109:@1583.4]
  wire  _T_208; // @[Controllers.scala 165:141:@1585.4]
  wire  _T_216; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  wire  _T_220; // @[Controllers.scala 167:54:@1600.4]
  wire  _T_221; // @[Controllers.scala 167:52:@1601.4]
  wire  _T_228; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  wire  _T_246; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  wire  _T_250; // @[Controllers.scala 169:67:@1632.4]
  wire  _T_251; // @[Controllers.scala 169:86:@1633.4]
  wire  _T_265; // @[Controllers.scala 213:68:@1649.4]
  wire  _T_267; // @[Controllers.scala 213:90:@1651.4]
  wire  _T_269; // @[Controllers.scala 213:132:@1653.4]
  wire  _T_273; // @[Controllers.scala 213:68:@1658.4]
  wire  _T_275; // @[Controllers.scala 213:90:@1660.4]
  wire  _T_282; // @[package.scala 100:49:@1666.4]
  reg  _T_285; // @[package.scala 48:56:@1667.4]
  reg [31:0] _RAND_0;
  wire  _T_286; // @[package.scala 100:41:@1669.4]
  reg  _T_299; // @[package.scala 48:56:@1685.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@1441.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@1444.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@1447.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@1450.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@1479.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@1482.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@1523.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@1537.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@1555.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@1592.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@1606.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@1624.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@1671.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@1688.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  assign allDone = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@1453.4]
  assign _T_127 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@1507.4]
  assign _T_129 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@1508.4]
  assign _T_130 = _T_127 & _T_129; // @[Controllers.scala 165:58:@1509.4]
  assign _T_132 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@1510.4]
  assign _T_133 = _T_130 & _T_132; // @[Controllers.scala 165:74:@1511.4]
  assign _T_137 = _T_133 & io_enable; // @[Controllers.scala 165:109:@1514.4]
  assign _T_140 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@1516.4]
  assign _T_148 = RetimeWrapper_io_out; // @[package.scala 96:25:@1528.4 package.scala 96:25:@1529.4]
  assign _T_152 = _T_148 == 1'h0; // @[Controllers.scala 167:54:@1531.4]
  assign _T_153 = io_doneIn_0 | _T_152; // @[Controllers.scala 167:52:@1532.4]
  assign _T_160 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@1542.4 package.scala 96:25:@1543.4]
  assign _T_178 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@1560.4 package.scala 96:25:@1561.4]
  assign _T_182 = _T_178 == 1'h0; // @[Controllers.scala 169:67:@1563.4]
  assign _T_183 = _T_182 & io_enable; // @[Controllers.scala 169:86:@1564.4]
  assign _T_195 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@1576.4]
  assign _T_197 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@1577.4]
  assign _T_198 = _T_195 & _T_197; // @[Controllers.scala 165:58:@1578.4]
  assign _T_200 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@1579.4]
  assign _T_201 = _T_198 & _T_200; // @[Controllers.scala 165:74:@1580.4]
  assign _T_205 = _T_201 & io_enable; // @[Controllers.scala 165:109:@1583.4]
  assign _T_208 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@1585.4]
  assign _T_216 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@1597.4 package.scala 96:25:@1598.4]
  assign _T_220 = _T_216 == 1'h0; // @[Controllers.scala 167:54:@1600.4]
  assign _T_221 = io_doneIn_1 | _T_220; // @[Controllers.scala 167:52:@1601.4]
  assign _T_228 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@1611.4 package.scala 96:25:@1612.4]
  assign _T_246 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@1629.4 package.scala 96:25:@1630.4]
  assign _T_250 = _T_246 == 1'h0; // @[Controllers.scala 169:67:@1632.4]
  assign _T_251 = _T_250 & io_enable; // @[Controllers.scala 169:86:@1633.4]
  assign _T_265 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@1649.4]
  assign _T_267 = _T_265 & _T_127; // @[Controllers.scala 213:90:@1651.4]
  assign _T_269 = ~ allDone; // @[Controllers.scala 213:132:@1653.4]
  assign _T_273 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@1658.4]
  assign _T_275 = _T_273 & _T_195; // @[Controllers.scala 213:90:@1660.4]
  assign _T_282 = allDone == 1'h0; // @[package.scala 100:49:@1666.4]
  assign _T_286 = allDone & _T_285; // @[package.scala 100:41:@1669.4]
  assign io_done = RetimeWrapper_7_io_out; // @[Controllers.scala 245:13:@1695.4]
  assign io_enableOut_0 = _T_267 & _T_269; // @[Controllers.scala 213:55:@1657.4]
  assign io_enableOut_1 = _T_275 & _T_269; // @[Controllers.scala 213:55:@1665.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@1646.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@1648.4]
  assign active_0_clock = clock; // @[:@1442.4]
  assign active_0_reset = reset; // @[:@1443.4]
  assign active_0_io_input_set = _T_137 & _T_140; // @[Controllers.scala 165:32:@1518.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@1522.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1456.4]
  assign active_1_clock = clock; // @[:@1445.4]
  assign active_1_reset = reset; // @[:@1446.4]
  assign active_1_io_input_set = _T_205 & _T_208; // @[Controllers.scala 165:32:@1587.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@1591.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@1457.4]
  assign done_0_clock = clock; // @[:@1448.4]
  assign done_0_reset = reset; // @[:@1449.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_183; // @[Controllers.scala 169:30:@1568.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1468.4 Controllers.scala 170:32:@1575.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1458.4]
  assign done_1_clock = clock; // @[:@1451.4]
  assign done_1_reset = reset; // @[:@1452.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_251; // @[Controllers.scala 169:30:@1637.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@1477.4 Controllers.scala 170:32:@1644.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@1459.4]
  assign iterDone_0_clock = clock; // @[:@1480.4]
  assign iterDone_0_reset = reset; // @[:@1481.4]
  assign iterDone_0_io_input_set = _T_153 & io_enable; // @[Controllers.scala 167:34:@1536.4]
  assign iterDone_0_io_input_reset = _T_160 | io_parentAck; // @[Controllers.scala 92:37:@1495.4 Controllers.scala 168:36:@1552.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1485.4]
  assign iterDone_1_clock = clock; // @[:@1483.4]
  assign iterDone_1_reset = reset; // @[:@1484.4]
  assign iterDone_1_io_input_set = _T_221 & io_enable; // @[Controllers.scala 167:34:@1605.4]
  assign iterDone_1_io_input_reset = _T_228 | io_parentAck; // @[Controllers.scala 92:37:@1504.4 Controllers.scala 168:36:@1621.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@1486.4]
  assign RetimeWrapper_clock = clock; // @[:@1524.4]
  assign RetimeWrapper_reset = reset; // @[:@1525.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@1527.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@1526.4]
  assign RetimeWrapper_1_clock = clock; // @[:@1538.4]
  assign RetimeWrapper_1_reset = reset; // @[:@1539.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@1541.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@1540.4]
  assign RetimeWrapper_2_clock = clock; // @[:@1556.4]
  assign RetimeWrapper_2_reset = reset; // @[:@1557.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@1559.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@1558.4]
  assign RetimeWrapper_3_clock = clock; // @[:@1593.4]
  assign RetimeWrapper_3_reset = reset; // @[:@1594.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@1596.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@1595.4]
  assign RetimeWrapper_4_clock = clock; // @[:@1607.4]
  assign RetimeWrapper_4_reset = reset; // @[:@1608.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@1610.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@1609.4]
  assign RetimeWrapper_5_clock = clock; // @[:@1625.4]
  assign RetimeWrapper_5_reset = reset; // @[:@1626.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@1628.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@1627.4]
  assign RetimeWrapper_6_clock = clock; // @[:@1672.4]
  assign RetimeWrapper_6_reset = reset; // @[:@1673.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@1675.4]
  assign RetimeWrapper_6_io_in = _T_286 | io_parentAck; // @[package.scala 94:16:@1674.4]
  assign RetimeWrapper_7_clock = clock; // @[:@1689.4]
  assign RetimeWrapper_7_reset = reset; // @[:@1690.4]
  assign RetimeWrapper_7_io_flow = io_enable; // @[package.scala 95:18:@1692.4]
  assign RetimeWrapper_7_io_in = allDone & _T_299; // @[package.scala 94:16:@1691.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_285 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_299 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_285 <= 1'h0;
    end else begin
      _T_285 <= _T_282;
    end
    if (reset) begin
      _T_299 <= 1'h0;
    end else begin
      _T_299 <= _T_282;
    end
  end
endmodule
module CompactingIncDincCtr( // @[:@1924.2]
  input   clock, // @[:@1925.4]
  input   reset, // @[:@1926.4]
  input   io_input_inc_en_0, // @[:@1927.4]
  input   io_input_dinc_en_0, // @[:@1927.4]
  output  io_output_full // @[:@1927.4]
);
  reg [31:0] cnt; // @[Counter.scala 170:20:@1929.4]
  reg [31:0] _RAND_0;
  wire [14:0] numPushed; // @[Counter.scala 172:47:@1930.4]
  wire [14:0] numPopped; // @[Counter.scala 173:48:@1931.4]
  wire [31:0] _GEN_0; // @[Counter.scala 174:14:@1932.4]
  wire [32:0] _T_37; // @[Counter.scala 174:14:@1932.4]
  wire [31:0] _T_38; // @[Counter.scala 174:14:@1933.4]
  wire [31:0] _T_39; // @[Counter.scala 174:14:@1934.4]
  wire [31:0] _GEN_1; // @[Counter.scala 174:26:@1935.4]
  wire [32:0] _T_40; // @[Counter.scala 174:26:@1935.4]
  wire [31:0] _T_41; // @[Counter.scala 174:26:@1936.4]
  wire [31:0] _T_42; // @[Counter.scala 174:26:@1937.4]
  assign numPushed = io_input_inc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 172:47:@1930.4]
  assign numPopped = io_input_dinc_en_0 ? $signed(15'sh1) : $signed(15'sh0); // @[Counter.scala 173:48:@1931.4]
  assign _GEN_0 = {{17{numPushed[14]}},numPushed}; // @[Counter.scala 174:14:@1932.4]
  assign _T_37 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1932.4]
  assign _T_38 = $signed(cnt) + $signed(_GEN_0); // @[Counter.scala 174:14:@1933.4]
  assign _T_39 = $signed(_T_38); // @[Counter.scala 174:14:@1934.4]
  assign _GEN_1 = {{17{numPopped[14]}},numPopped}; // @[Counter.scala 174:26:@1935.4]
  assign _T_40 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1935.4]
  assign _T_41 = $signed(_T_39) - $signed(_GEN_1); // @[Counter.scala 174:26:@1936.4]
  assign _T_42 = $signed(_T_41); // @[Counter.scala 174:26:@1937.4]
  assign io_output_full = $signed(cnt) > $signed(32'sh1dff); // @[Counter.scala 180:18:@1951.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  cnt = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cnt <= 32'sh0;
    end else begin
      cnt <= _T_42;
    end
  end
endmodule
module x224_fifoinraw_0( // @[:@2074.2]
  input   clock, // @[:@2075.4]
  input   reset // @[:@2076.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2121.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2121.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2121.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign elements_clock = clock; // @[:@2122.4]
  assign elements_reset = reset; // @[:@2123.4]
  assign elements_io_input_inc_en_0 = 1'h0; // @[MemPrimitives.scala 394:79:@2133.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2134.4]
endmodule
module x225_fifoinpacked_0( // @[:@2497.2]
  input   clock, // @[:@2498.4]
  input   reset, // @[:@2499.4]
  input   io_wPort_0_en_0, // @[:@2500.4]
  output  io_full, // @[:@2500.4]
  input   io_active_0_in, // @[:@2500.4]
  output  io_active_0_out // @[:@2500.4]
);
  wire  elements_clock; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_reset; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_inc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_input_dinc_en_0; // @[MemPrimitives.scala 392:24:@2544.4]
  wire  elements_io_output_full; // @[MemPrimitives.scala 392:24:@2544.4]
  CompactingIncDincCtr elements ( // @[MemPrimitives.scala 392:24:@2544.4]
    .clock(elements_clock),
    .reset(elements_reset),
    .io_input_inc_en_0(elements_io_input_inc_en_0),
    .io_input_dinc_en_0(elements_io_input_dinc_en_0),
    .io_output_full(elements_io_output_full)
  );
  assign io_full = elements_io_output_full; // @[MemPrimitives.scala 439:39:@2618.4]
  assign io_active_0_out = io_active_0_in; // @[MemPrimitives.scala 437:129:@2616.4]
  assign elements_clock = clock; // @[:@2545.4]
  assign elements_reset = reset; // @[:@2546.4]
  assign elements_io_input_inc_en_0 = io_wPort_0_en_0; // @[MemPrimitives.scala 394:79:@2556.4]
  assign elements_io_input_dinc_en_0 = 1'h0; // @[MemPrimitives.scala 395:80:@2557.4]
endmodule
module FF_7( // @[:@3047.2]
  input         clock, // @[:@3048.4]
  input         reset, // @[:@3049.4]
  output [12:0] io_rPort_0_output_0, // @[:@3050.4]
  input  [12:0] io_wPort_0_data_0, // @[:@3050.4]
  input         io_wPort_0_reset, // @[:@3050.4]
  input         io_wPort_0_en_0 // @[:@3050.4]
);
  reg [12:0] ff; // @[MemPrimitives.scala 321:19:@3065.4]
  reg [31:0] _RAND_0;
  wire [12:0] _T_68; // @[MemPrimitives.scala 325:32:@3067.4]
  wire [12:0] _T_69; // @[MemPrimitives.scala 325:12:@3068.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@3067.4]
  assign _T_69 = io_wPort_0_reset ? 13'h0 : _T_68; // @[MemPrimitives.scala 325:12:@3068.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@3070.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 13'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 13'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_1( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input         io_setup_saturate, // @[:@3088.4]
  input         io_input_reset, // @[:@3088.4]
  input         io_input_enable, // @[:@3088.4]
  output [12:0] io_output_count_0, // @[:@3088.4]
  output        io_output_oobs_0, // @[:@3088.4]
  output        io_output_done, // @[:@3088.4]
  output        io_output_saturated // @[:@3088.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3101.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3101.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3101.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3117.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3117.4]
  wire  _T_36; // @[Counter.scala 264:45:@3120.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3145.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3146.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3147.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3148.4]
  wire  _T_57; // @[Counter.scala 293:18:@3150.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3158.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3160.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3161.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3162.4]
  wire  _T_75; // @[Counter.scala 322:102:@3166.4]
  wire  _T_77; // @[Counter.scala 322:130:@3167.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3101.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3117.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3120.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3145.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3146.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh1); // @[Counter.scala 291:33:@3147.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3148.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh438); // @[Counter.scala 293:18:@3150.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3158.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3160.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3161.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3162.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3166.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh438); // @[Counter.scala 322:130:@3167.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3165.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3169.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3171.4]
  assign io_output_saturated = io_setup_saturate & _T_57; // @[Counter.scala 340:25:@3174.4]
  assign bases_0_clock = clock; // @[:@3102.4]
  assign bases_0_reset = reset; // @[:@3103.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3164.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3143.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3144.4]
  assign SRFF_clock = clock; // @[:@3118.4]
  assign SRFF_reset = reset; // @[:@3119.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3122.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3124.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3125.4]
endmodule
module SingleCounter_2( // @[:@3214.2]
  input         clock, // @[:@3215.4]
  input         reset, // @[:@3216.4]
  input         io_setup_saturate, // @[:@3217.4]
  input         io_input_reset, // @[:@3217.4]
  input         io_input_enable, // @[:@3217.4]
  output [12:0] io_output_count_0, // @[:@3217.4]
  output        io_output_oobs_0, // @[:@3217.4]
  output        io_output_done // @[:@3217.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@3230.4]
  wire [12:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@3230.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@3230.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@3246.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@3246.4]
  wire  _T_36; // @[Counter.scala 264:45:@3249.4]
  wire [12:0] _T_48; // @[Counter.scala 287:52:@3274.4]
  wire [13:0] _T_50; // @[Counter.scala 291:33:@3275.4]
  wire [12:0] _T_51; // @[Counter.scala 291:33:@3276.4]
  wire [12:0] _T_52; // @[Counter.scala 291:33:@3277.4]
  wire  _T_57; // @[Counter.scala 293:18:@3279.4]
  wire [12:0] _T_68; // @[Counter.scala 299:115:@3287.4]
  wire [12:0] _T_70; // @[Counter.scala 299:85:@3289.4]
  wire [12:0] _T_71; // @[Counter.scala 299:152:@3290.4]
  wire [12:0] _T_72; // @[Counter.scala 299:74:@3291.4]
  wire  _T_75; // @[Counter.scala 322:102:@3295.4]
  wire  _T_77; // @[Counter.scala 322:130:@3296.4]
  FF_7 bases_0 ( // @[Counter.scala 261:53:@3230.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@3246.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@3249.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@3274.4]
  assign _T_50 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3275.4]
  assign _T_51 = $signed(_T_48) + $signed(13'sh2); // @[Counter.scala 291:33:@3276.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@3277.4]
  assign _T_57 = $signed(_T_52) >= $signed(13'sh780); // @[Counter.scala 293:18:@3279.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@3287.4]
  assign _T_70 = io_setup_saturate ? _T_68 : 13'h0; // @[Counter.scala 299:85:@3289.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@3290.4]
  assign _T_72 = _T_57 ? _T_70 : _T_71; // @[Counter.scala 299:74:@3291.4]
  assign _T_75 = $signed(_T_48) < $signed(13'sh0); // @[Counter.scala 322:102:@3295.4]
  assign _T_77 = $signed(_T_48) >= $signed(13'sh780); // @[Counter.scala 322:130:@3296.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@3294.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@3298.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@3300.4]
  assign bases_0_clock = clock; // @[:@3231.4]
  assign bases_0_reset = reset; // @[:@3232.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 13'h0 : _T_72; // @[Counter.scala 299:31:@3293.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@3272.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@3273.4]
  assign SRFF_clock = clock; // @[:@3247.4]
  assign SRFF_reset = reset; // @[:@3248.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@3251.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@3253.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@3254.4]
endmodule
module x229_ctrchain( // @[:@3305.2]
  input         clock, // @[:@3306.4]
  input         reset, // @[:@3307.4]
  input         io_input_reset, // @[:@3308.4]
  input         io_input_enable, // @[:@3308.4]
  output [12:0] io_output_counts_1, // @[:@3308.4]
  output [12:0] io_output_counts_0, // @[:@3308.4]
  output        io_output_oobs_0, // @[:@3308.4]
  output        io_output_oobs_1, // @[:@3308.4]
  output        io_output_done // @[:@3308.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_setup_saturate; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@3310.4]
  wire [12:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_0_io_output_saturated; // @[Counter.scala 513:46:@3310.4]
  wire  ctrs_1_clock; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_setup_saturate; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_reset; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_input_enable; // @[Counter.scala 513:46:@3313.4]
  wire [12:0] ctrs_1_io_output_count_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_oobs_0; // @[Counter.scala 513:46:@3313.4]
  wire  ctrs_1_io_output_done; // @[Counter.scala 513:46:@3313.4]
  wire  isDone; // @[Counter.scala 541:51:@3330.4]
  reg  wasDone; // @[Counter.scala 542:24:@3331.4]
  reg [31:0] _RAND_0;
  wire  _T_64; // @[Counter.scala 546:69:@3339.4]
  wire  _T_66; // @[Counter.scala 546:80:@3340.4]
  reg  doneLatch; // @[Counter.scala 550:26:@3345.4]
  reg [31:0] _RAND_1;
  wire  _T_73; // @[Counter.scala 551:48:@3346.4]
  wire  _T_74; // @[Counter.scala 551:19:@3347.4]
  SingleCounter_1 ctrs_0 ( // @[Counter.scala 513:46:@3310.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_setup_saturate(ctrs_0_io_setup_saturate),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done),
    .io_output_saturated(ctrs_0_io_output_saturated)
  );
  SingleCounter_2 ctrs_1 ( // @[Counter.scala 513:46:@3313.4]
    .clock(ctrs_1_clock),
    .reset(ctrs_1_reset),
    .io_setup_saturate(ctrs_1_io_setup_saturate),
    .io_input_reset(ctrs_1_io_input_reset),
    .io_input_enable(ctrs_1_io_input_enable),
    .io_output_count_0(ctrs_1_io_output_count_0),
    .io_output_oobs_0(ctrs_1_io_output_oobs_0),
    .io_output_done(ctrs_1_io_output_done)
  );
  assign isDone = ctrs_0_io_output_done & ctrs_1_io_output_done; // @[Counter.scala 541:51:@3330.4]
  assign _T_64 = io_input_enable & isDone; // @[Counter.scala 546:69:@3339.4]
  assign _T_66 = wasDone == 1'h0; // @[Counter.scala 546:80:@3340.4]
  assign _T_73 = isDone ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@3346.4]
  assign _T_74 = io_input_reset ? 1'h0 : _T_73; // @[Counter.scala 551:19:@3347.4]
  assign io_output_counts_1 = ctrs_1_io_output_count_0; // @[Counter.scala 557:32:@3352.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@3349.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3351.4]
  assign io_output_oobs_1 = ctrs_1_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@3354.4]
  assign io_output_done = _T_64 & _T_66; // @[Counter.scala 546:18:@3342.4]
  assign ctrs_0_clock = clock; // @[:@3311.4]
  assign ctrs_0_reset = reset; // @[:@3312.4]
  assign ctrs_0_io_setup_saturate = 1'h1; // @[Counter.scala 530:29:@3327.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3319.4]
  assign ctrs_0_io_input_enable = ctrs_1_io_output_done & io_input_enable; // @[Counter.scala 526:29:@3326.4]
  assign ctrs_1_clock = clock; // @[:@3314.4]
  assign ctrs_1_reset = reset; // @[:@3315.4]
  assign ctrs_1_io_setup_saturate = ctrs_0_io_output_saturated; // @[Counter.scala 532:31:@3329.4]
  assign ctrs_1_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@3323.4]
  assign ctrs_1_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@3324.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= isDone;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (isDone) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module RetimeWrapper_21( // @[:@3394.2]
  input   clock, // @[:@3395.4]
  input   reset, // @[:@3396.4]
  input   io_flow, // @[:@3397.4]
  input   io_in, // @[:@3397.4]
  output  io_out // @[:@3397.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3399.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(5)) sr ( // @[RetimeShiftRegister.scala 15:20:@3399.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3412.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3411.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3410.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3409.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3408.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3406.4]
endmodule
module RetimeWrapper_25( // @[:@3522.2]
  input   clock, // @[:@3523.4]
  input   reset, // @[:@3524.4]
  input   io_flow, // @[:@3525.4]
  input   io_in, // @[:@3525.4]
  output  io_out // @[:@3525.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3527.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(4)) sr ( // @[RetimeShiftRegister.scala 15:20:@3527.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3540.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3539.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@3538.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3537.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3536.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3534.4]
endmodule
module x247_inr_Foreach_sm( // @[:@3542.2]
  input   clock, // @[:@3543.4]
  input   reset, // @[:@3544.4]
  input   io_enable, // @[:@3545.4]
  output  io_done, // @[:@3545.4]
  output  io_doneLatch, // @[:@3545.4]
  input   io_ctrDone, // @[:@3545.4]
  output  io_datapathEn, // @[:@3545.4]
  output  io_ctrInc, // @[:@3545.4]
  output  io_ctrRst, // @[:@3545.4]
  input   io_parentAck, // @[:@3545.4]
  input   io_backpressure, // @[:@3545.4]
  input   io_break // @[:@3545.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@3547.4]
  wire  active_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@3547.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@3547.4]
  wire  done_clock; // @[Controllers.scala 262:20:@3550.4]
  wire  done_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@3550.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@3550.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@3584.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@3606.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@3618.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@3626.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@3642.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@3642.4]
  wire  _T_80; // @[Controllers.scala 264:48:@3555.4]
  wire  _T_81; // @[Controllers.scala 264:46:@3556.4]
  wire  _T_82; // @[Controllers.scala 264:62:@3557.4]
  wire  _T_83; // @[Controllers.scala 264:60:@3558.4]
  wire  _T_100; // @[package.scala 100:49:@3575.4]
  reg  _T_103; // @[package.scala 48:56:@3576.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  wire  _T_110; // @[package.scala 100:49:@3591.4]
  reg  _T_113; // @[package.scala 48:56:@3592.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@3594.4]
  wire  _T_118; // @[Controllers.scala 283:41:@3599.4]
  wire  _T_119; // @[Controllers.scala 283:59:@3600.4]
  wire  _T_121; // @[Controllers.scala 284:37:@3603.4]
  wire  _T_124; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  wire  _T_126; // @[package.scala 100:49:@3613.4]
  reg  _T_129; // @[package.scala 48:56:@3614.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@3636.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@3638.4]
  reg  _T_153; // @[package.scala 48:56:@3639.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  wire  _T_158; // @[Controllers.scala 292:61:@3649.4]
  wire  _T_159; // @[Controllers.scala 292:24:@3650.4]
  SRFF active ( // @[Controllers.scala 261:22:@3547.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@3550.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_21 RetimeWrapper ( // @[package.scala 93:22:@3584.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_21 RetimeWrapper_1 ( // @[package.scala 93:22:@3606.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@3618.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@3626.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_4 ( // @[package.scala 93:22:@3642.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@3555.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@3556.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@3557.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@3558.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@3575.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@3589.4 package.scala 96:25:@3590.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@3591.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@3594.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@3599.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@3600.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@3603.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@3611.4 package.scala 96:25:@3612.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@3613.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@3638.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@3647.4 package.scala 96:25:@3648.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@3649.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@3650.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@3617.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@3652.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@3602.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@3605.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@3597.4]
  assign active_clock = clock; // @[:@3548.4]
  assign active_reset = reset; // @[:@3549.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@3560.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@3564.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@3565.4]
  assign done_clock = clock; // @[:@3551.4]
  assign done_reset = reset; // @[:@3552.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@3580.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@3573.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@3574.4]
  assign RetimeWrapper_clock = clock; // @[:@3585.4]
  assign RetimeWrapper_reset = reset; // @[:@3586.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@3588.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@3587.4]
  assign RetimeWrapper_1_clock = clock; // @[:@3607.4]
  assign RetimeWrapper_1_reset = reset; // @[:@3608.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@3610.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@3609.4]
  assign RetimeWrapper_2_clock = clock; // @[:@3619.4]
  assign RetimeWrapper_2_reset = reset; // @[:@3620.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@3622.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@3621.4]
  assign RetimeWrapper_3_clock = clock; // @[:@3627.4]
  assign RetimeWrapper_3_reset = reset; // @[:@3628.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@3630.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@3629.4]
  assign RetimeWrapper_4_clock = clock; // @[:@3643.4]
  assign RetimeWrapper_4_reset = reset; // @[:@3644.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@3646.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@3645.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module fix2fixBox( // @[:@3759.2]
  input  [31:0] io_a, // @[:@3762.4]
  output [31:0] io_b // @[:@3762.4]
);
  assign io_b = io_a; // @[Converter.scala 95:38:@3775.4]
endmodule
module _( // @[:@3777.2]
  input  [31:0] io_b, // @[:@3780.4]
  output [31:0] io_result // @[:@3780.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3785.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3785.4]
  fix2fixBox fix2fixBox ( // @[BigIPZynq.scala 219:30:@3785.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3793.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3788.4]
endmodule
module fix2fixBox_2( // @[:@3831.2]
  input  [31:0] io_a, // @[:@3834.4]
  output [32:0] io_b // @[:@3834.4]
);
  wire  _T_20; // @[implicits.scala 69:16:@3844.4]
  assign _T_20 = io_a[31]; // @[implicits.scala 69:16:@3844.4]
  assign io_b = {_T_20,io_a}; // @[Converter.scala 95:38:@3849.4]
endmodule
module __2( // @[:@3851.2]
  input  [31:0] io_b, // @[:@3854.4]
  output [32:0] io_result // @[:@3854.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@3859.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@3859.4]
  fix2fixBox_2 fix2fixBox ( // @[BigIPZynq.scala 219:30:@3859.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@3867.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@3862.4]
endmodule
module RetimeWrapper_29( // @[:@3919.2]
  input         clock, // @[:@3920.4]
  input         reset, // @[:@3921.4]
  input         io_flow, // @[:@3922.4]
  input  [31:0] io_in, // @[:@3922.4]
  output [31:0] io_out // @[:@3922.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@3924.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@3924.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@3937.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@3936.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@3935.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@3934.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@3933.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@3931.4]
endmodule
module fix2fixBox_4( // @[:@3939.2]
  input         clock, // @[:@3940.4]
  input         reset, // @[:@3941.4]
  input  [32:0] io_a, // @[:@3942.4]
  input         io_flow, // @[:@3942.4]
  output [31:0] io_b // @[:@3942.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@3955.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@3955.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@3955.4]
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@3955.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign io_b = RetimeWrapper_io_out; // @[Converter.scala 95:38:@3962.4]
  assign RetimeWrapper_clock = clock; // @[:@3956.4]
  assign RetimeWrapper_reset = reset; // @[:@3957.4]
  assign RetimeWrapper_io_flow = io_flow; // @[package.scala 95:18:@3959.4]
  assign RetimeWrapper_io_in = io_a[31:0]; // @[package.scala 94:16:@3958.4]
endmodule
module x452_sub( // @[:@3964.2]
  input         clock, // @[:@3965.4]
  input         reset, // @[:@3966.4]
  input  [31:0] io_a, // @[:@3967.4]
  input  [31:0] io_b, // @[:@3967.4]
  input         io_flow, // @[:@3967.4]
  output [31:0] io_result // @[:@3967.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@3975.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@3975.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@3982.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@3982.4]
  wire  fix2fixBox_clock; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_reset; // @[Math.scala 182:30:@4001.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 182:30:@4001.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 182:30:@4001.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 182:30:@4001.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  wire [33:0] _T_21; // @[Math.scala 177:37:@3989.4]
  wire [33:0] _T_22; // @[Math.scala 177:37:@3990.4]
  __2 _ ( // @[Math.scala 720:24:@3975.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@3982.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 182:30:@4001.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@3980.4 Math.scala 724:14:@3981.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@3987.4 Math.scala 724:14:@3988.4]
  assign _T_21 = a_upcast_number - b_upcast_number; // @[Math.scala 177:37:@3989.4]
  assign _T_22 = $unsigned(_T_21); // @[Math.scala 177:37:@3990.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 188:17:@4009.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@3978.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@3985.4]
  assign fix2fixBox_clock = clock; // @[:@4002.4]
  assign fix2fixBox_reset = reset; // @[:@4003.4]
  assign fix2fixBox_io_a = _T_22[32:0]; // @[Math.scala 183:23:@4004.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 186:26:@4007.4]
endmodule
module x235_sum( // @[:@4176.2]
  input         clock, // @[:@4177.4]
  input         reset, // @[:@4178.4]
  input  [31:0] io_a, // @[:@4179.4]
  input  [31:0] io_b, // @[:@4179.4]
  input         io_flow, // @[:@4179.4]
  output [31:0] io_result // @[:@4179.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@4187.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@4187.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@4194.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@4194.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@4212.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@4212.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@4212.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@4212.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@4201.4]
  __2 _ ( // @[Math.scala 720:24:@4187.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __2 __1 ( // @[Math.scala 720:24:@4194.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@4212.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@4192.4 Math.scala 724:14:@4193.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@4199.4 Math.scala 724:14:@4200.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@4201.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@4220.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@4190.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@4197.4]
  assign fix2fixBox_clock = clock; // @[:@4213.4]
  assign fix2fixBox_reset = reset; // @[:@4214.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@4215.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@4218.4]
endmodule
module x247_inr_Foreach_kernelx247_inr_Foreach_concrete1( // @[:@5106.2]
  input         clock, // @[:@5107.4]
  input         reset, // @[:@5108.4]
  output        io_in_x225_fifoinpacked_0_wPort_0_en_0, // @[:@5109.4]
  input         io_in_x225_fifoinpacked_0_full, // @[:@5109.4]
  output        io_in_x225_fifoinpacked_0_active_0_in, // @[:@5109.4]
  input         io_in_x225_fifoinpacked_0_active_0_out, // @[:@5109.4]
  input         io_sigsIn_backpressure, // @[:@5109.4]
  input         io_sigsIn_datapathEn, // @[:@5109.4]
  input         io_sigsIn_break, // @[:@5109.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_1, // @[:@5109.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@5109.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@5109.4]
  input         io_sigsIn_cchainOutputs_0_oobs_1, // @[:@5109.4]
  input         io_rr // @[:@5109.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@5143.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@5143.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@5155.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@5155.4]
  wire  x452_sub_1_clock; // @[Math.scala 191:24:@5182.4]
  wire  x452_sub_1_reset; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x452_sub_1_io_a; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x452_sub_1_io_b; // @[Math.scala 191:24:@5182.4]
  wire  x452_sub_1_io_flow; // @[Math.scala 191:24:@5182.4]
  wire [31:0] x452_sub_1_io_result; // @[Math.scala 191:24:@5182.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@5192.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@5192.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@5192.4]
  wire [31:0] RetimeWrapper_io_in; // @[package.scala 93:22:@5192.4]
  wire [31:0] RetimeWrapper_io_out; // @[package.scala 93:22:@5192.4]
  wire  x235_sum_1_clock; // @[Math.scala 150:24:@5201.4]
  wire  x235_sum_1_reset; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x235_sum_1_io_a; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x235_sum_1_io_b; // @[Math.scala 150:24:@5201.4]
  wire  x235_sum_1_io_flow; // @[Math.scala 150:24:@5201.4]
  wire [31:0] x235_sum_1_io_result; // @[Math.scala 150:24:@5201.4]
  wire  x236_sum_1_clock; // @[Math.scala 150:24:@5213.4]
  wire  x236_sum_1_reset; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x236_sum_1_io_a; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x236_sum_1_io_b; // @[Math.scala 150:24:@5213.4]
  wire  x236_sum_1_io_flow; // @[Math.scala 150:24:@5213.4]
  wire [31:0] x236_sum_1_io_result; // @[Math.scala 150:24:@5213.4]
  wire  x454_sum_1_clock; // @[Math.scala 150:24:@5228.4]
  wire  x454_sum_1_reset; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x454_sum_1_io_a; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x454_sum_1_io_b; // @[Math.scala 150:24:@5228.4]
  wire  x454_sum_1_io_flow; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x454_sum_1_io_result; // @[Math.scala 150:24:@5228.4]
  wire [31:0] x239_1_io_b; // @[Math.scala 720:24:@5249.4]
  wire [31:0] x239_1_io_result; // @[Math.scala 720:24:@5249.4]
  wire  x240_sum_1_clock; // @[Math.scala 150:24:@5260.4]
  wire  x240_sum_1_reset; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x240_sum_1_io_a; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x240_sum_1_io_b; // @[Math.scala 150:24:@5260.4]
  wire  x240_sum_1_io_flow; // @[Math.scala 150:24:@5260.4]
  wire [31:0] x240_sum_1_io_result; // @[Math.scala 150:24:@5260.4]
  wire  x457_sum_1_clock; // @[Math.scala 150:24:@5275.4]
  wire  x457_sum_1_reset; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x457_sum_1_io_a; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x457_sum_1_io_b; // @[Math.scala 150:24:@5275.4]
  wire  x457_sum_1_io_flow; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x457_sum_1_io_result; // @[Math.scala 150:24:@5275.4]
  wire [31:0] x243_1_io_b; // @[Math.scala 720:24:@5296.4]
  wire [31:0] x243_1_io_result; // @[Math.scala 720:24:@5296.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@5311.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@5320.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@5331.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@5331.4]
  wire  _T_327; // @[sm_x247_inr_Foreach.scala 62:18:@5168.4]
  wire  _T_328; // @[sm_x247_inr_Foreach.scala 62:55:@5169.4]
  wire [31:0] b230_number; // @[Math.scala 723:22:@5148.4 Math.scala 724:14:@5149.4]
  wire [42:0] _GEN_0; // @[Math.scala 461:32:@5173.4]
  wire [42:0] _T_331; // @[Math.scala 461:32:@5173.4]
  wire [38:0] _GEN_1; // @[Math.scala 461:32:@5178.4]
  wire [38:0] _T_334; // @[Math.scala 461:32:@5178.4]
  wire [31:0] x236_sum_number; // @[Math.scala 154:22:@5219.4 Math.scala 155:14:@5220.4]
  wire [33:0] _GEN_2; // @[Math.scala 461:32:@5224.4]
  wire [33:0] _T_353; // @[Math.scala 461:32:@5224.4]
  wire [31:0] x454_sum_number; // @[Math.scala 154:22:@5234.4 Math.scala 155:14:@5235.4]
  wire [31:0] _T_364; // @[Math.scala 406:49:@5241.4]
  wire [31:0] _T_366; // @[Math.scala 406:56:@5243.4]
  wire [31:0] _T_367; // @[Math.scala 406:56:@5244.4]
  wire [31:0] x240_sum_number; // @[Math.scala 154:22:@5266.4 Math.scala 155:14:@5267.4]
  wire [33:0] _GEN_3; // @[Math.scala 461:32:@5271.4]
  wire [33:0] _T_381; // @[Math.scala 461:32:@5271.4]
  wire [31:0] x457_sum_number; // @[Math.scala 154:22:@5281.4 Math.scala 155:14:@5282.4]
  wire [31:0] _T_392; // @[Math.scala 406:49:@5288.4]
  wire [31:0] _T_394; // @[Math.scala 406:56:@5290.4]
  wire [31:0] _T_395; // @[Math.scala 406:56:@5291.4]
  wire  _T_415; // @[sm_x247_inr_Foreach.scala 103:131:@5328.4]
  wire  _T_419; // @[package.scala 96:25:@5336.4 package.scala 96:25:@5337.4]
  wire  _T_421; // @[implicits.scala 55:10:@5338.4]
  wire  _T_422; // @[sm_x247_inr_Foreach.scala 103:148:@5339.4]
  wire  _T_424; // @[sm_x247_inr_Foreach.scala 103:236:@5341.4]
  wire  _T_425; // @[sm_x247_inr_Foreach.scala 103:255:@5342.4]
  wire  x481_b232_D4; // @[package.scala 96:25:@5316.4 package.scala 96:25:@5317.4]
  wire  _T_428; // @[sm_x247_inr_Foreach.scala 103:291:@5344.4]
  wire  x482_b233_D4; // @[package.scala 96:25:@5325.4 package.scala 96:25:@5326.4]
  _ _ ( // @[Math.scala 720:24:@5143.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@5155.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  x452_sub x452_sub_1 ( // @[Math.scala 191:24:@5182.4]
    .clock(x452_sub_1_clock),
    .reset(x452_sub_1_reset),
    .io_a(x452_sub_1_io_a),
    .io_b(x452_sub_1_io_b),
    .io_flow(x452_sub_1_io_flow),
    .io_result(x452_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper ( // @[package.scala 93:22:@5192.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x235_sum x235_sum_1 ( // @[Math.scala 150:24:@5201.4]
    .clock(x235_sum_1_clock),
    .reset(x235_sum_1_reset),
    .io_a(x235_sum_1_io_a),
    .io_b(x235_sum_1_io_b),
    .io_flow(x235_sum_1_io_flow),
    .io_result(x235_sum_1_io_result)
  );
  x235_sum x236_sum_1 ( // @[Math.scala 150:24:@5213.4]
    .clock(x236_sum_1_clock),
    .reset(x236_sum_1_reset),
    .io_a(x236_sum_1_io_a),
    .io_b(x236_sum_1_io_b),
    .io_flow(x236_sum_1_io_flow),
    .io_result(x236_sum_1_io_result)
  );
  x235_sum x454_sum_1 ( // @[Math.scala 150:24:@5228.4]
    .clock(x454_sum_1_clock),
    .reset(x454_sum_1_reset),
    .io_a(x454_sum_1_io_a),
    .io_b(x454_sum_1_io_b),
    .io_flow(x454_sum_1_io_flow),
    .io_result(x454_sum_1_io_result)
  );
  _ x239_1 ( // @[Math.scala 720:24:@5249.4]
    .io_b(x239_1_io_b),
    .io_result(x239_1_io_result)
  );
  x235_sum x240_sum_1 ( // @[Math.scala 150:24:@5260.4]
    .clock(x240_sum_1_clock),
    .reset(x240_sum_1_reset),
    .io_a(x240_sum_1_io_a),
    .io_b(x240_sum_1_io_b),
    .io_flow(x240_sum_1_io_flow),
    .io_result(x240_sum_1_io_result)
  );
  x235_sum x457_sum_1 ( // @[Math.scala 150:24:@5275.4]
    .clock(x457_sum_1_clock),
    .reset(x457_sum_1_reset),
    .io_a(x457_sum_1_io_a),
    .io_b(x457_sum_1_io_b),
    .io_flow(x457_sum_1_io_flow),
    .io_result(x457_sum_1_io_result)
  );
  _ x243_1 ( // @[Math.scala 720:24:@5296.4]
    .io_b(x243_1_io_b),
    .io_result(x243_1_io_result)
  );
  RetimeWrapper_25 RetimeWrapper_1 ( // @[package.scala 93:22:@5311.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_2 ( // @[package.scala 93:22:@5320.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_25 RetimeWrapper_3 ( // @[package.scala 93:22:@5331.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_327 = ~ io_in_x225_fifoinpacked_0_full; // @[sm_x247_inr_Foreach.scala 62:18:@5168.4]
  assign _T_328 = ~ io_in_x225_fifoinpacked_0_active_0_out; // @[sm_x247_inr_Foreach.scala 62:55:@5169.4]
  assign b230_number = __io_result; // @[Math.scala 723:22:@5148.4 Math.scala 724:14:@5149.4]
  assign _GEN_0 = {{11'd0}, b230_number}; // @[Math.scala 461:32:@5173.4]
  assign _T_331 = _GEN_0 << 11; // @[Math.scala 461:32:@5173.4]
  assign _GEN_1 = {{7'd0}, b230_number}; // @[Math.scala 461:32:@5178.4]
  assign _T_334 = _GEN_1 << 7; // @[Math.scala 461:32:@5178.4]
  assign x236_sum_number = x236_sum_1_io_result; // @[Math.scala 154:22:@5219.4 Math.scala 155:14:@5220.4]
  assign _GEN_2 = {{2'd0}, x236_sum_number}; // @[Math.scala 461:32:@5224.4]
  assign _T_353 = _GEN_2 << 2; // @[Math.scala 461:32:@5224.4]
  assign x454_sum_number = x454_sum_1_io_result; // @[Math.scala 154:22:@5234.4 Math.scala 155:14:@5235.4]
  assign _T_364 = $signed(x454_sum_number); // @[Math.scala 406:49:@5241.4]
  assign _T_366 = $signed(_T_364) & $signed(32'shff); // @[Math.scala 406:56:@5243.4]
  assign _T_367 = $signed(_T_366); // @[Math.scala 406:56:@5244.4]
  assign x240_sum_number = x240_sum_1_io_result; // @[Math.scala 154:22:@5266.4 Math.scala 155:14:@5267.4]
  assign _GEN_3 = {{2'd0}, x240_sum_number}; // @[Math.scala 461:32:@5271.4]
  assign _T_381 = _GEN_3 << 2; // @[Math.scala 461:32:@5271.4]
  assign x457_sum_number = x457_sum_1_io_result; // @[Math.scala 154:22:@5281.4 Math.scala 155:14:@5282.4]
  assign _T_392 = $signed(x457_sum_number); // @[Math.scala 406:49:@5288.4]
  assign _T_394 = $signed(_T_392) & $signed(32'shff); // @[Math.scala 406:56:@5290.4]
  assign _T_395 = $signed(_T_394); // @[Math.scala 406:56:@5291.4]
  assign _T_415 = ~ io_sigsIn_break; // @[sm_x247_inr_Foreach.scala 103:131:@5328.4]
  assign _T_419 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@5336.4 package.scala 96:25:@5337.4]
  assign _T_421 = io_rr ? _T_419 : 1'h0; // @[implicits.scala 55:10:@5338.4]
  assign _T_422 = _T_415 & _T_421; // @[sm_x247_inr_Foreach.scala 103:148:@5339.4]
  assign _T_424 = _T_422 & _T_415; // @[sm_x247_inr_Foreach.scala 103:236:@5341.4]
  assign _T_425 = _T_424 & io_sigsIn_backpressure; // @[sm_x247_inr_Foreach.scala 103:255:@5342.4]
  assign x481_b232_D4 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@5316.4 package.scala 96:25:@5317.4]
  assign _T_428 = _T_425 & x481_b232_D4; // @[sm_x247_inr_Foreach.scala 103:291:@5344.4]
  assign x482_b233_D4 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@5325.4 package.scala 96:25:@5326.4]
  assign io_in_x225_fifoinpacked_0_wPort_0_en_0 = _T_428 & x482_b233_D4; // @[MemInterfaceType.scala 93:57:@5348.4]
  assign io_in_x225_fifoinpacked_0_active_0_in = x481_b232_D4 & x482_b233_D4; // @[MemInterfaceType.scala 147:18:@5351.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@5146.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@5158.4]
  assign x452_sub_1_clock = clock; // @[:@5183.4]
  assign x452_sub_1_reset = reset; // @[:@5184.4]
  assign x452_sub_1_io_a = _T_331[31:0]; // @[Math.scala 192:17:@5185.4]
  assign x452_sub_1_io_b = _T_334[31:0]; // @[Math.scala 193:17:@5186.4]
  assign x452_sub_1_io_flow = _T_327 | _T_328; // @[Math.scala 194:20:@5187.4]
  assign RetimeWrapper_clock = clock; // @[:@5193.4]
  assign RetimeWrapper_reset = reset; // @[:@5194.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5196.4]
  assign RetimeWrapper_io_in = __1_io_result; // @[package.scala 94:16:@5195.4]
  assign x235_sum_1_clock = clock; // @[:@5202.4]
  assign x235_sum_1_reset = reset; // @[:@5203.4]
  assign x235_sum_1_io_a = x452_sub_1_io_result; // @[Math.scala 151:17:@5204.4]
  assign x235_sum_1_io_b = RetimeWrapper_io_out; // @[Math.scala 152:17:@5205.4]
  assign x235_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5206.4]
  assign x236_sum_1_clock = clock; // @[:@5214.4]
  assign x236_sum_1_reset = reset; // @[:@5215.4]
  assign x236_sum_1_io_a = x235_sum_1_io_result; // @[Math.scala 151:17:@5216.4]
  assign x236_sum_1_io_b = 32'h1; // @[Math.scala 152:17:@5217.4]
  assign x236_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5218.4]
  assign x454_sum_1_clock = clock; // @[:@5229.4]
  assign x454_sum_1_reset = reset; // @[:@5230.4]
  assign x454_sum_1_io_a = _T_353[31:0]; // @[Math.scala 151:17:@5231.4]
  assign x454_sum_1_io_b = x236_sum_1_io_result; // @[Math.scala 152:17:@5232.4]
  assign x454_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5233.4]
  assign x239_1_io_b = $unsigned(_T_367); // @[Math.scala 721:17:@5252.4]
  assign x240_sum_1_clock = clock; // @[:@5261.4]
  assign x240_sum_1_reset = reset; // @[:@5262.4]
  assign x240_sum_1_io_a = x235_sum_1_io_result; // @[Math.scala 151:17:@5263.4]
  assign x240_sum_1_io_b = 32'h2; // @[Math.scala 152:17:@5264.4]
  assign x240_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5265.4]
  assign x457_sum_1_clock = clock; // @[:@5276.4]
  assign x457_sum_1_reset = reset; // @[:@5277.4]
  assign x457_sum_1_io_a = _T_381[31:0]; // @[Math.scala 151:17:@5278.4]
  assign x457_sum_1_io_b = x240_sum_1_io_result; // @[Math.scala 152:17:@5279.4]
  assign x457_sum_1_io_flow = _T_327 | _T_328; // @[Math.scala 153:20:@5280.4]
  assign x243_1_io_b = $unsigned(_T_395); // @[Math.scala 721:17:@5299.4]
  assign RetimeWrapper_1_clock = clock; // @[:@5312.4]
  assign RetimeWrapper_1_reset = reset; // @[:@5313.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5315.4]
  assign RetimeWrapper_1_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@5314.4]
  assign RetimeWrapper_2_clock = clock; // @[:@5321.4]
  assign RetimeWrapper_2_reset = reset; // @[:@5322.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5324.4]
  assign RetimeWrapper_2_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@5323.4]
  assign RetimeWrapper_3_clock = clock; // @[:@5332.4]
  assign RetimeWrapper_3_reset = reset; // @[:@5333.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@5335.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@5334.4]
endmodule
module RetimeWrapper_44( // @[:@6469.2]
  input   clock, // @[:@6470.4]
  input   reset, // @[:@6471.4]
  input   io_flow, // @[:@6472.4]
  input   io_in, // @[:@6472.4]
  output  io_out // @[:@6472.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6474.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(31)) sr ( // @[RetimeShiftRegister.scala 15:20:@6474.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6487.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6486.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6485.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6484.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6483.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6481.4]
endmodule
module RetimeWrapper_48( // @[:@6597.2]
  input   clock, // @[:@6598.4]
  input   reset, // @[:@6599.4]
  input   io_flow, // @[:@6600.4]
  input   io_in, // @[:@6600.4]
  output  io_out // @[:@6600.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6602.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(30)) sr ( // @[RetimeShiftRegister.scala 15:20:@6602.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6615.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6614.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@6613.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6612.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6611.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6609.4]
endmodule
module x401_inr_Foreach_SAMPLER_BOX_sm( // @[:@6617.2]
  input   clock, // @[:@6618.4]
  input   reset, // @[:@6619.4]
  input   io_enable, // @[:@6620.4]
  output  io_done, // @[:@6620.4]
  output  io_doneLatch, // @[:@6620.4]
  input   io_ctrDone, // @[:@6620.4]
  output  io_datapathEn, // @[:@6620.4]
  output  io_ctrInc, // @[:@6620.4]
  output  io_ctrRst, // @[:@6620.4]
  input   io_parentAck, // @[:@6620.4]
  input   io_backpressure, // @[:@6620.4]
  input   io_break // @[:@6620.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@6622.4]
  wire  active_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@6622.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@6622.4]
  wire  done_clock; // @[Controllers.scala 262:20:@6625.4]
  wire  done_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@6625.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@6625.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@6659.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@6681.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@6693.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@6701.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@6717.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@6717.4]
  wire  _T_80; // @[Controllers.scala 264:48:@6630.4]
  wire  _T_81; // @[Controllers.scala 264:46:@6631.4]
  wire  _T_82; // @[Controllers.scala 264:62:@6632.4]
  wire  _T_83; // @[Controllers.scala 264:60:@6633.4]
  wire  _T_100; // @[package.scala 100:49:@6650.4]
  reg  _T_103; // @[package.scala 48:56:@6651.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@6664.4 package.scala 96:25:@6665.4]
  wire  _T_110; // @[package.scala 100:49:@6666.4]
  reg  _T_113; // @[package.scala 48:56:@6667.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@6669.4]
  wire  _T_118; // @[Controllers.scala 283:41:@6674.4]
  wire  _T_119; // @[Controllers.scala 283:59:@6675.4]
  wire  _T_121; // @[Controllers.scala 284:37:@6678.4]
  wire  _T_124; // @[package.scala 96:25:@6686.4 package.scala 96:25:@6687.4]
  wire  _T_126; // @[package.scala 100:49:@6688.4]
  reg  _T_129; // @[package.scala 48:56:@6689.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@6711.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@6713.4]
  reg  _T_153; // @[package.scala 48:56:@6714.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@6722.4 package.scala 96:25:@6723.4]
  wire  _T_158; // @[Controllers.scala 292:61:@6724.4]
  wire  _T_159; // @[Controllers.scala 292:24:@6725.4]
  SRFF active ( // @[Controllers.scala 261:22:@6622.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@6625.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_44 RetimeWrapper ( // @[package.scala 93:22:@6659.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_44 RetimeWrapper_1 ( // @[package.scala 93:22:@6681.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@6693.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@6701.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_4 ( // @[package.scala 93:22:@6717.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@6630.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@6631.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@6632.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@6633.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@6650.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@6664.4 package.scala 96:25:@6665.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@6666.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@6669.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@6674.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@6675.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@6678.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@6686.4 package.scala 96:25:@6687.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@6688.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@6713.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@6722.4 package.scala 96:25:@6723.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@6724.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@6725.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@6692.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@6727.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@6677.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@6680.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@6672.4]
  assign active_clock = clock; // @[:@6623.4]
  assign active_reset = reset; // @[:@6624.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@6635.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@6639.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@6640.4]
  assign done_clock = clock; // @[:@6626.4]
  assign done_reset = reset; // @[:@6627.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@6655.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@6648.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@6649.4]
  assign RetimeWrapper_clock = clock; // @[:@6660.4]
  assign RetimeWrapper_reset = reset; // @[:@6661.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@6663.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@6662.4]
  assign RetimeWrapper_1_clock = clock; // @[:@6682.4]
  assign RetimeWrapper_1_reset = reset; // @[:@6683.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@6685.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@6684.4]
  assign RetimeWrapper_2_clock = clock; // @[:@6694.4]
  assign RetimeWrapper_2_reset = reset; // @[:@6695.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@6697.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@6696.4]
  assign RetimeWrapper_3_clock = clock; // @[:@6702.4]
  assign RetimeWrapper_3_reset = reset; // @[:@6703.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@6705.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@6704.4]
  assign RetimeWrapper_4_clock = clock; // @[:@6718.4]
  assign RetimeWrapper_4_reset = reset; // @[:@6719.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@6721.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@6720.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module RetimeWrapper_52( // @[:@6918.2]
  input         clock, // @[:@6919.4]
  input         reset, // @[:@6920.4]
  input         io_flow, // @[:@6921.4]
  input  [63:0] io_in, // @[:@6921.4]
  output [63:0] io_out // @[:@6921.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@6923.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@6923.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@6936.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@6935.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@6934.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@6933.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@6932.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@6930.4]
endmodule
module SRAM_1( // @[:@6954.2]
  input         clock, // @[:@6955.4]
  input         reset, // @[:@6956.4]
  input  [8:0]  io_raddr, // @[:@6957.4]
  input         io_wen, // @[:@6957.4]
  input  [8:0]  io_waddr, // @[:@6957.4]
  input  [31:0] io_wdata, // @[:@6957.4]
  output [31:0] io_rdata, // @[:@6957.4]
  input         io_backpressure // @[:@6957.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@6959.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@6959.4]
  wire [8:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@6959.4]
  wire [8:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@6959.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@6959.4]
  wire  _T_19; // @[SRAM.scala 182:49:@6977.4]
  wire  _T_20; // @[SRAM.scala 182:37:@6978.4]
  reg  _T_23; // @[SRAM.scala 182:29:@6979.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@6981.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(480), .AWIDTH(9)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@6959.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@6977.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@6978.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@6986.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@6973.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@6974.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@6971.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@6976.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@6975.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@6972.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@6970.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@6969.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module RetimeWrapper_53( // @[:@7000.2]
  input        clock, // @[:@7001.4]
  input        reset, // @[:@7002.4]
  input        io_flow, // @[:@7003.4]
  input  [8:0] io_in, // @[:@7003.4]
  output [8:0] io_out // @[:@7003.4]
);
  wire [8:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire [8:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire [8:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@7005.4]
  RetimeShiftRegister #(.WIDTH(9), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@7005.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@7018.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@7017.4]
  assign sr_init = 9'h0; // @[RetimeShiftRegister.scala 19:16:@7016.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@7015.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@7014.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@7012.4]
endmodule
module Mem1D_5( // @[:@7020.2]
  input         clock, // @[:@7021.4]
  input         reset, // @[:@7022.4]
  input  [8:0]  io_r_ofs_0, // @[:@7023.4]
  input         io_r_backpressure, // @[:@7023.4]
  input  [8:0]  io_w_ofs_0, // @[:@7023.4]
  input  [31:0] io_w_data_0, // @[:@7023.4]
  input         io_w_en_0, // @[:@7023.4]
  output [31:0] io_output // @[:@7023.4]
);
  wire  SRAM_clock; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_reset; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [8:0] SRAM_io_raddr; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_io_wen; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [8:0] SRAM_io_waddr; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [31:0] SRAM_io_wdata; // @[MemPrimitives.scala 715:21:@7027.4]
  wire [31:0] SRAM_io_rdata; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  SRAM_io_backpressure; // @[MemPrimitives.scala 715:21:@7027.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@7030.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@7030.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@7030.4]
  wire [8:0] RetimeWrapper_io_in; // @[package.scala 93:22:@7030.4]
  wire [8:0] RetimeWrapper_io_out; // @[package.scala 93:22:@7030.4]
  wire  wInBound; // @[MemPrimitives.scala 702:32:@7025.4]
  SRAM_1 SRAM ( // @[MemPrimitives.scala 715:21:@7027.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  RetimeWrapper_53 RetimeWrapper ( // @[package.scala 93:22:@7030.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign wInBound = io_w_ofs_0 <= 9'h1e0; // @[MemPrimitives.scala 702:32:@7025.4]
  assign io_output = SRAM_io_rdata; // @[MemPrimitives.scala 722:17:@7043.4]
  assign SRAM_clock = clock; // @[:@7028.4]
  assign SRAM_reset = reset; // @[:@7029.4]
  assign SRAM_io_raddr = RetimeWrapper_io_out; // @[MemPrimitives.scala 716:37:@7037.4]
  assign SRAM_io_wen = io_w_en_0 & wInBound; // @[MemPrimitives.scala 719:22:@7040.4]
  assign SRAM_io_waddr = io_w_ofs_0; // @[MemPrimitives.scala 718:22:@7038.4]
  assign SRAM_io_wdata = io_w_data_0; // @[MemPrimitives.scala 720:22:@7041.4]
  assign SRAM_io_backpressure = io_r_backpressure; // @[MemPrimitives.scala 721:30:@7042.4]
  assign RetimeWrapper_clock = clock; // @[:@7031.4]
  assign RetimeWrapper_reset = reset; // @[:@7032.4]
  assign RetimeWrapper_io_flow = io_r_backpressure; // @[package.scala 95:18:@7034.4]
  assign RetimeWrapper_io_in = io_r_ofs_0; // @[package.scala 94:16:@7033.4]
endmodule
module StickySelects_1( // @[:@8650.2]
  input   clock, // @[:@8651.4]
  input   reset, // @[:@8652.4]
  input   io_ins_0, // @[:@8653.4]
  input   io_ins_1, // @[:@8653.4]
  input   io_ins_2, // @[:@8653.4]
  input   io_ins_3, // @[:@8653.4]
  input   io_ins_4, // @[:@8653.4]
  input   io_ins_5, // @[:@8653.4]
  output  io_outs_0, // @[:@8653.4]
  output  io_outs_1, // @[:@8653.4]
  output  io_outs_2, // @[:@8653.4]
  output  io_outs_3, // @[:@8653.4]
  output  io_outs_4, // @[:@8653.4]
  output  io_outs_5 // @[:@8653.4]
);
  reg  _T_19; // @[StickySelects.scala 37:46:@8655.4]
  reg [31:0] _RAND_0;
  reg  _T_22; // @[StickySelects.scala 37:46:@8656.4]
  reg [31:0] _RAND_1;
  reg  _T_25; // @[StickySelects.scala 37:46:@8657.4]
  reg [31:0] _RAND_2;
  reg  _T_28; // @[StickySelects.scala 37:46:@8658.4]
  reg [31:0] _RAND_3;
  reg  _T_31; // @[StickySelects.scala 37:46:@8659.4]
  reg [31:0] _RAND_4;
  reg  _T_34; // @[StickySelects.scala 37:46:@8660.4]
  reg [31:0] _RAND_5;
  wire  _T_35; // @[StickySelects.scala 47:46:@8661.4]
  wire  _T_36; // @[StickySelects.scala 47:46:@8662.4]
  wire  _T_37; // @[StickySelects.scala 47:46:@8663.4]
  wire  _T_38; // @[StickySelects.scala 47:46:@8664.4]
  wire  _T_39; // @[StickySelects.scala 49:53:@8665.4]
  wire  _T_40; // @[StickySelects.scala 49:21:@8666.4]
  wire  _T_41; // @[StickySelects.scala 47:46:@8668.4]
  wire  _T_42; // @[StickySelects.scala 47:46:@8669.4]
  wire  _T_43; // @[StickySelects.scala 47:46:@8670.4]
  wire  _T_44; // @[StickySelects.scala 47:46:@8671.4]
  wire  _T_45; // @[StickySelects.scala 49:53:@8672.4]
  wire  _T_46; // @[StickySelects.scala 49:21:@8673.4]
  wire  _T_47; // @[StickySelects.scala 47:46:@8675.4]
  wire  _T_48; // @[StickySelects.scala 47:46:@8676.4]
  wire  _T_49; // @[StickySelects.scala 47:46:@8677.4]
  wire  _T_50; // @[StickySelects.scala 47:46:@8678.4]
  wire  _T_51; // @[StickySelects.scala 49:53:@8679.4]
  wire  _T_52; // @[StickySelects.scala 49:21:@8680.4]
  wire  _T_54; // @[StickySelects.scala 47:46:@8683.4]
  wire  _T_55; // @[StickySelects.scala 47:46:@8684.4]
  wire  _T_56; // @[StickySelects.scala 47:46:@8685.4]
  wire  _T_57; // @[StickySelects.scala 49:53:@8686.4]
  wire  _T_58; // @[StickySelects.scala 49:21:@8687.4]
  wire  _T_61; // @[StickySelects.scala 47:46:@8691.4]
  wire  _T_62; // @[StickySelects.scala 47:46:@8692.4]
  wire  _T_63; // @[StickySelects.scala 49:53:@8693.4]
  wire  _T_64; // @[StickySelects.scala 49:21:@8694.4]
  wire  _T_68; // @[StickySelects.scala 47:46:@8699.4]
  wire  _T_69; // @[StickySelects.scala 49:53:@8700.4]
  wire  _T_70; // @[StickySelects.scala 49:21:@8701.4]
  assign _T_35 = io_ins_1 | io_ins_2; // @[StickySelects.scala 47:46:@8661.4]
  assign _T_36 = _T_35 | io_ins_3; // @[StickySelects.scala 47:46:@8662.4]
  assign _T_37 = _T_36 | io_ins_4; // @[StickySelects.scala 47:46:@8663.4]
  assign _T_38 = _T_37 | io_ins_5; // @[StickySelects.scala 47:46:@8664.4]
  assign _T_39 = io_ins_0 | _T_19; // @[StickySelects.scala 49:53:@8665.4]
  assign _T_40 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 49:21:@8666.4]
  assign _T_41 = io_ins_0 | io_ins_2; // @[StickySelects.scala 47:46:@8668.4]
  assign _T_42 = _T_41 | io_ins_3; // @[StickySelects.scala 47:46:@8669.4]
  assign _T_43 = _T_42 | io_ins_4; // @[StickySelects.scala 47:46:@8670.4]
  assign _T_44 = _T_43 | io_ins_5; // @[StickySelects.scala 47:46:@8671.4]
  assign _T_45 = io_ins_1 | _T_22; // @[StickySelects.scala 49:53:@8672.4]
  assign _T_46 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 49:21:@8673.4]
  assign _T_47 = io_ins_0 | io_ins_1; // @[StickySelects.scala 47:46:@8675.4]
  assign _T_48 = _T_47 | io_ins_3; // @[StickySelects.scala 47:46:@8676.4]
  assign _T_49 = _T_48 | io_ins_4; // @[StickySelects.scala 47:46:@8677.4]
  assign _T_50 = _T_49 | io_ins_5; // @[StickySelects.scala 47:46:@8678.4]
  assign _T_51 = io_ins_2 | _T_25; // @[StickySelects.scala 49:53:@8679.4]
  assign _T_52 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 49:21:@8680.4]
  assign _T_54 = _T_47 | io_ins_2; // @[StickySelects.scala 47:46:@8683.4]
  assign _T_55 = _T_54 | io_ins_4; // @[StickySelects.scala 47:46:@8684.4]
  assign _T_56 = _T_55 | io_ins_5; // @[StickySelects.scala 47:46:@8685.4]
  assign _T_57 = io_ins_3 | _T_28; // @[StickySelects.scala 49:53:@8686.4]
  assign _T_58 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 49:21:@8687.4]
  assign _T_61 = _T_54 | io_ins_3; // @[StickySelects.scala 47:46:@8691.4]
  assign _T_62 = _T_61 | io_ins_5; // @[StickySelects.scala 47:46:@8692.4]
  assign _T_63 = io_ins_4 | _T_31; // @[StickySelects.scala 49:53:@8693.4]
  assign _T_64 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 49:21:@8694.4]
  assign _T_68 = _T_61 | io_ins_4; // @[StickySelects.scala 47:46:@8699.4]
  assign _T_69 = io_ins_5 | _T_34; // @[StickySelects.scala 49:53:@8700.4]
  assign _T_70 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 49:21:@8701.4]
  assign io_outs_0 = _T_38 ? io_ins_0 : _T_39; // @[StickySelects.scala 53:57:@8703.4]
  assign io_outs_1 = _T_44 ? io_ins_1 : _T_45; // @[StickySelects.scala 53:57:@8704.4]
  assign io_outs_2 = _T_50 ? io_ins_2 : _T_51; // @[StickySelects.scala 53:57:@8705.4]
  assign io_outs_3 = _T_56 ? io_ins_3 : _T_57; // @[StickySelects.scala 53:57:@8706.4]
  assign io_outs_4 = _T_62 ? io_ins_4 : _T_63; // @[StickySelects.scala 53:57:@8707.4]
  assign io_outs_5 = _T_68 ? io_ins_5 : _T_69; // @[StickySelects.scala 53:57:@8708.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_19 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_22 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_25 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_28 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_31 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_19 <= 1'h0;
    end else begin
      if (_T_38) begin
        _T_19 <= io_ins_0;
      end else begin
        _T_19 <= _T_39;
      end
    end
    if (reset) begin
      _T_22 <= 1'h0;
    end else begin
      if (_T_44) begin
        _T_22 <= io_ins_1;
      end else begin
        _T_22 <= _T_45;
      end
    end
    if (reset) begin
      _T_25 <= 1'h0;
    end else begin
      if (_T_50) begin
        _T_25 <= io_ins_2;
      end else begin
        _T_25 <= _T_51;
      end
    end
    if (reset) begin
      _T_28 <= 1'h0;
    end else begin
      if (_T_56) begin
        _T_28 <= io_ins_3;
      end else begin
        _T_28 <= _T_57;
      end
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else begin
      if (_T_62) begin
        _T_31 <= io_ins_4;
      end else begin
        _T_31 <= _T_63;
      end
    end
    if (reset) begin
      _T_34 <= 1'h0;
    end else begin
      if (_T_68) begin
        _T_34 <= io_ins_5;
      end else begin
        _T_34 <= _T_69;
      end
    end
  end
endmodule
module x258_lb_0( // @[:@12682.2]
  input         clock, // @[:@12683.4]
  input         reset, // @[:@12684.4]
  input  [2:0]  io_rPort_11_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_11_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_11_ofs_0, // @[:@12685.4]
  input         io_rPort_11_en_0, // @[:@12685.4]
  input         io_rPort_11_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_11_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_10_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_10_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_10_ofs_0, // @[:@12685.4]
  input         io_rPort_10_en_0, // @[:@12685.4]
  input         io_rPort_10_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_10_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_9_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_9_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_9_ofs_0, // @[:@12685.4]
  input         io_rPort_9_en_0, // @[:@12685.4]
  input         io_rPort_9_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_9_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_8_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_8_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_8_ofs_0, // @[:@12685.4]
  input         io_rPort_8_en_0, // @[:@12685.4]
  input         io_rPort_8_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_8_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_7_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_7_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_7_ofs_0, // @[:@12685.4]
  input         io_rPort_7_en_0, // @[:@12685.4]
  input         io_rPort_7_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_7_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_6_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_6_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_6_ofs_0, // @[:@12685.4]
  input         io_rPort_6_en_0, // @[:@12685.4]
  input         io_rPort_6_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_6_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_5_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_5_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_5_ofs_0, // @[:@12685.4]
  input         io_rPort_5_en_0, // @[:@12685.4]
  input         io_rPort_5_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_5_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_4_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_4_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_4_ofs_0, // @[:@12685.4]
  input         io_rPort_4_en_0, // @[:@12685.4]
  input         io_rPort_4_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_4_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_3_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_3_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_3_ofs_0, // @[:@12685.4]
  input         io_rPort_3_en_0, // @[:@12685.4]
  input         io_rPort_3_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_3_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_2_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_2_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_2_ofs_0, // @[:@12685.4]
  input         io_rPort_2_en_0, // @[:@12685.4]
  input         io_rPort_2_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_2_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_1_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_1_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_1_ofs_0, // @[:@12685.4]
  input         io_rPort_1_en_0, // @[:@12685.4]
  input         io_rPort_1_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_1_output_0, // @[:@12685.4]
  input  [2:0]  io_rPort_0_banks_1, // @[:@12685.4]
  input  [2:0]  io_rPort_0_banks_0, // @[:@12685.4]
  input  [8:0]  io_rPort_0_ofs_0, // @[:@12685.4]
  input         io_rPort_0_en_0, // @[:@12685.4]
  input         io_rPort_0_backpressure, // @[:@12685.4]
  output [31:0] io_rPort_0_output_0, // @[:@12685.4]
  input  [2:0]  io_wPort_1_banks_1, // @[:@12685.4]
  input  [2:0]  io_wPort_1_banks_0, // @[:@12685.4]
  input  [8:0]  io_wPort_1_ofs_0, // @[:@12685.4]
  input  [31:0] io_wPort_1_data_0, // @[:@12685.4]
  input         io_wPort_1_en_0, // @[:@12685.4]
  input  [2:0]  io_wPort_0_banks_1, // @[:@12685.4]
  input  [2:0]  io_wPort_0_banks_0, // @[:@12685.4]
  input  [8:0]  io_wPort_0_ofs_0, // @[:@12685.4]
  input  [31:0] io_wPort_0_data_0, // @[:@12685.4]
  input         io_wPort_0_en_0 // @[:@12685.4]
);
  wire  Mem1D_clock; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_reset; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [8:0] Mem1D_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [8:0] Mem1D_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [31:0] Mem1D_io_w_data_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_io_w_en_0; // @[MemPrimitives.scala 64:21:@12776.4]
  wire [31:0] Mem1D_io_output; // @[MemPrimitives.scala 64:21:@12776.4]
  wire  Mem1D_1_clock; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_reset; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [8:0] Mem1D_1_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [8:0] Mem1D_1_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [31:0] Mem1D_1_io_w_data_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_1_io_w_en_0; // @[MemPrimitives.scala 64:21:@12792.4]
  wire [31:0] Mem1D_1_io_output; // @[MemPrimitives.scala 64:21:@12792.4]
  wire  Mem1D_2_clock; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_reset; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [8:0] Mem1D_2_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [8:0] Mem1D_2_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [31:0] Mem1D_2_io_w_data_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_2_io_w_en_0; // @[MemPrimitives.scala 64:21:@12808.4]
  wire [31:0] Mem1D_2_io_output; // @[MemPrimitives.scala 64:21:@12808.4]
  wire  Mem1D_3_clock; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_reset; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [8:0] Mem1D_3_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [8:0] Mem1D_3_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [31:0] Mem1D_3_io_w_data_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_3_io_w_en_0; // @[MemPrimitives.scala 64:21:@12824.4]
  wire [31:0] Mem1D_3_io_output; // @[MemPrimitives.scala 64:21:@12824.4]
  wire  Mem1D_4_clock; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_reset; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [8:0] Mem1D_4_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [8:0] Mem1D_4_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [31:0] Mem1D_4_io_w_data_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_4_io_w_en_0; // @[MemPrimitives.scala 64:21:@12840.4]
  wire [31:0] Mem1D_4_io_output; // @[MemPrimitives.scala 64:21:@12840.4]
  wire  Mem1D_5_clock; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_reset; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [8:0] Mem1D_5_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [8:0] Mem1D_5_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [31:0] Mem1D_5_io_w_data_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_5_io_w_en_0; // @[MemPrimitives.scala 64:21:@12856.4]
  wire [31:0] Mem1D_5_io_output; // @[MemPrimitives.scala 64:21:@12856.4]
  wire  Mem1D_6_clock; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_reset; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [8:0] Mem1D_6_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [8:0] Mem1D_6_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [31:0] Mem1D_6_io_w_data_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_6_io_w_en_0; // @[MemPrimitives.scala 64:21:@12872.4]
  wire [31:0] Mem1D_6_io_output; // @[MemPrimitives.scala 64:21:@12872.4]
  wire  Mem1D_7_clock; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_reset; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [8:0] Mem1D_7_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [8:0] Mem1D_7_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [31:0] Mem1D_7_io_w_data_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_7_io_w_en_0; // @[MemPrimitives.scala 64:21:@12888.4]
  wire [31:0] Mem1D_7_io_output; // @[MemPrimitives.scala 64:21:@12888.4]
  wire  Mem1D_8_clock; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_reset; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [8:0] Mem1D_8_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [8:0] Mem1D_8_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [31:0] Mem1D_8_io_w_data_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_8_io_w_en_0; // @[MemPrimitives.scala 64:21:@12904.4]
  wire [31:0] Mem1D_8_io_output; // @[MemPrimitives.scala 64:21:@12904.4]
  wire  Mem1D_9_clock; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_reset; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [8:0] Mem1D_9_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [8:0] Mem1D_9_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [31:0] Mem1D_9_io_w_data_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_9_io_w_en_0; // @[MemPrimitives.scala 64:21:@12920.4]
  wire [31:0] Mem1D_9_io_output; // @[MemPrimitives.scala 64:21:@12920.4]
  wire  Mem1D_10_clock; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_reset; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [8:0] Mem1D_10_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [8:0] Mem1D_10_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [31:0] Mem1D_10_io_w_data_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_10_io_w_en_0; // @[MemPrimitives.scala 64:21:@12936.4]
  wire [31:0] Mem1D_10_io_output; // @[MemPrimitives.scala 64:21:@12936.4]
  wire  Mem1D_11_clock; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_reset; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [8:0] Mem1D_11_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [8:0] Mem1D_11_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [31:0] Mem1D_11_io_w_data_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_11_io_w_en_0; // @[MemPrimitives.scala 64:21:@12952.4]
  wire [31:0] Mem1D_11_io_output; // @[MemPrimitives.scala 64:21:@12952.4]
  wire  Mem1D_12_clock; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_reset; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [8:0] Mem1D_12_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [8:0] Mem1D_12_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [31:0] Mem1D_12_io_w_data_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_12_io_w_en_0; // @[MemPrimitives.scala 64:21:@12968.4]
  wire [31:0] Mem1D_12_io_output; // @[MemPrimitives.scala 64:21:@12968.4]
  wire  Mem1D_13_clock; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_reset; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [8:0] Mem1D_13_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_io_r_backpressure; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [8:0] Mem1D_13_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [31:0] Mem1D_13_io_w_data_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_13_io_w_en_0; // @[MemPrimitives.scala 64:21:@12984.4]
  wire [31:0] Mem1D_13_io_output; // @[MemPrimitives.scala 64:21:@12984.4]
  wire  Mem1D_14_clock; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_reset; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [8:0] Mem1D_14_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [8:0] Mem1D_14_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [31:0] Mem1D_14_io_w_data_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_14_io_w_en_0; // @[MemPrimitives.scala 64:21:@13000.4]
  wire [31:0] Mem1D_14_io_output; // @[MemPrimitives.scala 64:21:@13000.4]
  wire  Mem1D_15_clock; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_reset; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [8:0] Mem1D_15_io_r_ofs_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_io_r_backpressure; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [8:0] Mem1D_15_io_w_ofs_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [31:0] Mem1D_15_io_w_data_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  Mem1D_15_io_w_en_0; // @[MemPrimitives.scala 64:21:@13016.4]
  wire [31:0] Mem1D_15_io_output; // @[MemPrimitives.scala 64:21:@13016.4]
  wire  StickySelects_clock; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_reset; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_0; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_1; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_2; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_3; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_4; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_ins_5; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_0; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_1; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_2; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_3; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_4; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_io_outs_5; // @[MemPrimitives.scala 124:33:@13248.4]
  wire  StickySelects_1_clock; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_reset; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_ins_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_0; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_1; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_2; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_3; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_4; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_1_io_outs_5; // @[MemPrimitives.scala 124:33:@13310.4]
  wire  StickySelects_2_clock; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_reset; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_0; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_1; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_2; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_3; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_4; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_ins_5; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_0; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_1; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_2; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_3; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_4; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_2_io_outs_5; // @[MemPrimitives.scala 124:33:@13372.4]
  wire  StickySelects_3_clock; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_reset; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_0; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_1; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_2; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_3; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_4; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_ins_5; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_0; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_1; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_2; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_3; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_4; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_3_io_outs_5; // @[MemPrimitives.scala 124:33:@13434.4]
  wire  StickySelects_4_clock; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_reset; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_0; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_1; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_2; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_3; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_4; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_ins_5; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_0; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_1; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_2; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_3; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_4; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_4_io_outs_5; // @[MemPrimitives.scala 124:33:@13496.4]
  wire  StickySelects_5_clock; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_reset; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_0; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_1; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_2; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_3; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_4; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_ins_5; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_0; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_1; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_2; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_3; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_4; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_5_io_outs_5; // @[MemPrimitives.scala 124:33:@13558.4]
  wire  StickySelects_6_clock; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_reset; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_0; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_1; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_2; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_3; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_4; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_ins_5; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_0; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_1; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_2; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_3; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_4; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_6_io_outs_5; // @[MemPrimitives.scala 124:33:@13620.4]
  wire  StickySelects_7_clock; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_reset; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_0; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_1; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_2; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_3; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_4; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_ins_5; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_0; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_1; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_2; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_3; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_4; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_7_io_outs_5; // @[MemPrimitives.scala 124:33:@13682.4]
  wire  StickySelects_8_clock; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_reset; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_0; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_1; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_2; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_3; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_4; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_ins_5; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_0; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_1; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_2; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_3; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_4; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_8_io_outs_5; // @[MemPrimitives.scala 124:33:@13744.4]
  wire  StickySelects_9_clock; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_reset; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_0; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_1; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_2; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_3; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_4; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_ins_5; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_0; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_1; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_2; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_3; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_4; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_9_io_outs_5; // @[MemPrimitives.scala 124:33:@13806.4]
  wire  StickySelects_10_clock; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_reset; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_0; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_1; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_2; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_3; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_4; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_ins_5; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_0; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_1; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_2; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_3; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_4; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_10_io_outs_5; // @[MemPrimitives.scala 124:33:@13868.4]
  wire  StickySelects_11_clock; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_reset; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_0; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_1; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_2; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_3; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_4; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_ins_5; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_0; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_1; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_2; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_3; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_4; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_11_io_outs_5; // @[MemPrimitives.scala 124:33:@13930.4]
  wire  StickySelects_12_clock; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_reset; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_0; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_1; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_2; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_3; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_4; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_ins_5; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_0; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_1; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_2; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_3; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_4; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_12_io_outs_5; // @[MemPrimitives.scala 124:33:@13992.4]
  wire  StickySelects_13_clock; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_reset; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_0; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_1; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_2; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_3; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_4; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_ins_5; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_0; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_1; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_2; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_3; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_4; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_13_io_outs_5; // @[MemPrimitives.scala 124:33:@14054.4]
  wire  StickySelects_14_clock; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_reset; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_0; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_1; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_2; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_3; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_4; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_ins_5; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_0; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_1; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_2; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_3; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_4; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_14_io_outs_5; // @[MemPrimitives.scala 124:33:@14116.4]
  wire  StickySelects_15_clock; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_reset; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_0; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_1; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_2; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_3; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_4; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_ins_5; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_0; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_1; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_2; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_3; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_4; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  StickySelects_15_io_outs_5; // @[MemPrimitives.scala 124:33:@14178.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@14241.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@14249.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@14257.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@14265.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@14273.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@14281.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@14289.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@14297.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@14337.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@14345.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@14353.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_in; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_11_io_out; // @[package.scala 93:22:@14361.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@14369.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_in; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_13_io_out; // @[package.scala 93:22:@14377.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_in; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_14_io_out; // @[package.scala 93:22:@14385.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@14393.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_in; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_16_io_out; // @[package.scala 93:22:@14433.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@14441.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@14449.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_in; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_19_io_out; // @[package.scala 93:22:@14457.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_in; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_20_io_out; // @[package.scala 93:22:@14465.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@14473.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@14481.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_in; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_23_io_out; // @[package.scala 93:22:@14489.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@14529.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_in; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_25_io_out; // @[package.scala 93:22:@14537.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_in; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_26_io_out; // @[package.scala 93:22:@14545.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@14553.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_in; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_28_io_out; // @[package.scala 93:22:@14561.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_in; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_29_io_out; // @[package.scala 93:22:@14569.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_in; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_30_io_out; // @[package.scala 93:22:@14577.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@14585.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@14625.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_in; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_33_io_out; // @[package.scala 93:22:@14633.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_in; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_34_io_out; // @[package.scala 93:22:@14641.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@14649.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@14657.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_in; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_37_io_out; // @[package.scala 93:22:@14665.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_in; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_38_io_out; // @[package.scala 93:22:@14673.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@14681.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@14721.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@14729.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_in; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_42_io_out; // @[package.scala 93:22:@14737.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@14745.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@14753.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_in; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_45_io_out; // @[package.scala 93:22:@14761.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@14769.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@14777.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_in; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_48_io_out; // @[package.scala 93:22:@14817.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@14825.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@14833.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@14841.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_in; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_52_io_out; // @[package.scala 93:22:@14849.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@14857.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@14865.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@14873.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@14913.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@14921.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@14929.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@14937.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_in; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_60_io_out; // @[package.scala 93:22:@14945.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_in; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_61_io_out; // @[package.scala 93:22:@14953.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_in; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_62_io_out; // @[package.scala 93:22:@14961.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@14969.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@15009.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@15017.4]
  wire  RetimeWrapper_66_clock; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_reset; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_flow; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_in; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_66_io_out; // @[package.scala 93:22:@15025.4]
  wire  RetimeWrapper_67_clock; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_reset; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_flow; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_in; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_67_io_out; // @[package.scala 93:22:@15033.4]
  wire  RetimeWrapper_68_clock; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_reset; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_flow; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_in; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_68_io_out; // @[package.scala 93:22:@15041.4]
  wire  RetimeWrapper_69_clock; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_reset; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_flow; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_in; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_69_io_out; // @[package.scala 93:22:@15049.4]
  wire  RetimeWrapper_70_clock; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_reset; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_flow; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_in; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_70_io_out; // @[package.scala 93:22:@15057.4]
  wire  RetimeWrapper_71_clock; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_reset; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_flow; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_in; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_71_io_out; // @[package.scala 93:22:@15065.4]
  wire  RetimeWrapper_72_clock; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_reset; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_flow; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_in; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_72_io_out; // @[package.scala 93:22:@15105.4]
  wire  RetimeWrapper_73_clock; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_reset; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_flow; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_in; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_73_io_out; // @[package.scala 93:22:@15113.4]
  wire  RetimeWrapper_74_clock; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_reset; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_flow; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_in; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_74_io_out; // @[package.scala 93:22:@15121.4]
  wire  RetimeWrapper_75_clock; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_reset; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_flow; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_in; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_75_io_out; // @[package.scala 93:22:@15129.4]
  wire  RetimeWrapper_76_clock; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_reset; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_flow; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_in; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_76_io_out; // @[package.scala 93:22:@15137.4]
  wire  RetimeWrapper_77_clock; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_reset; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_flow; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_in; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_77_io_out; // @[package.scala 93:22:@15145.4]
  wire  RetimeWrapper_78_clock; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_reset; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_flow; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_in; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_78_io_out; // @[package.scala 93:22:@15153.4]
  wire  RetimeWrapper_79_clock; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_reset; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_flow; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_in; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_79_io_out; // @[package.scala 93:22:@15161.4]
  wire  RetimeWrapper_80_clock; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_reset; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_flow; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_in; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_80_io_out; // @[package.scala 93:22:@15201.4]
  wire  RetimeWrapper_81_clock; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_reset; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_flow; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_in; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_81_io_out; // @[package.scala 93:22:@15209.4]
  wire  RetimeWrapper_82_clock; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_reset; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_flow; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_in; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_82_io_out; // @[package.scala 93:22:@15217.4]
  wire  RetimeWrapper_83_clock; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_reset; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_flow; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_in; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_83_io_out; // @[package.scala 93:22:@15225.4]
  wire  RetimeWrapper_84_clock; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_reset; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_flow; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_in; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_84_io_out; // @[package.scala 93:22:@15233.4]
  wire  RetimeWrapper_85_clock; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_reset; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_flow; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_in; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_85_io_out; // @[package.scala 93:22:@15241.4]
  wire  RetimeWrapper_86_clock; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_reset; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_flow; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_in; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_86_io_out; // @[package.scala 93:22:@15249.4]
  wire  RetimeWrapper_87_clock; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_reset; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_flow; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_in; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_87_io_out; // @[package.scala 93:22:@15257.4]
  wire  RetimeWrapper_88_clock; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_reset; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_flow; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_in; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_88_io_out; // @[package.scala 93:22:@15297.4]
  wire  RetimeWrapper_89_clock; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_reset; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_flow; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_in; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_89_io_out; // @[package.scala 93:22:@15305.4]
  wire  RetimeWrapper_90_clock; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_reset; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_flow; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_in; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_90_io_out; // @[package.scala 93:22:@15313.4]
  wire  RetimeWrapper_91_clock; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_reset; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_flow; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_in; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_91_io_out; // @[package.scala 93:22:@15321.4]
  wire  RetimeWrapper_92_clock; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_reset; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_flow; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_in; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_92_io_out; // @[package.scala 93:22:@15329.4]
  wire  RetimeWrapper_93_clock; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_reset; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_flow; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_in; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_93_io_out; // @[package.scala 93:22:@15337.4]
  wire  RetimeWrapper_94_clock; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_reset; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_flow; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_in; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_94_io_out; // @[package.scala 93:22:@15345.4]
  wire  RetimeWrapper_95_clock; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_reset; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_flow; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_in; // @[package.scala 93:22:@15353.4]
  wire  RetimeWrapper_95_io_out; // @[package.scala 93:22:@15353.4]
  wire  _T_444; // @[MemPrimitives.scala 82:210:@13032.4]
  wire  _T_446; // @[MemPrimitives.scala 82:210:@13033.4]
  wire  _T_447; // @[MemPrimitives.scala 82:228:@13034.4]
  wire  _T_448; // @[MemPrimitives.scala 83:102:@13035.4]
  wire [41:0] _T_450; // @[Cat.scala 30:58:@13037.4]
  wire  _T_455; // @[MemPrimitives.scala 82:210:@13044.4]
  wire  _T_457; // @[MemPrimitives.scala 82:210:@13045.4]
  wire  _T_458; // @[MemPrimitives.scala 82:228:@13046.4]
  wire  _T_459; // @[MemPrimitives.scala 83:102:@13047.4]
  wire [41:0] _T_461; // @[Cat.scala 30:58:@13049.4]
  wire  _T_468; // @[MemPrimitives.scala 82:210:@13057.4]
  wire  _T_469; // @[MemPrimitives.scala 82:228:@13058.4]
  wire  _T_470; // @[MemPrimitives.scala 83:102:@13059.4]
  wire [41:0] _T_472; // @[Cat.scala 30:58:@13061.4]
  wire  _T_479; // @[MemPrimitives.scala 82:210:@13069.4]
  wire  _T_480; // @[MemPrimitives.scala 82:228:@13070.4]
  wire  _T_481; // @[MemPrimitives.scala 83:102:@13071.4]
  wire [41:0] _T_483; // @[Cat.scala 30:58:@13073.4]
  wire  _T_488; // @[MemPrimitives.scala 82:210:@13080.4]
  wire  _T_491; // @[MemPrimitives.scala 82:228:@13082.4]
  wire  _T_492; // @[MemPrimitives.scala 83:102:@13083.4]
  wire [41:0] _T_494; // @[Cat.scala 30:58:@13085.4]
  wire  _T_499; // @[MemPrimitives.scala 82:210:@13092.4]
  wire  _T_502; // @[MemPrimitives.scala 82:228:@13094.4]
  wire  _T_503; // @[MemPrimitives.scala 83:102:@13095.4]
  wire [41:0] _T_505; // @[Cat.scala 30:58:@13097.4]
  wire  _T_513; // @[MemPrimitives.scala 82:228:@13106.4]
  wire  _T_514; // @[MemPrimitives.scala 83:102:@13107.4]
  wire [41:0] _T_516; // @[Cat.scala 30:58:@13109.4]
  wire  _T_524; // @[MemPrimitives.scala 82:228:@13118.4]
  wire  _T_525; // @[MemPrimitives.scala 83:102:@13119.4]
  wire [41:0] _T_527; // @[Cat.scala 30:58:@13121.4]
  wire  _T_532; // @[MemPrimitives.scala 82:210:@13128.4]
  wire  _T_535; // @[MemPrimitives.scala 82:228:@13130.4]
  wire  _T_536; // @[MemPrimitives.scala 83:102:@13131.4]
  wire [41:0] _T_538; // @[Cat.scala 30:58:@13133.4]
  wire  _T_543; // @[MemPrimitives.scala 82:210:@13140.4]
  wire  _T_546; // @[MemPrimitives.scala 82:228:@13142.4]
  wire  _T_547; // @[MemPrimitives.scala 83:102:@13143.4]
  wire [41:0] _T_549; // @[Cat.scala 30:58:@13145.4]
  wire  _T_557; // @[MemPrimitives.scala 82:228:@13154.4]
  wire  _T_558; // @[MemPrimitives.scala 83:102:@13155.4]
  wire [41:0] _T_560; // @[Cat.scala 30:58:@13157.4]
  wire  _T_568; // @[MemPrimitives.scala 82:228:@13166.4]
  wire  _T_569; // @[MemPrimitives.scala 83:102:@13167.4]
  wire [41:0] _T_571; // @[Cat.scala 30:58:@13169.4]
  wire  _T_576; // @[MemPrimitives.scala 82:210:@13176.4]
  wire  _T_579; // @[MemPrimitives.scala 82:228:@13178.4]
  wire  _T_580; // @[MemPrimitives.scala 83:102:@13179.4]
  wire [41:0] _T_582; // @[Cat.scala 30:58:@13181.4]
  wire  _T_587; // @[MemPrimitives.scala 82:210:@13188.4]
  wire  _T_590; // @[MemPrimitives.scala 82:228:@13190.4]
  wire  _T_591; // @[MemPrimitives.scala 83:102:@13191.4]
  wire [41:0] _T_593; // @[Cat.scala 30:58:@13193.4]
  wire  _T_601; // @[MemPrimitives.scala 82:228:@13202.4]
  wire  _T_602; // @[MemPrimitives.scala 83:102:@13203.4]
  wire [41:0] _T_604; // @[Cat.scala 30:58:@13205.4]
  wire  _T_612; // @[MemPrimitives.scala 82:228:@13214.4]
  wire  _T_613; // @[MemPrimitives.scala 83:102:@13215.4]
  wire [41:0] _T_615; // @[Cat.scala 30:58:@13217.4]
  wire  _T_620; // @[MemPrimitives.scala 110:210:@13224.4]
  wire  _T_622; // @[MemPrimitives.scala 110:210:@13225.4]
  wire  _T_623; // @[MemPrimitives.scala 110:228:@13226.4]
  wire  _T_626; // @[MemPrimitives.scala 110:210:@13228.4]
  wire  _T_628; // @[MemPrimitives.scala 110:210:@13229.4]
  wire  _T_629; // @[MemPrimitives.scala 110:228:@13230.4]
  wire  _T_632; // @[MemPrimitives.scala 110:210:@13232.4]
  wire  _T_634; // @[MemPrimitives.scala 110:210:@13233.4]
  wire  _T_635; // @[MemPrimitives.scala 110:228:@13234.4]
  wire  _T_638; // @[MemPrimitives.scala 110:210:@13236.4]
  wire  _T_640; // @[MemPrimitives.scala 110:210:@13237.4]
  wire  _T_641; // @[MemPrimitives.scala 110:228:@13238.4]
  wire  _T_644; // @[MemPrimitives.scala 110:210:@13240.4]
  wire  _T_646; // @[MemPrimitives.scala 110:210:@13241.4]
  wire  _T_647; // @[MemPrimitives.scala 110:228:@13242.4]
  wire  _T_650; // @[MemPrimitives.scala 110:210:@13244.4]
  wire  _T_652; // @[MemPrimitives.scala 110:210:@13245.4]
  wire  _T_653; // @[MemPrimitives.scala 110:228:@13246.4]
  wire  _T_655; // @[MemPrimitives.scala 126:35:@13257.4]
  wire  _T_656; // @[MemPrimitives.scala 126:35:@13258.4]
  wire  _T_657; // @[MemPrimitives.scala 126:35:@13259.4]
  wire  _T_658; // @[MemPrimitives.scala 126:35:@13260.4]
  wire  _T_659; // @[MemPrimitives.scala 126:35:@13261.4]
  wire  _T_660; // @[MemPrimitives.scala 126:35:@13262.4]
  wire [10:0] _T_662; // @[Cat.scala 30:58:@13264.4]
  wire [10:0] _T_664; // @[Cat.scala 30:58:@13266.4]
  wire [10:0] _T_666; // @[Cat.scala 30:58:@13268.4]
  wire [10:0] _T_668; // @[Cat.scala 30:58:@13270.4]
  wire [10:0] _T_670; // @[Cat.scala 30:58:@13272.4]
  wire [10:0] _T_672; // @[Cat.scala 30:58:@13274.4]
  wire [10:0] _T_673; // @[Mux.scala 31:69:@13275.4]
  wire [10:0] _T_674; // @[Mux.scala 31:69:@13276.4]
  wire [10:0] _T_675; // @[Mux.scala 31:69:@13277.4]
  wire [10:0] _T_676; // @[Mux.scala 31:69:@13278.4]
  wire [10:0] _T_677; // @[Mux.scala 31:69:@13279.4]
  wire  _T_682; // @[MemPrimitives.scala 110:210:@13286.4]
  wire  _T_684; // @[MemPrimitives.scala 110:210:@13287.4]
  wire  _T_685; // @[MemPrimitives.scala 110:228:@13288.4]
  wire  _T_688; // @[MemPrimitives.scala 110:210:@13290.4]
  wire  _T_690; // @[MemPrimitives.scala 110:210:@13291.4]
  wire  _T_691; // @[MemPrimitives.scala 110:228:@13292.4]
  wire  _T_694; // @[MemPrimitives.scala 110:210:@13294.4]
  wire  _T_696; // @[MemPrimitives.scala 110:210:@13295.4]
  wire  _T_697; // @[MemPrimitives.scala 110:228:@13296.4]
  wire  _T_700; // @[MemPrimitives.scala 110:210:@13298.4]
  wire  _T_702; // @[MemPrimitives.scala 110:210:@13299.4]
  wire  _T_703; // @[MemPrimitives.scala 110:228:@13300.4]
  wire  _T_706; // @[MemPrimitives.scala 110:210:@13302.4]
  wire  _T_708; // @[MemPrimitives.scala 110:210:@13303.4]
  wire  _T_709; // @[MemPrimitives.scala 110:228:@13304.4]
  wire  _T_712; // @[MemPrimitives.scala 110:210:@13306.4]
  wire  _T_714; // @[MemPrimitives.scala 110:210:@13307.4]
  wire  _T_715; // @[MemPrimitives.scala 110:228:@13308.4]
  wire  _T_717; // @[MemPrimitives.scala 126:35:@13319.4]
  wire  _T_718; // @[MemPrimitives.scala 126:35:@13320.4]
  wire  _T_719; // @[MemPrimitives.scala 126:35:@13321.4]
  wire  _T_720; // @[MemPrimitives.scala 126:35:@13322.4]
  wire  _T_721; // @[MemPrimitives.scala 126:35:@13323.4]
  wire  _T_722; // @[MemPrimitives.scala 126:35:@13324.4]
  wire [10:0] _T_724; // @[Cat.scala 30:58:@13326.4]
  wire [10:0] _T_726; // @[Cat.scala 30:58:@13328.4]
  wire [10:0] _T_728; // @[Cat.scala 30:58:@13330.4]
  wire [10:0] _T_730; // @[Cat.scala 30:58:@13332.4]
  wire [10:0] _T_732; // @[Cat.scala 30:58:@13334.4]
  wire [10:0] _T_734; // @[Cat.scala 30:58:@13336.4]
  wire [10:0] _T_735; // @[Mux.scala 31:69:@13337.4]
  wire [10:0] _T_736; // @[Mux.scala 31:69:@13338.4]
  wire [10:0] _T_737; // @[Mux.scala 31:69:@13339.4]
  wire [10:0] _T_738; // @[Mux.scala 31:69:@13340.4]
  wire [10:0] _T_739; // @[Mux.scala 31:69:@13341.4]
  wire  _T_746; // @[MemPrimitives.scala 110:210:@13349.4]
  wire  _T_747; // @[MemPrimitives.scala 110:228:@13350.4]
  wire  _T_752; // @[MemPrimitives.scala 110:210:@13353.4]
  wire  _T_753; // @[MemPrimitives.scala 110:228:@13354.4]
  wire  _T_758; // @[MemPrimitives.scala 110:210:@13357.4]
  wire  _T_759; // @[MemPrimitives.scala 110:228:@13358.4]
  wire  _T_764; // @[MemPrimitives.scala 110:210:@13361.4]
  wire  _T_765; // @[MemPrimitives.scala 110:228:@13362.4]
  wire  _T_770; // @[MemPrimitives.scala 110:210:@13365.4]
  wire  _T_771; // @[MemPrimitives.scala 110:228:@13366.4]
  wire  _T_776; // @[MemPrimitives.scala 110:210:@13369.4]
  wire  _T_777; // @[MemPrimitives.scala 110:228:@13370.4]
  wire  _T_779; // @[MemPrimitives.scala 126:35:@13381.4]
  wire  _T_780; // @[MemPrimitives.scala 126:35:@13382.4]
  wire  _T_781; // @[MemPrimitives.scala 126:35:@13383.4]
  wire  _T_782; // @[MemPrimitives.scala 126:35:@13384.4]
  wire  _T_783; // @[MemPrimitives.scala 126:35:@13385.4]
  wire  _T_784; // @[MemPrimitives.scala 126:35:@13386.4]
  wire [10:0] _T_786; // @[Cat.scala 30:58:@13388.4]
  wire [10:0] _T_788; // @[Cat.scala 30:58:@13390.4]
  wire [10:0] _T_790; // @[Cat.scala 30:58:@13392.4]
  wire [10:0] _T_792; // @[Cat.scala 30:58:@13394.4]
  wire [10:0] _T_794; // @[Cat.scala 30:58:@13396.4]
  wire [10:0] _T_796; // @[Cat.scala 30:58:@13398.4]
  wire [10:0] _T_797; // @[Mux.scala 31:69:@13399.4]
  wire [10:0] _T_798; // @[Mux.scala 31:69:@13400.4]
  wire [10:0] _T_799; // @[Mux.scala 31:69:@13401.4]
  wire [10:0] _T_800; // @[Mux.scala 31:69:@13402.4]
  wire [10:0] _T_801; // @[Mux.scala 31:69:@13403.4]
  wire  _T_808; // @[MemPrimitives.scala 110:210:@13411.4]
  wire  _T_809; // @[MemPrimitives.scala 110:228:@13412.4]
  wire  _T_814; // @[MemPrimitives.scala 110:210:@13415.4]
  wire  _T_815; // @[MemPrimitives.scala 110:228:@13416.4]
  wire  _T_820; // @[MemPrimitives.scala 110:210:@13419.4]
  wire  _T_821; // @[MemPrimitives.scala 110:228:@13420.4]
  wire  _T_826; // @[MemPrimitives.scala 110:210:@13423.4]
  wire  _T_827; // @[MemPrimitives.scala 110:228:@13424.4]
  wire  _T_832; // @[MemPrimitives.scala 110:210:@13427.4]
  wire  _T_833; // @[MemPrimitives.scala 110:228:@13428.4]
  wire  _T_838; // @[MemPrimitives.scala 110:210:@13431.4]
  wire  _T_839; // @[MemPrimitives.scala 110:228:@13432.4]
  wire  _T_841; // @[MemPrimitives.scala 126:35:@13443.4]
  wire  _T_842; // @[MemPrimitives.scala 126:35:@13444.4]
  wire  _T_843; // @[MemPrimitives.scala 126:35:@13445.4]
  wire  _T_844; // @[MemPrimitives.scala 126:35:@13446.4]
  wire  _T_845; // @[MemPrimitives.scala 126:35:@13447.4]
  wire  _T_846; // @[MemPrimitives.scala 126:35:@13448.4]
  wire [10:0] _T_848; // @[Cat.scala 30:58:@13450.4]
  wire [10:0] _T_850; // @[Cat.scala 30:58:@13452.4]
  wire [10:0] _T_852; // @[Cat.scala 30:58:@13454.4]
  wire [10:0] _T_854; // @[Cat.scala 30:58:@13456.4]
  wire [10:0] _T_856; // @[Cat.scala 30:58:@13458.4]
  wire [10:0] _T_858; // @[Cat.scala 30:58:@13460.4]
  wire [10:0] _T_859; // @[Mux.scala 31:69:@13461.4]
  wire [10:0] _T_860; // @[Mux.scala 31:69:@13462.4]
  wire [10:0] _T_861; // @[Mux.scala 31:69:@13463.4]
  wire [10:0] _T_862; // @[Mux.scala 31:69:@13464.4]
  wire [10:0] _T_863; // @[Mux.scala 31:69:@13465.4]
  wire  _T_868; // @[MemPrimitives.scala 110:210:@13472.4]
  wire  _T_871; // @[MemPrimitives.scala 110:228:@13474.4]
  wire  _T_874; // @[MemPrimitives.scala 110:210:@13476.4]
  wire  _T_877; // @[MemPrimitives.scala 110:228:@13478.4]
  wire  _T_880; // @[MemPrimitives.scala 110:210:@13480.4]
  wire  _T_883; // @[MemPrimitives.scala 110:228:@13482.4]
  wire  _T_886; // @[MemPrimitives.scala 110:210:@13484.4]
  wire  _T_889; // @[MemPrimitives.scala 110:228:@13486.4]
  wire  _T_892; // @[MemPrimitives.scala 110:210:@13488.4]
  wire  _T_895; // @[MemPrimitives.scala 110:228:@13490.4]
  wire  _T_898; // @[MemPrimitives.scala 110:210:@13492.4]
  wire  _T_901; // @[MemPrimitives.scala 110:228:@13494.4]
  wire  _T_903; // @[MemPrimitives.scala 126:35:@13505.4]
  wire  _T_904; // @[MemPrimitives.scala 126:35:@13506.4]
  wire  _T_905; // @[MemPrimitives.scala 126:35:@13507.4]
  wire  _T_906; // @[MemPrimitives.scala 126:35:@13508.4]
  wire  _T_907; // @[MemPrimitives.scala 126:35:@13509.4]
  wire  _T_908; // @[MemPrimitives.scala 126:35:@13510.4]
  wire [10:0] _T_910; // @[Cat.scala 30:58:@13512.4]
  wire [10:0] _T_912; // @[Cat.scala 30:58:@13514.4]
  wire [10:0] _T_914; // @[Cat.scala 30:58:@13516.4]
  wire [10:0] _T_916; // @[Cat.scala 30:58:@13518.4]
  wire [10:0] _T_918; // @[Cat.scala 30:58:@13520.4]
  wire [10:0] _T_920; // @[Cat.scala 30:58:@13522.4]
  wire [10:0] _T_921; // @[Mux.scala 31:69:@13523.4]
  wire [10:0] _T_922; // @[Mux.scala 31:69:@13524.4]
  wire [10:0] _T_923; // @[Mux.scala 31:69:@13525.4]
  wire [10:0] _T_924; // @[Mux.scala 31:69:@13526.4]
  wire [10:0] _T_925; // @[Mux.scala 31:69:@13527.4]
  wire  _T_930; // @[MemPrimitives.scala 110:210:@13534.4]
  wire  _T_933; // @[MemPrimitives.scala 110:228:@13536.4]
  wire  _T_936; // @[MemPrimitives.scala 110:210:@13538.4]
  wire  _T_939; // @[MemPrimitives.scala 110:228:@13540.4]
  wire  _T_942; // @[MemPrimitives.scala 110:210:@13542.4]
  wire  _T_945; // @[MemPrimitives.scala 110:228:@13544.4]
  wire  _T_948; // @[MemPrimitives.scala 110:210:@13546.4]
  wire  _T_951; // @[MemPrimitives.scala 110:228:@13548.4]
  wire  _T_954; // @[MemPrimitives.scala 110:210:@13550.4]
  wire  _T_957; // @[MemPrimitives.scala 110:228:@13552.4]
  wire  _T_960; // @[MemPrimitives.scala 110:210:@13554.4]
  wire  _T_963; // @[MemPrimitives.scala 110:228:@13556.4]
  wire  _T_965; // @[MemPrimitives.scala 126:35:@13567.4]
  wire  _T_966; // @[MemPrimitives.scala 126:35:@13568.4]
  wire  _T_967; // @[MemPrimitives.scala 126:35:@13569.4]
  wire  _T_968; // @[MemPrimitives.scala 126:35:@13570.4]
  wire  _T_969; // @[MemPrimitives.scala 126:35:@13571.4]
  wire  _T_970; // @[MemPrimitives.scala 126:35:@13572.4]
  wire [10:0] _T_972; // @[Cat.scala 30:58:@13574.4]
  wire [10:0] _T_974; // @[Cat.scala 30:58:@13576.4]
  wire [10:0] _T_976; // @[Cat.scala 30:58:@13578.4]
  wire [10:0] _T_978; // @[Cat.scala 30:58:@13580.4]
  wire [10:0] _T_980; // @[Cat.scala 30:58:@13582.4]
  wire [10:0] _T_982; // @[Cat.scala 30:58:@13584.4]
  wire [10:0] _T_983; // @[Mux.scala 31:69:@13585.4]
  wire [10:0] _T_984; // @[Mux.scala 31:69:@13586.4]
  wire [10:0] _T_985; // @[Mux.scala 31:69:@13587.4]
  wire [10:0] _T_986; // @[Mux.scala 31:69:@13588.4]
  wire [10:0] _T_987; // @[Mux.scala 31:69:@13589.4]
  wire  _T_995; // @[MemPrimitives.scala 110:228:@13598.4]
  wire  _T_1001; // @[MemPrimitives.scala 110:228:@13602.4]
  wire  _T_1007; // @[MemPrimitives.scala 110:228:@13606.4]
  wire  _T_1013; // @[MemPrimitives.scala 110:228:@13610.4]
  wire  _T_1019; // @[MemPrimitives.scala 110:228:@13614.4]
  wire  _T_1025; // @[MemPrimitives.scala 110:228:@13618.4]
  wire  _T_1027; // @[MemPrimitives.scala 126:35:@13629.4]
  wire  _T_1028; // @[MemPrimitives.scala 126:35:@13630.4]
  wire  _T_1029; // @[MemPrimitives.scala 126:35:@13631.4]
  wire  _T_1030; // @[MemPrimitives.scala 126:35:@13632.4]
  wire  _T_1031; // @[MemPrimitives.scala 126:35:@13633.4]
  wire  _T_1032; // @[MemPrimitives.scala 126:35:@13634.4]
  wire [10:0] _T_1034; // @[Cat.scala 30:58:@13636.4]
  wire [10:0] _T_1036; // @[Cat.scala 30:58:@13638.4]
  wire [10:0] _T_1038; // @[Cat.scala 30:58:@13640.4]
  wire [10:0] _T_1040; // @[Cat.scala 30:58:@13642.4]
  wire [10:0] _T_1042; // @[Cat.scala 30:58:@13644.4]
  wire [10:0] _T_1044; // @[Cat.scala 30:58:@13646.4]
  wire [10:0] _T_1045; // @[Mux.scala 31:69:@13647.4]
  wire [10:0] _T_1046; // @[Mux.scala 31:69:@13648.4]
  wire [10:0] _T_1047; // @[Mux.scala 31:69:@13649.4]
  wire [10:0] _T_1048; // @[Mux.scala 31:69:@13650.4]
  wire [10:0] _T_1049; // @[Mux.scala 31:69:@13651.4]
  wire  _T_1057; // @[MemPrimitives.scala 110:228:@13660.4]
  wire  _T_1063; // @[MemPrimitives.scala 110:228:@13664.4]
  wire  _T_1069; // @[MemPrimitives.scala 110:228:@13668.4]
  wire  _T_1075; // @[MemPrimitives.scala 110:228:@13672.4]
  wire  _T_1081; // @[MemPrimitives.scala 110:228:@13676.4]
  wire  _T_1087; // @[MemPrimitives.scala 110:228:@13680.4]
  wire  _T_1089; // @[MemPrimitives.scala 126:35:@13691.4]
  wire  _T_1090; // @[MemPrimitives.scala 126:35:@13692.4]
  wire  _T_1091; // @[MemPrimitives.scala 126:35:@13693.4]
  wire  _T_1092; // @[MemPrimitives.scala 126:35:@13694.4]
  wire  _T_1093; // @[MemPrimitives.scala 126:35:@13695.4]
  wire  _T_1094; // @[MemPrimitives.scala 126:35:@13696.4]
  wire [10:0] _T_1096; // @[Cat.scala 30:58:@13698.4]
  wire [10:0] _T_1098; // @[Cat.scala 30:58:@13700.4]
  wire [10:0] _T_1100; // @[Cat.scala 30:58:@13702.4]
  wire [10:0] _T_1102; // @[Cat.scala 30:58:@13704.4]
  wire [10:0] _T_1104; // @[Cat.scala 30:58:@13706.4]
  wire [10:0] _T_1106; // @[Cat.scala 30:58:@13708.4]
  wire [10:0] _T_1107; // @[Mux.scala 31:69:@13709.4]
  wire [10:0] _T_1108; // @[Mux.scala 31:69:@13710.4]
  wire [10:0] _T_1109; // @[Mux.scala 31:69:@13711.4]
  wire [10:0] _T_1110; // @[Mux.scala 31:69:@13712.4]
  wire [10:0] _T_1111; // @[Mux.scala 31:69:@13713.4]
  wire  _T_1116; // @[MemPrimitives.scala 110:210:@13720.4]
  wire  _T_1119; // @[MemPrimitives.scala 110:228:@13722.4]
  wire  _T_1122; // @[MemPrimitives.scala 110:210:@13724.4]
  wire  _T_1125; // @[MemPrimitives.scala 110:228:@13726.4]
  wire  _T_1128; // @[MemPrimitives.scala 110:210:@13728.4]
  wire  _T_1131; // @[MemPrimitives.scala 110:228:@13730.4]
  wire  _T_1134; // @[MemPrimitives.scala 110:210:@13732.4]
  wire  _T_1137; // @[MemPrimitives.scala 110:228:@13734.4]
  wire  _T_1140; // @[MemPrimitives.scala 110:210:@13736.4]
  wire  _T_1143; // @[MemPrimitives.scala 110:228:@13738.4]
  wire  _T_1146; // @[MemPrimitives.scala 110:210:@13740.4]
  wire  _T_1149; // @[MemPrimitives.scala 110:228:@13742.4]
  wire  _T_1151; // @[MemPrimitives.scala 126:35:@13753.4]
  wire  _T_1152; // @[MemPrimitives.scala 126:35:@13754.4]
  wire  _T_1153; // @[MemPrimitives.scala 126:35:@13755.4]
  wire  _T_1154; // @[MemPrimitives.scala 126:35:@13756.4]
  wire  _T_1155; // @[MemPrimitives.scala 126:35:@13757.4]
  wire  _T_1156; // @[MemPrimitives.scala 126:35:@13758.4]
  wire [10:0] _T_1158; // @[Cat.scala 30:58:@13760.4]
  wire [10:0] _T_1160; // @[Cat.scala 30:58:@13762.4]
  wire [10:0] _T_1162; // @[Cat.scala 30:58:@13764.4]
  wire [10:0] _T_1164; // @[Cat.scala 30:58:@13766.4]
  wire [10:0] _T_1166; // @[Cat.scala 30:58:@13768.4]
  wire [10:0] _T_1168; // @[Cat.scala 30:58:@13770.4]
  wire [10:0] _T_1169; // @[Mux.scala 31:69:@13771.4]
  wire [10:0] _T_1170; // @[Mux.scala 31:69:@13772.4]
  wire [10:0] _T_1171; // @[Mux.scala 31:69:@13773.4]
  wire [10:0] _T_1172; // @[Mux.scala 31:69:@13774.4]
  wire [10:0] _T_1173; // @[Mux.scala 31:69:@13775.4]
  wire  _T_1178; // @[MemPrimitives.scala 110:210:@13782.4]
  wire  _T_1181; // @[MemPrimitives.scala 110:228:@13784.4]
  wire  _T_1184; // @[MemPrimitives.scala 110:210:@13786.4]
  wire  _T_1187; // @[MemPrimitives.scala 110:228:@13788.4]
  wire  _T_1190; // @[MemPrimitives.scala 110:210:@13790.4]
  wire  _T_1193; // @[MemPrimitives.scala 110:228:@13792.4]
  wire  _T_1196; // @[MemPrimitives.scala 110:210:@13794.4]
  wire  _T_1199; // @[MemPrimitives.scala 110:228:@13796.4]
  wire  _T_1202; // @[MemPrimitives.scala 110:210:@13798.4]
  wire  _T_1205; // @[MemPrimitives.scala 110:228:@13800.4]
  wire  _T_1208; // @[MemPrimitives.scala 110:210:@13802.4]
  wire  _T_1211; // @[MemPrimitives.scala 110:228:@13804.4]
  wire  _T_1213; // @[MemPrimitives.scala 126:35:@13815.4]
  wire  _T_1214; // @[MemPrimitives.scala 126:35:@13816.4]
  wire  _T_1215; // @[MemPrimitives.scala 126:35:@13817.4]
  wire  _T_1216; // @[MemPrimitives.scala 126:35:@13818.4]
  wire  _T_1217; // @[MemPrimitives.scala 126:35:@13819.4]
  wire  _T_1218; // @[MemPrimitives.scala 126:35:@13820.4]
  wire [10:0] _T_1220; // @[Cat.scala 30:58:@13822.4]
  wire [10:0] _T_1222; // @[Cat.scala 30:58:@13824.4]
  wire [10:0] _T_1224; // @[Cat.scala 30:58:@13826.4]
  wire [10:0] _T_1226; // @[Cat.scala 30:58:@13828.4]
  wire [10:0] _T_1228; // @[Cat.scala 30:58:@13830.4]
  wire [10:0] _T_1230; // @[Cat.scala 30:58:@13832.4]
  wire [10:0] _T_1231; // @[Mux.scala 31:69:@13833.4]
  wire [10:0] _T_1232; // @[Mux.scala 31:69:@13834.4]
  wire [10:0] _T_1233; // @[Mux.scala 31:69:@13835.4]
  wire [10:0] _T_1234; // @[Mux.scala 31:69:@13836.4]
  wire [10:0] _T_1235; // @[Mux.scala 31:69:@13837.4]
  wire  _T_1243; // @[MemPrimitives.scala 110:228:@13846.4]
  wire  _T_1249; // @[MemPrimitives.scala 110:228:@13850.4]
  wire  _T_1255; // @[MemPrimitives.scala 110:228:@13854.4]
  wire  _T_1261; // @[MemPrimitives.scala 110:228:@13858.4]
  wire  _T_1267; // @[MemPrimitives.scala 110:228:@13862.4]
  wire  _T_1273; // @[MemPrimitives.scala 110:228:@13866.4]
  wire  _T_1275; // @[MemPrimitives.scala 126:35:@13877.4]
  wire  _T_1276; // @[MemPrimitives.scala 126:35:@13878.4]
  wire  _T_1277; // @[MemPrimitives.scala 126:35:@13879.4]
  wire  _T_1278; // @[MemPrimitives.scala 126:35:@13880.4]
  wire  _T_1279; // @[MemPrimitives.scala 126:35:@13881.4]
  wire  _T_1280; // @[MemPrimitives.scala 126:35:@13882.4]
  wire [10:0] _T_1282; // @[Cat.scala 30:58:@13884.4]
  wire [10:0] _T_1284; // @[Cat.scala 30:58:@13886.4]
  wire [10:0] _T_1286; // @[Cat.scala 30:58:@13888.4]
  wire [10:0] _T_1288; // @[Cat.scala 30:58:@13890.4]
  wire [10:0] _T_1290; // @[Cat.scala 30:58:@13892.4]
  wire [10:0] _T_1292; // @[Cat.scala 30:58:@13894.4]
  wire [10:0] _T_1293; // @[Mux.scala 31:69:@13895.4]
  wire [10:0] _T_1294; // @[Mux.scala 31:69:@13896.4]
  wire [10:0] _T_1295; // @[Mux.scala 31:69:@13897.4]
  wire [10:0] _T_1296; // @[Mux.scala 31:69:@13898.4]
  wire [10:0] _T_1297; // @[Mux.scala 31:69:@13899.4]
  wire  _T_1305; // @[MemPrimitives.scala 110:228:@13908.4]
  wire  _T_1311; // @[MemPrimitives.scala 110:228:@13912.4]
  wire  _T_1317; // @[MemPrimitives.scala 110:228:@13916.4]
  wire  _T_1323; // @[MemPrimitives.scala 110:228:@13920.4]
  wire  _T_1329; // @[MemPrimitives.scala 110:228:@13924.4]
  wire  _T_1335; // @[MemPrimitives.scala 110:228:@13928.4]
  wire  _T_1337; // @[MemPrimitives.scala 126:35:@13939.4]
  wire  _T_1338; // @[MemPrimitives.scala 126:35:@13940.4]
  wire  _T_1339; // @[MemPrimitives.scala 126:35:@13941.4]
  wire  _T_1340; // @[MemPrimitives.scala 126:35:@13942.4]
  wire  _T_1341; // @[MemPrimitives.scala 126:35:@13943.4]
  wire  _T_1342; // @[MemPrimitives.scala 126:35:@13944.4]
  wire [10:0] _T_1344; // @[Cat.scala 30:58:@13946.4]
  wire [10:0] _T_1346; // @[Cat.scala 30:58:@13948.4]
  wire [10:0] _T_1348; // @[Cat.scala 30:58:@13950.4]
  wire [10:0] _T_1350; // @[Cat.scala 30:58:@13952.4]
  wire [10:0] _T_1352; // @[Cat.scala 30:58:@13954.4]
  wire [10:0] _T_1354; // @[Cat.scala 30:58:@13956.4]
  wire [10:0] _T_1355; // @[Mux.scala 31:69:@13957.4]
  wire [10:0] _T_1356; // @[Mux.scala 31:69:@13958.4]
  wire [10:0] _T_1357; // @[Mux.scala 31:69:@13959.4]
  wire [10:0] _T_1358; // @[Mux.scala 31:69:@13960.4]
  wire [10:0] _T_1359; // @[Mux.scala 31:69:@13961.4]
  wire  _T_1364; // @[MemPrimitives.scala 110:210:@13968.4]
  wire  _T_1367; // @[MemPrimitives.scala 110:228:@13970.4]
  wire  _T_1370; // @[MemPrimitives.scala 110:210:@13972.4]
  wire  _T_1373; // @[MemPrimitives.scala 110:228:@13974.4]
  wire  _T_1376; // @[MemPrimitives.scala 110:210:@13976.4]
  wire  _T_1379; // @[MemPrimitives.scala 110:228:@13978.4]
  wire  _T_1382; // @[MemPrimitives.scala 110:210:@13980.4]
  wire  _T_1385; // @[MemPrimitives.scala 110:228:@13982.4]
  wire  _T_1388; // @[MemPrimitives.scala 110:210:@13984.4]
  wire  _T_1391; // @[MemPrimitives.scala 110:228:@13986.4]
  wire  _T_1394; // @[MemPrimitives.scala 110:210:@13988.4]
  wire  _T_1397; // @[MemPrimitives.scala 110:228:@13990.4]
  wire  _T_1399; // @[MemPrimitives.scala 126:35:@14001.4]
  wire  _T_1400; // @[MemPrimitives.scala 126:35:@14002.4]
  wire  _T_1401; // @[MemPrimitives.scala 126:35:@14003.4]
  wire  _T_1402; // @[MemPrimitives.scala 126:35:@14004.4]
  wire  _T_1403; // @[MemPrimitives.scala 126:35:@14005.4]
  wire  _T_1404; // @[MemPrimitives.scala 126:35:@14006.4]
  wire [10:0] _T_1406; // @[Cat.scala 30:58:@14008.4]
  wire [10:0] _T_1408; // @[Cat.scala 30:58:@14010.4]
  wire [10:0] _T_1410; // @[Cat.scala 30:58:@14012.4]
  wire [10:0] _T_1412; // @[Cat.scala 30:58:@14014.4]
  wire [10:0] _T_1414; // @[Cat.scala 30:58:@14016.4]
  wire [10:0] _T_1416; // @[Cat.scala 30:58:@14018.4]
  wire [10:0] _T_1417; // @[Mux.scala 31:69:@14019.4]
  wire [10:0] _T_1418; // @[Mux.scala 31:69:@14020.4]
  wire [10:0] _T_1419; // @[Mux.scala 31:69:@14021.4]
  wire [10:0] _T_1420; // @[Mux.scala 31:69:@14022.4]
  wire [10:0] _T_1421; // @[Mux.scala 31:69:@14023.4]
  wire  _T_1426; // @[MemPrimitives.scala 110:210:@14030.4]
  wire  _T_1429; // @[MemPrimitives.scala 110:228:@14032.4]
  wire  _T_1432; // @[MemPrimitives.scala 110:210:@14034.4]
  wire  _T_1435; // @[MemPrimitives.scala 110:228:@14036.4]
  wire  _T_1438; // @[MemPrimitives.scala 110:210:@14038.4]
  wire  _T_1441; // @[MemPrimitives.scala 110:228:@14040.4]
  wire  _T_1444; // @[MemPrimitives.scala 110:210:@14042.4]
  wire  _T_1447; // @[MemPrimitives.scala 110:228:@14044.4]
  wire  _T_1450; // @[MemPrimitives.scala 110:210:@14046.4]
  wire  _T_1453; // @[MemPrimitives.scala 110:228:@14048.4]
  wire  _T_1456; // @[MemPrimitives.scala 110:210:@14050.4]
  wire  _T_1459; // @[MemPrimitives.scala 110:228:@14052.4]
  wire  _T_1461; // @[MemPrimitives.scala 126:35:@14063.4]
  wire  _T_1462; // @[MemPrimitives.scala 126:35:@14064.4]
  wire  _T_1463; // @[MemPrimitives.scala 126:35:@14065.4]
  wire  _T_1464; // @[MemPrimitives.scala 126:35:@14066.4]
  wire  _T_1465; // @[MemPrimitives.scala 126:35:@14067.4]
  wire  _T_1466; // @[MemPrimitives.scala 126:35:@14068.4]
  wire [10:0] _T_1468; // @[Cat.scala 30:58:@14070.4]
  wire [10:0] _T_1470; // @[Cat.scala 30:58:@14072.4]
  wire [10:0] _T_1472; // @[Cat.scala 30:58:@14074.4]
  wire [10:0] _T_1474; // @[Cat.scala 30:58:@14076.4]
  wire [10:0] _T_1476; // @[Cat.scala 30:58:@14078.4]
  wire [10:0] _T_1478; // @[Cat.scala 30:58:@14080.4]
  wire [10:0] _T_1479; // @[Mux.scala 31:69:@14081.4]
  wire [10:0] _T_1480; // @[Mux.scala 31:69:@14082.4]
  wire [10:0] _T_1481; // @[Mux.scala 31:69:@14083.4]
  wire [10:0] _T_1482; // @[Mux.scala 31:69:@14084.4]
  wire [10:0] _T_1483; // @[Mux.scala 31:69:@14085.4]
  wire  _T_1491; // @[MemPrimitives.scala 110:228:@14094.4]
  wire  _T_1497; // @[MemPrimitives.scala 110:228:@14098.4]
  wire  _T_1503; // @[MemPrimitives.scala 110:228:@14102.4]
  wire  _T_1509; // @[MemPrimitives.scala 110:228:@14106.4]
  wire  _T_1515; // @[MemPrimitives.scala 110:228:@14110.4]
  wire  _T_1521; // @[MemPrimitives.scala 110:228:@14114.4]
  wire  _T_1523; // @[MemPrimitives.scala 126:35:@14125.4]
  wire  _T_1524; // @[MemPrimitives.scala 126:35:@14126.4]
  wire  _T_1525; // @[MemPrimitives.scala 126:35:@14127.4]
  wire  _T_1526; // @[MemPrimitives.scala 126:35:@14128.4]
  wire  _T_1527; // @[MemPrimitives.scala 126:35:@14129.4]
  wire  _T_1528; // @[MemPrimitives.scala 126:35:@14130.4]
  wire [10:0] _T_1530; // @[Cat.scala 30:58:@14132.4]
  wire [10:0] _T_1532; // @[Cat.scala 30:58:@14134.4]
  wire [10:0] _T_1534; // @[Cat.scala 30:58:@14136.4]
  wire [10:0] _T_1536; // @[Cat.scala 30:58:@14138.4]
  wire [10:0] _T_1538; // @[Cat.scala 30:58:@14140.4]
  wire [10:0] _T_1540; // @[Cat.scala 30:58:@14142.4]
  wire [10:0] _T_1541; // @[Mux.scala 31:69:@14143.4]
  wire [10:0] _T_1542; // @[Mux.scala 31:69:@14144.4]
  wire [10:0] _T_1543; // @[Mux.scala 31:69:@14145.4]
  wire [10:0] _T_1544; // @[Mux.scala 31:69:@14146.4]
  wire [10:0] _T_1545; // @[Mux.scala 31:69:@14147.4]
  wire  _T_1553; // @[MemPrimitives.scala 110:228:@14156.4]
  wire  _T_1559; // @[MemPrimitives.scala 110:228:@14160.4]
  wire  _T_1565; // @[MemPrimitives.scala 110:228:@14164.4]
  wire  _T_1571; // @[MemPrimitives.scala 110:228:@14168.4]
  wire  _T_1577; // @[MemPrimitives.scala 110:228:@14172.4]
  wire  _T_1583; // @[MemPrimitives.scala 110:228:@14176.4]
  wire  _T_1585; // @[MemPrimitives.scala 126:35:@14187.4]
  wire  _T_1586; // @[MemPrimitives.scala 126:35:@14188.4]
  wire  _T_1587; // @[MemPrimitives.scala 126:35:@14189.4]
  wire  _T_1588; // @[MemPrimitives.scala 126:35:@14190.4]
  wire  _T_1589; // @[MemPrimitives.scala 126:35:@14191.4]
  wire  _T_1590; // @[MemPrimitives.scala 126:35:@14192.4]
  wire [10:0] _T_1592; // @[Cat.scala 30:58:@14194.4]
  wire [10:0] _T_1594; // @[Cat.scala 30:58:@14196.4]
  wire [10:0] _T_1596; // @[Cat.scala 30:58:@14198.4]
  wire [10:0] _T_1598; // @[Cat.scala 30:58:@14200.4]
  wire [10:0] _T_1600; // @[Cat.scala 30:58:@14202.4]
  wire [10:0] _T_1602; // @[Cat.scala 30:58:@14204.4]
  wire [10:0] _T_1603; // @[Mux.scala 31:69:@14205.4]
  wire [10:0] _T_1604; // @[Mux.scala 31:69:@14206.4]
  wire [10:0] _T_1605; // @[Mux.scala 31:69:@14207.4]
  wire [10:0] _T_1606; // @[Mux.scala 31:69:@14208.4]
  wire [10:0] _T_1607; // @[Mux.scala 31:69:@14209.4]
  wire  _T_1671; // @[package.scala 96:25:@14294.4 package.scala 96:25:@14295.4]
  wire [31:0] _T_1675; // @[Mux.scala 31:69:@14304.4]
  wire  _T_1668; // @[package.scala 96:25:@14286.4 package.scala 96:25:@14287.4]
  wire [31:0] _T_1676; // @[Mux.scala 31:69:@14305.4]
  wire  _T_1665; // @[package.scala 96:25:@14278.4 package.scala 96:25:@14279.4]
  wire [31:0] _T_1677; // @[Mux.scala 31:69:@14306.4]
  wire  _T_1662; // @[package.scala 96:25:@14270.4 package.scala 96:25:@14271.4]
  wire [31:0] _T_1678; // @[Mux.scala 31:69:@14307.4]
  wire  _T_1659; // @[package.scala 96:25:@14262.4 package.scala 96:25:@14263.4]
  wire [31:0] _T_1679; // @[Mux.scala 31:69:@14308.4]
  wire  _T_1656; // @[package.scala 96:25:@14254.4 package.scala 96:25:@14255.4]
  wire [31:0] _T_1680; // @[Mux.scala 31:69:@14309.4]
  wire  _T_1653; // @[package.scala 96:25:@14246.4 package.scala 96:25:@14247.4]
  wire  _T_1742; // @[package.scala 96:25:@14390.4 package.scala 96:25:@14391.4]
  wire [31:0] _T_1746; // @[Mux.scala 31:69:@14400.4]
  wire  _T_1739; // @[package.scala 96:25:@14382.4 package.scala 96:25:@14383.4]
  wire [31:0] _T_1747; // @[Mux.scala 31:69:@14401.4]
  wire  _T_1736; // @[package.scala 96:25:@14374.4 package.scala 96:25:@14375.4]
  wire [31:0] _T_1748; // @[Mux.scala 31:69:@14402.4]
  wire  _T_1733; // @[package.scala 96:25:@14366.4 package.scala 96:25:@14367.4]
  wire [31:0] _T_1749; // @[Mux.scala 31:69:@14403.4]
  wire  _T_1730; // @[package.scala 96:25:@14358.4 package.scala 96:25:@14359.4]
  wire [31:0] _T_1750; // @[Mux.scala 31:69:@14404.4]
  wire  _T_1727; // @[package.scala 96:25:@14350.4 package.scala 96:25:@14351.4]
  wire [31:0] _T_1751; // @[Mux.scala 31:69:@14405.4]
  wire  _T_1724; // @[package.scala 96:25:@14342.4 package.scala 96:25:@14343.4]
  wire  _T_1813; // @[package.scala 96:25:@14486.4 package.scala 96:25:@14487.4]
  wire [31:0] _T_1817; // @[Mux.scala 31:69:@14496.4]
  wire  _T_1810; // @[package.scala 96:25:@14478.4 package.scala 96:25:@14479.4]
  wire [31:0] _T_1818; // @[Mux.scala 31:69:@14497.4]
  wire  _T_1807; // @[package.scala 96:25:@14470.4 package.scala 96:25:@14471.4]
  wire [31:0] _T_1819; // @[Mux.scala 31:69:@14498.4]
  wire  _T_1804; // @[package.scala 96:25:@14462.4 package.scala 96:25:@14463.4]
  wire [31:0] _T_1820; // @[Mux.scala 31:69:@14499.4]
  wire  _T_1801; // @[package.scala 96:25:@14454.4 package.scala 96:25:@14455.4]
  wire [31:0] _T_1821; // @[Mux.scala 31:69:@14500.4]
  wire  _T_1798; // @[package.scala 96:25:@14446.4 package.scala 96:25:@14447.4]
  wire [31:0] _T_1822; // @[Mux.scala 31:69:@14501.4]
  wire  _T_1795; // @[package.scala 96:25:@14438.4 package.scala 96:25:@14439.4]
  wire  _T_1884; // @[package.scala 96:25:@14582.4 package.scala 96:25:@14583.4]
  wire [31:0] _T_1888; // @[Mux.scala 31:69:@14592.4]
  wire  _T_1881; // @[package.scala 96:25:@14574.4 package.scala 96:25:@14575.4]
  wire [31:0] _T_1889; // @[Mux.scala 31:69:@14593.4]
  wire  _T_1878; // @[package.scala 96:25:@14566.4 package.scala 96:25:@14567.4]
  wire [31:0] _T_1890; // @[Mux.scala 31:69:@14594.4]
  wire  _T_1875; // @[package.scala 96:25:@14558.4 package.scala 96:25:@14559.4]
  wire [31:0] _T_1891; // @[Mux.scala 31:69:@14595.4]
  wire  _T_1872; // @[package.scala 96:25:@14550.4 package.scala 96:25:@14551.4]
  wire [31:0] _T_1892; // @[Mux.scala 31:69:@14596.4]
  wire  _T_1869; // @[package.scala 96:25:@14542.4 package.scala 96:25:@14543.4]
  wire [31:0] _T_1893; // @[Mux.scala 31:69:@14597.4]
  wire  _T_1866; // @[package.scala 96:25:@14534.4 package.scala 96:25:@14535.4]
  wire  _T_1955; // @[package.scala 96:25:@14678.4 package.scala 96:25:@14679.4]
  wire [31:0] _T_1959; // @[Mux.scala 31:69:@14688.4]
  wire  _T_1952; // @[package.scala 96:25:@14670.4 package.scala 96:25:@14671.4]
  wire [31:0] _T_1960; // @[Mux.scala 31:69:@14689.4]
  wire  _T_1949; // @[package.scala 96:25:@14662.4 package.scala 96:25:@14663.4]
  wire [31:0] _T_1961; // @[Mux.scala 31:69:@14690.4]
  wire  _T_1946; // @[package.scala 96:25:@14654.4 package.scala 96:25:@14655.4]
  wire [31:0] _T_1962; // @[Mux.scala 31:69:@14691.4]
  wire  _T_1943; // @[package.scala 96:25:@14646.4 package.scala 96:25:@14647.4]
  wire [31:0] _T_1963; // @[Mux.scala 31:69:@14692.4]
  wire  _T_1940; // @[package.scala 96:25:@14638.4 package.scala 96:25:@14639.4]
  wire [31:0] _T_1964; // @[Mux.scala 31:69:@14693.4]
  wire  _T_1937; // @[package.scala 96:25:@14630.4 package.scala 96:25:@14631.4]
  wire  _T_2026; // @[package.scala 96:25:@14774.4 package.scala 96:25:@14775.4]
  wire [31:0] _T_2030; // @[Mux.scala 31:69:@14784.4]
  wire  _T_2023; // @[package.scala 96:25:@14766.4 package.scala 96:25:@14767.4]
  wire [31:0] _T_2031; // @[Mux.scala 31:69:@14785.4]
  wire  _T_2020; // @[package.scala 96:25:@14758.4 package.scala 96:25:@14759.4]
  wire [31:0] _T_2032; // @[Mux.scala 31:69:@14786.4]
  wire  _T_2017; // @[package.scala 96:25:@14750.4 package.scala 96:25:@14751.4]
  wire [31:0] _T_2033; // @[Mux.scala 31:69:@14787.4]
  wire  _T_2014; // @[package.scala 96:25:@14742.4 package.scala 96:25:@14743.4]
  wire [31:0] _T_2034; // @[Mux.scala 31:69:@14788.4]
  wire  _T_2011; // @[package.scala 96:25:@14734.4 package.scala 96:25:@14735.4]
  wire [31:0] _T_2035; // @[Mux.scala 31:69:@14789.4]
  wire  _T_2008; // @[package.scala 96:25:@14726.4 package.scala 96:25:@14727.4]
  wire  _T_2097; // @[package.scala 96:25:@14870.4 package.scala 96:25:@14871.4]
  wire [31:0] _T_2101; // @[Mux.scala 31:69:@14880.4]
  wire  _T_2094; // @[package.scala 96:25:@14862.4 package.scala 96:25:@14863.4]
  wire [31:0] _T_2102; // @[Mux.scala 31:69:@14881.4]
  wire  _T_2091; // @[package.scala 96:25:@14854.4 package.scala 96:25:@14855.4]
  wire [31:0] _T_2103; // @[Mux.scala 31:69:@14882.4]
  wire  _T_2088; // @[package.scala 96:25:@14846.4 package.scala 96:25:@14847.4]
  wire [31:0] _T_2104; // @[Mux.scala 31:69:@14883.4]
  wire  _T_2085; // @[package.scala 96:25:@14838.4 package.scala 96:25:@14839.4]
  wire [31:0] _T_2105; // @[Mux.scala 31:69:@14884.4]
  wire  _T_2082; // @[package.scala 96:25:@14830.4 package.scala 96:25:@14831.4]
  wire [31:0] _T_2106; // @[Mux.scala 31:69:@14885.4]
  wire  _T_2079; // @[package.scala 96:25:@14822.4 package.scala 96:25:@14823.4]
  wire  _T_2168; // @[package.scala 96:25:@14966.4 package.scala 96:25:@14967.4]
  wire [31:0] _T_2172; // @[Mux.scala 31:69:@14976.4]
  wire  _T_2165; // @[package.scala 96:25:@14958.4 package.scala 96:25:@14959.4]
  wire [31:0] _T_2173; // @[Mux.scala 31:69:@14977.4]
  wire  _T_2162; // @[package.scala 96:25:@14950.4 package.scala 96:25:@14951.4]
  wire [31:0] _T_2174; // @[Mux.scala 31:69:@14978.4]
  wire  _T_2159; // @[package.scala 96:25:@14942.4 package.scala 96:25:@14943.4]
  wire [31:0] _T_2175; // @[Mux.scala 31:69:@14979.4]
  wire  _T_2156; // @[package.scala 96:25:@14934.4 package.scala 96:25:@14935.4]
  wire [31:0] _T_2176; // @[Mux.scala 31:69:@14980.4]
  wire  _T_2153; // @[package.scala 96:25:@14926.4 package.scala 96:25:@14927.4]
  wire [31:0] _T_2177; // @[Mux.scala 31:69:@14981.4]
  wire  _T_2150; // @[package.scala 96:25:@14918.4 package.scala 96:25:@14919.4]
  wire  _T_2239; // @[package.scala 96:25:@15062.4 package.scala 96:25:@15063.4]
  wire [31:0] _T_2243; // @[Mux.scala 31:69:@15072.4]
  wire  _T_2236; // @[package.scala 96:25:@15054.4 package.scala 96:25:@15055.4]
  wire [31:0] _T_2244; // @[Mux.scala 31:69:@15073.4]
  wire  _T_2233; // @[package.scala 96:25:@15046.4 package.scala 96:25:@15047.4]
  wire [31:0] _T_2245; // @[Mux.scala 31:69:@15074.4]
  wire  _T_2230; // @[package.scala 96:25:@15038.4 package.scala 96:25:@15039.4]
  wire [31:0] _T_2246; // @[Mux.scala 31:69:@15075.4]
  wire  _T_2227; // @[package.scala 96:25:@15030.4 package.scala 96:25:@15031.4]
  wire [31:0] _T_2247; // @[Mux.scala 31:69:@15076.4]
  wire  _T_2224; // @[package.scala 96:25:@15022.4 package.scala 96:25:@15023.4]
  wire [31:0] _T_2248; // @[Mux.scala 31:69:@15077.4]
  wire  _T_2221; // @[package.scala 96:25:@15014.4 package.scala 96:25:@15015.4]
  wire  _T_2310; // @[package.scala 96:25:@15158.4 package.scala 96:25:@15159.4]
  wire [31:0] _T_2314; // @[Mux.scala 31:69:@15168.4]
  wire  _T_2307; // @[package.scala 96:25:@15150.4 package.scala 96:25:@15151.4]
  wire [31:0] _T_2315; // @[Mux.scala 31:69:@15169.4]
  wire  _T_2304; // @[package.scala 96:25:@15142.4 package.scala 96:25:@15143.4]
  wire [31:0] _T_2316; // @[Mux.scala 31:69:@15170.4]
  wire  _T_2301; // @[package.scala 96:25:@15134.4 package.scala 96:25:@15135.4]
  wire [31:0] _T_2317; // @[Mux.scala 31:69:@15171.4]
  wire  _T_2298; // @[package.scala 96:25:@15126.4 package.scala 96:25:@15127.4]
  wire [31:0] _T_2318; // @[Mux.scala 31:69:@15172.4]
  wire  _T_2295; // @[package.scala 96:25:@15118.4 package.scala 96:25:@15119.4]
  wire [31:0] _T_2319; // @[Mux.scala 31:69:@15173.4]
  wire  _T_2292; // @[package.scala 96:25:@15110.4 package.scala 96:25:@15111.4]
  wire  _T_2381; // @[package.scala 96:25:@15254.4 package.scala 96:25:@15255.4]
  wire [31:0] _T_2385; // @[Mux.scala 31:69:@15264.4]
  wire  _T_2378; // @[package.scala 96:25:@15246.4 package.scala 96:25:@15247.4]
  wire [31:0] _T_2386; // @[Mux.scala 31:69:@15265.4]
  wire  _T_2375; // @[package.scala 96:25:@15238.4 package.scala 96:25:@15239.4]
  wire [31:0] _T_2387; // @[Mux.scala 31:69:@15266.4]
  wire  _T_2372; // @[package.scala 96:25:@15230.4 package.scala 96:25:@15231.4]
  wire [31:0] _T_2388; // @[Mux.scala 31:69:@15267.4]
  wire  _T_2369; // @[package.scala 96:25:@15222.4 package.scala 96:25:@15223.4]
  wire [31:0] _T_2389; // @[Mux.scala 31:69:@15268.4]
  wire  _T_2366; // @[package.scala 96:25:@15214.4 package.scala 96:25:@15215.4]
  wire [31:0] _T_2390; // @[Mux.scala 31:69:@15269.4]
  wire  _T_2363; // @[package.scala 96:25:@15206.4 package.scala 96:25:@15207.4]
  wire  _T_2452; // @[package.scala 96:25:@15350.4 package.scala 96:25:@15351.4]
  wire [31:0] _T_2456; // @[Mux.scala 31:69:@15360.4]
  wire  _T_2449; // @[package.scala 96:25:@15342.4 package.scala 96:25:@15343.4]
  wire [31:0] _T_2457; // @[Mux.scala 31:69:@15361.4]
  wire  _T_2446; // @[package.scala 96:25:@15334.4 package.scala 96:25:@15335.4]
  wire [31:0] _T_2458; // @[Mux.scala 31:69:@15362.4]
  wire  _T_2443; // @[package.scala 96:25:@15326.4 package.scala 96:25:@15327.4]
  wire [31:0] _T_2459; // @[Mux.scala 31:69:@15363.4]
  wire  _T_2440; // @[package.scala 96:25:@15318.4 package.scala 96:25:@15319.4]
  wire [31:0] _T_2460; // @[Mux.scala 31:69:@15364.4]
  wire  _T_2437; // @[package.scala 96:25:@15310.4 package.scala 96:25:@15311.4]
  wire [31:0] _T_2461; // @[Mux.scala 31:69:@15365.4]
  wire  _T_2434; // @[package.scala 96:25:@15302.4 package.scala 96:25:@15303.4]
  Mem1D_5 Mem1D ( // @[MemPrimitives.scala 64:21:@12776.4]
    .clock(Mem1D_clock),
    .reset(Mem1D_reset),
    .io_r_ofs_0(Mem1D_io_r_ofs_0),
    .io_r_backpressure(Mem1D_io_r_backpressure),
    .io_w_ofs_0(Mem1D_io_w_ofs_0),
    .io_w_data_0(Mem1D_io_w_data_0),
    .io_w_en_0(Mem1D_io_w_en_0),
    .io_output(Mem1D_io_output)
  );
  Mem1D_5 Mem1D_1 ( // @[MemPrimitives.scala 64:21:@12792.4]
    .clock(Mem1D_1_clock),
    .reset(Mem1D_1_reset),
    .io_r_ofs_0(Mem1D_1_io_r_ofs_0),
    .io_r_backpressure(Mem1D_1_io_r_backpressure),
    .io_w_ofs_0(Mem1D_1_io_w_ofs_0),
    .io_w_data_0(Mem1D_1_io_w_data_0),
    .io_w_en_0(Mem1D_1_io_w_en_0),
    .io_output(Mem1D_1_io_output)
  );
  Mem1D_5 Mem1D_2 ( // @[MemPrimitives.scala 64:21:@12808.4]
    .clock(Mem1D_2_clock),
    .reset(Mem1D_2_reset),
    .io_r_ofs_0(Mem1D_2_io_r_ofs_0),
    .io_r_backpressure(Mem1D_2_io_r_backpressure),
    .io_w_ofs_0(Mem1D_2_io_w_ofs_0),
    .io_w_data_0(Mem1D_2_io_w_data_0),
    .io_w_en_0(Mem1D_2_io_w_en_0),
    .io_output(Mem1D_2_io_output)
  );
  Mem1D_5 Mem1D_3 ( // @[MemPrimitives.scala 64:21:@12824.4]
    .clock(Mem1D_3_clock),
    .reset(Mem1D_3_reset),
    .io_r_ofs_0(Mem1D_3_io_r_ofs_0),
    .io_r_backpressure(Mem1D_3_io_r_backpressure),
    .io_w_ofs_0(Mem1D_3_io_w_ofs_0),
    .io_w_data_0(Mem1D_3_io_w_data_0),
    .io_w_en_0(Mem1D_3_io_w_en_0),
    .io_output(Mem1D_3_io_output)
  );
  Mem1D_5 Mem1D_4 ( // @[MemPrimitives.scala 64:21:@12840.4]
    .clock(Mem1D_4_clock),
    .reset(Mem1D_4_reset),
    .io_r_ofs_0(Mem1D_4_io_r_ofs_0),
    .io_r_backpressure(Mem1D_4_io_r_backpressure),
    .io_w_ofs_0(Mem1D_4_io_w_ofs_0),
    .io_w_data_0(Mem1D_4_io_w_data_0),
    .io_w_en_0(Mem1D_4_io_w_en_0),
    .io_output(Mem1D_4_io_output)
  );
  Mem1D_5 Mem1D_5 ( // @[MemPrimitives.scala 64:21:@12856.4]
    .clock(Mem1D_5_clock),
    .reset(Mem1D_5_reset),
    .io_r_ofs_0(Mem1D_5_io_r_ofs_0),
    .io_r_backpressure(Mem1D_5_io_r_backpressure),
    .io_w_ofs_0(Mem1D_5_io_w_ofs_0),
    .io_w_data_0(Mem1D_5_io_w_data_0),
    .io_w_en_0(Mem1D_5_io_w_en_0),
    .io_output(Mem1D_5_io_output)
  );
  Mem1D_5 Mem1D_6 ( // @[MemPrimitives.scala 64:21:@12872.4]
    .clock(Mem1D_6_clock),
    .reset(Mem1D_6_reset),
    .io_r_ofs_0(Mem1D_6_io_r_ofs_0),
    .io_r_backpressure(Mem1D_6_io_r_backpressure),
    .io_w_ofs_0(Mem1D_6_io_w_ofs_0),
    .io_w_data_0(Mem1D_6_io_w_data_0),
    .io_w_en_0(Mem1D_6_io_w_en_0),
    .io_output(Mem1D_6_io_output)
  );
  Mem1D_5 Mem1D_7 ( // @[MemPrimitives.scala 64:21:@12888.4]
    .clock(Mem1D_7_clock),
    .reset(Mem1D_7_reset),
    .io_r_ofs_0(Mem1D_7_io_r_ofs_0),
    .io_r_backpressure(Mem1D_7_io_r_backpressure),
    .io_w_ofs_0(Mem1D_7_io_w_ofs_0),
    .io_w_data_0(Mem1D_7_io_w_data_0),
    .io_w_en_0(Mem1D_7_io_w_en_0),
    .io_output(Mem1D_7_io_output)
  );
  Mem1D_5 Mem1D_8 ( // @[MemPrimitives.scala 64:21:@12904.4]
    .clock(Mem1D_8_clock),
    .reset(Mem1D_8_reset),
    .io_r_ofs_0(Mem1D_8_io_r_ofs_0),
    .io_r_backpressure(Mem1D_8_io_r_backpressure),
    .io_w_ofs_0(Mem1D_8_io_w_ofs_0),
    .io_w_data_0(Mem1D_8_io_w_data_0),
    .io_w_en_0(Mem1D_8_io_w_en_0),
    .io_output(Mem1D_8_io_output)
  );
  Mem1D_5 Mem1D_9 ( // @[MemPrimitives.scala 64:21:@12920.4]
    .clock(Mem1D_9_clock),
    .reset(Mem1D_9_reset),
    .io_r_ofs_0(Mem1D_9_io_r_ofs_0),
    .io_r_backpressure(Mem1D_9_io_r_backpressure),
    .io_w_ofs_0(Mem1D_9_io_w_ofs_0),
    .io_w_data_0(Mem1D_9_io_w_data_0),
    .io_w_en_0(Mem1D_9_io_w_en_0),
    .io_output(Mem1D_9_io_output)
  );
  Mem1D_5 Mem1D_10 ( // @[MemPrimitives.scala 64:21:@12936.4]
    .clock(Mem1D_10_clock),
    .reset(Mem1D_10_reset),
    .io_r_ofs_0(Mem1D_10_io_r_ofs_0),
    .io_r_backpressure(Mem1D_10_io_r_backpressure),
    .io_w_ofs_0(Mem1D_10_io_w_ofs_0),
    .io_w_data_0(Mem1D_10_io_w_data_0),
    .io_w_en_0(Mem1D_10_io_w_en_0),
    .io_output(Mem1D_10_io_output)
  );
  Mem1D_5 Mem1D_11 ( // @[MemPrimitives.scala 64:21:@12952.4]
    .clock(Mem1D_11_clock),
    .reset(Mem1D_11_reset),
    .io_r_ofs_0(Mem1D_11_io_r_ofs_0),
    .io_r_backpressure(Mem1D_11_io_r_backpressure),
    .io_w_ofs_0(Mem1D_11_io_w_ofs_0),
    .io_w_data_0(Mem1D_11_io_w_data_0),
    .io_w_en_0(Mem1D_11_io_w_en_0),
    .io_output(Mem1D_11_io_output)
  );
  Mem1D_5 Mem1D_12 ( // @[MemPrimitives.scala 64:21:@12968.4]
    .clock(Mem1D_12_clock),
    .reset(Mem1D_12_reset),
    .io_r_ofs_0(Mem1D_12_io_r_ofs_0),
    .io_r_backpressure(Mem1D_12_io_r_backpressure),
    .io_w_ofs_0(Mem1D_12_io_w_ofs_0),
    .io_w_data_0(Mem1D_12_io_w_data_0),
    .io_w_en_0(Mem1D_12_io_w_en_0),
    .io_output(Mem1D_12_io_output)
  );
  Mem1D_5 Mem1D_13 ( // @[MemPrimitives.scala 64:21:@12984.4]
    .clock(Mem1D_13_clock),
    .reset(Mem1D_13_reset),
    .io_r_ofs_0(Mem1D_13_io_r_ofs_0),
    .io_r_backpressure(Mem1D_13_io_r_backpressure),
    .io_w_ofs_0(Mem1D_13_io_w_ofs_0),
    .io_w_data_0(Mem1D_13_io_w_data_0),
    .io_w_en_0(Mem1D_13_io_w_en_0),
    .io_output(Mem1D_13_io_output)
  );
  Mem1D_5 Mem1D_14 ( // @[MemPrimitives.scala 64:21:@13000.4]
    .clock(Mem1D_14_clock),
    .reset(Mem1D_14_reset),
    .io_r_ofs_0(Mem1D_14_io_r_ofs_0),
    .io_r_backpressure(Mem1D_14_io_r_backpressure),
    .io_w_ofs_0(Mem1D_14_io_w_ofs_0),
    .io_w_data_0(Mem1D_14_io_w_data_0),
    .io_w_en_0(Mem1D_14_io_w_en_0),
    .io_output(Mem1D_14_io_output)
  );
  Mem1D_5 Mem1D_15 ( // @[MemPrimitives.scala 64:21:@13016.4]
    .clock(Mem1D_15_clock),
    .reset(Mem1D_15_reset),
    .io_r_ofs_0(Mem1D_15_io_r_ofs_0),
    .io_r_backpressure(Mem1D_15_io_r_backpressure),
    .io_w_ofs_0(Mem1D_15_io_w_ofs_0),
    .io_w_data_0(Mem1D_15_io_w_data_0),
    .io_w_en_0(Mem1D_15_io_w_en_0),
    .io_output(Mem1D_15_io_output)
  );
  StickySelects_1 StickySelects ( // @[MemPrimitives.scala 124:33:@13248.4]
    .clock(StickySelects_clock),
    .reset(StickySelects_reset),
    .io_ins_0(StickySelects_io_ins_0),
    .io_ins_1(StickySelects_io_ins_1),
    .io_ins_2(StickySelects_io_ins_2),
    .io_ins_3(StickySelects_io_ins_3),
    .io_ins_4(StickySelects_io_ins_4),
    .io_ins_5(StickySelects_io_ins_5),
    .io_outs_0(StickySelects_io_outs_0),
    .io_outs_1(StickySelects_io_outs_1),
    .io_outs_2(StickySelects_io_outs_2),
    .io_outs_3(StickySelects_io_outs_3),
    .io_outs_4(StickySelects_io_outs_4),
    .io_outs_5(StickySelects_io_outs_5)
  );
  StickySelects_1 StickySelects_1 ( // @[MemPrimitives.scala 124:33:@13310.4]
    .clock(StickySelects_1_clock),
    .reset(StickySelects_1_reset),
    .io_ins_0(StickySelects_1_io_ins_0),
    .io_ins_1(StickySelects_1_io_ins_1),
    .io_ins_2(StickySelects_1_io_ins_2),
    .io_ins_3(StickySelects_1_io_ins_3),
    .io_ins_4(StickySelects_1_io_ins_4),
    .io_ins_5(StickySelects_1_io_ins_5),
    .io_outs_0(StickySelects_1_io_outs_0),
    .io_outs_1(StickySelects_1_io_outs_1),
    .io_outs_2(StickySelects_1_io_outs_2),
    .io_outs_3(StickySelects_1_io_outs_3),
    .io_outs_4(StickySelects_1_io_outs_4),
    .io_outs_5(StickySelects_1_io_outs_5)
  );
  StickySelects_1 StickySelects_2 ( // @[MemPrimitives.scala 124:33:@13372.4]
    .clock(StickySelects_2_clock),
    .reset(StickySelects_2_reset),
    .io_ins_0(StickySelects_2_io_ins_0),
    .io_ins_1(StickySelects_2_io_ins_1),
    .io_ins_2(StickySelects_2_io_ins_2),
    .io_ins_3(StickySelects_2_io_ins_3),
    .io_ins_4(StickySelects_2_io_ins_4),
    .io_ins_5(StickySelects_2_io_ins_5),
    .io_outs_0(StickySelects_2_io_outs_0),
    .io_outs_1(StickySelects_2_io_outs_1),
    .io_outs_2(StickySelects_2_io_outs_2),
    .io_outs_3(StickySelects_2_io_outs_3),
    .io_outs_4(StickySelects_2_io_outs_4),
    .io_outs_5(StickySelects_2_io_outs_5)
  );
  StickySelects_1 StickySelects_3 ( // @[MemPrimitives.scala 124:33:@13434.4]
    .clock(StickySelects_3_clock),
    .reset(StickySelects_3_reset),
    .io_ins_0(StickySelects_3_io_ins_0),
    .io_ins_1(StickySelects_3_io_ins_1),
    .io_ins_2(StickySelects_3_io_ins_2),
    .io_ins_3(StickySelects_3_io_ins_3),
    .io_ins_4(StickySelects_3_io_ins_4),
    .io_ins_5(StickySelects_3_io_ins_5),
    .io_outs_0(StickySelects_3_io_outs_0),
    .io_outs_1(StickySelects_3_io_outs_1),
    .io_outs_2(StickySelects_3_io_outs_2),
    .io_outs_3(StickySelects_3_io_outs_3),
    .io_outs_4(StickySelects_3_io_outs_4),
    .io_outs_5(StickySelects_3_io_outs_5)
  );
  StickySelects_1 StickySelects_4 ( // @[MemPrimitives.scala 124:33:@13496.4]
    .clock(StickySelects_4_clock),
    .reset(StickySelects_4_reset),
    .io_ins_0(StickySelects_4_io_ins_0),
    .io_ins_1(StickySelects_4_io_ins_1),
    .io_ins_2(StickySelects_4_io_ins_2),
    .io_ins_3(StickySelects_4_io_ins_3),
    .io_ins_4(StickySelects_4_io_ins_4),
    .io_ins_5(StickySelects_4_io_ins_5),
    .io_outs_0(StickySelects_4_io_outs_0),
    .io_outs_1(StickySelects_4_io_outs_1),
    .io_outs_2(StickySelects_4_io_outs_2),
    .io_outs_3(StickySelects_4_io_outs_3),
    .io_outs_4(StickySelects_4_io_outs_4),
    .io_outs_5(StickySelects_4_io_outs_5)
  );
  StickySelects_1 StickySelects_5 ( // @[MemPrimitives.scala 124:33:@13558.4]
    .clock(StickySelects_5_clock),
    .reset(StickySelects_5_reset),
    .io_ins_0(StickySelects_5_io_ins_0),
    .io_ins_1(StickySelects_5_io_ins_1),
    .io_ins_2(StickySelects_5_io_ins_2),
    .io_ins_3(StickySelects_5_io_ins_3),
    .io_ins_4(StickySelects_5_io_ins_4),
    .io_ins_5(StickySelects_5_io_ins_5),
    .io_outs_0(StickySelects_5_io_outs_0),
    .io_outs_1(StickySelects_5_io_outs_1),
    .io_outs_2(StickySelects_5_io_outs_2),
    .io_outs_3(StickySelects_5_io_outs_3),
    .io_outs_4(StickySelects_5_io_outs_4),
    .io_outs_5(StickySelects_5_io_outs_5)
  );
  StickySelects_1 StickySelects_6 ( // @[MemPrimitives.scala 124:33:@13620.4]
    .clock(StickySelects_6_clock),
    .reset(StickySelects_6_reset),
    .io_ins_0(StickySelects_6_io_ins_0),
    .io_ins_1(StickySelects_6_io_ins_1),
    .io_ins_2(StickySelects_6_io_ins_2),
    .io_ins_3(StickySelects_6_io_ins_3),
    .io_ins_4(StickySelects_6_io_ins_4),
    .io_ins_5(StickySelects_6_io_ins_5),
    .io_outs_0(StickySelects_6_io_outs_0),
    .io_outs_1(StickySelects_6_io_outs_1),
    .io_outs_2(StickySelects_6_io_outs_2),
    .io_outs_3(StickySelects_6_io_outs_3),
    .io_outs_4(StickySelects_6_io_outs_4),
    .io_outs_5(StickySelects_6_io_outs_5)
  );
  StickySelects_1 StickySelects_7 ( // @[MemPrimitives.scala 124:33:@13682.4]
    .clock(StickySelects_7_clock),
    .reset(StickySelects_7_reset),
    .io_ins_0(StickySelects_7_io_ins_0),
    .io_ins_1(StickySelects_7_io_ins_1),
    .io_ins_2(StickySelects_7_io_ins_2),
    .io_ins_3(StickySelects_7_io_ins_3),
    .io_ins_4(StickySelects_7_io_ins_4),
    .io_ins_5(StickySelects_7_io_ins_5),
    .io_outs_0(StickySelects_7_io_outs_0),
    .io_outs_1(StickySelects_7_io_outs_1),
    .io_outs_2(StickySelects_7_io_outs_2),
    .io_outs_3(StickySelects_7_io_outs_3),
    .io_outs_4(StickySelects_7_io_outs_4),
    .io_outs_5(StickySelects_7_io_outs_5)
  );
  StickySelects_1 StickySelects_8 ( // @[MemPrimitives.scala 124:33:@13744.4]
    .clock(StickySelects_8_clock),
    .reset(StickySelects_8_reset),
    .io_ins_0(StickySelects_8_io_ins_0),
    .io_ins_1(StickySelects_8_io_ins_1),
    .io_ins_2(StickySelects_8_io_ins_2),
    .io_ins_3(StickySelects_8_io_ins_3),
    .io_ins_4(StickySelects_8_io_ins_4),
    .io_ins_5(StickySelects_8_io_ins_5),
    .io_outs_0(StickySelects_8_io_outs_0),
    .io_outs_1(StickySelects_8_io_outs_1),
    .io_outs_2(StickySelects_8_io_outs_2),
    .io_outs_3(StickySelects_8_io_outs_3),
    .io_outs_4(StickySelects_8_io_outs_4),
    .io_outs_5(StickySelects_8_io_outs_5)
  );
  StickySelects_1 StickySelects_9 ( // @[MemPrimitives.scala 124:33:@13806.4]
    .clock(StickySelects_9_clock),
    .reset(StickySelects_9_reset),
    .io_ins_0(StickySelects_9_io_ins_0),
    .io_ins_1(StickySelects_9_io_ins_1),
    .io_ins_2(StickySelects_9_io_ins_2),
    .io_ins_3(StickySelects_9_io_ins_3),
    .io_ins_4(StickySelects_9_io_ins_4),
    .io_ins_5(StickySelects_9_io_ins_5),
    .io_outs_0(StickySelects_9_io_outs_0),
    .io_outs_1(StickySelects_9_io_outs_1),
    .io_outs_2(StickySelects_9_io_outs_2),
    .io_outs_3(StickySelects_9_io_outs_3),
    .io_outs_4(StickySelects_9_io_outs_4),
    .io_outs_5(StickySelects_9_io_outs_5)
  );
  StickySelects_1 StickySelects_10 ( // @[MemPrimitives.scala 124:33:@13868.4]
    .clock(StickySelects_10_clock),
    .reset(StickySelects_10_reset),
    .io_ins_0(StickySelects_10_io_ins_0),
    .io_ins_1(StickySelects_10_io_ins_1),
    .io_ins_2(StickySelects_10_io_ins_2),
    .io_ins_3(StickySelects_10_io_ins_3),
    .io_ins_4(StickySelects_10_io_ins_4),
    .io_ins_5(StickySelects_10_io_ins_5),
    .io_outs_0(StickySelects_10_io_outs_0),
    .io_outs_1(StickySelects_10_io_outs_1),
    .io_outs_2(StickySelects_10_io_outs_2),
    .io_outs_3(StickySelects_10_io_outs_3),
    .io_outs_4(StickySelects_10_io_outs_4),
    .io_outs_5(StickySelects_10_io_outs_5)
  );
  StickySelects_1 StickySelects_11 ( // @[MemPrimitives.scala 124:33:@13930.4]
    .clock(StickySelects_11_clock),
    .reset(StickySelects_11_reset),
    .io_ins_0(StickySelects_11_io_ins_0),
    .io_ins_1(StickySelects_11_io_ins_1),
    .io_ins_2(StickySelects_11_io_ins_2),
    .io_ins_3(StickySelects_11_io_ins_3),
    .io_ins_4(StickySelects_11_io_ins_4),
    .io_ins_5(StickySelects_11_io_ins_5),
    .io_outs_0(StickySelects_11_io_outs_0),
    .io_outs_1(StickySelects_11_io_outs_1),
    .io_outs_2(StickySelects_11_io_outs_2),
    .io_outs_3(StickySelects_11_io_outs_3),
    .io_outs_4(StickySelects_11_io_outs_4),
    .io_outs_5(StickySelects_11_io_outs_5)
  );
  StickySelects_1 StickySelects_12 ( // @[MemPrimitives.scala 124:33:@13992.4]
    .clock(StickySelects_12_clock),
    .reset(StickySelects_12_reset),
    .io_ins_0(StickySelects_12_io_ins_0),
    .io_ins_1(StickySelects_12_io_ins_1),
    .io_ins_2(StickySelects_12_io_ins_2),
    .io_ins_3(StickySelects_12_io_ins_3),
    .io_ins_4(StickySelects_12_io_ins_4),
    .io_ins_5(StickySelects_12_io_ins_5),
    .io_outs_0(StickySelects_12_io_outs_0),
    .io_outs_1(StickySelects_12_io_outs_1),
    .io_outs_2(StickySelects_12_io_outs_2),
    .io_outs_3(StickySelects_12_io_outs_3),
    .io_outs_4(StickySelects_12_io_outs_4),
    .io_outs_5(StickySelects_12_io_outs_5)
  );
  StickySelects_1 StickySelects_13 ( // @[MemPrimitives.scala 124:33:@14054.4]
    .clock(StickySelects_13_clock),
    .reset(StickySelects_13_reset),
    .io_ins_0(StickySelects_13_io_ins_0),
    .io_ins_1(StickySelects_13_io_ins_1),
    .io_ins_2(StickySelects_13_io_ins_2),
    .io_ins_3(StickySelects_13_io_ins_3),
    .io_ins_4(StickySelects_13_io_ins_4),
    .io_ins_5(StickySelects_13_io_ins_5),
    .io_outs_0(StickySelects_13_io_outs_0),
    .io_outs_1(StickySelects_13_io_outs_1),
    .io_outs_2(StickySelects_13_io_outs_2),
    .io_outs_3(StickySelects_13_io_outs_3),
    .io_outs_4(StickySelects_13_io_outs_4),
    .io_outs_5(StickySelects_13_io_outs_5)
  );
  StickySelects_1 StickySelects_14 ( // @[MemPrimitives.scala 124:33:@14116.4]
    .clock(StickySelects_14_clock),
    .reset(StickySelects_14_reset),
    .io_ins_0(StickySelects_14_io_ins_0),
    .io_ins_1(StickySelects_14_io_ins_1),
    .io_ins_2(StickySelects_14_io_ins_2),
    .io_ins_3(StickySelects_14_io_ins_3),
    .io_ins_4(StickySelects_14_io_ins_4),
    .io_ins_5(StickySelects_14_io_ins_5),
    .io_outs_0(StickySelects_14_io_outs_0),
    .io_outs_1(StickySelects_14_io_outs_1),
    .io_outs_2(StickySelects_14_io_outs_2),
    .io_outs_3(StickySelects_14_io_outs_3),
    .io_outs_4(StickySelects_14_io_outs_4),
    .io_outs_5(StickySelects_14_io_outs_5)
  );
  StickySelects_1 StickySelects_15 ( // @[MemPrimitives.scala 124:33:@14178.4]
    .clock(StickySelects_15_clock),
    .reset(StickySelects_15_reset),
    .io_ins_0(StickySelects_15_io_ins_0),
    .io_ins_1(StickySelects_15_io_ins_1),
    .io_ins_2(StickySelects_15_io_ins_2),
    .io_ins_3(StickySelects_15_io_ins_3),
    .io_ins_4(StickySelects_15_io_ins_4),
    .io_ins_5(StickySelects_15_io_ins_5),
    .io_outs_0(StickySelects_15_io_outs_0),
    .io_outs_1(StickySelects_15_io_outs_1),
    .io_outs_2(StickySelects_15_io_outs_2),
    .io_outs_3(StickySelects_15_io_outs_3),
    .io_outs_4(StickySelects_15_io_outs_4),
    .io_outs_5(StickySelects_15_io_outs_5)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@14241.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@14249.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_2 ( // @[package.scala 93:22:@14257.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_3 ( // @[package.scala 93:22:@14265.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_4 ( // @[package.scala 93:22:@14273.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_5 ( // @[package.scala 93:22:@14281.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_6 ( // @[package.scala 93:22:@14289.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_7 ( // @[package.scala 93:22:@14297.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_8 ( // @[package.scala 93:22:@14337.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_9 ( // @[package.scala 93:22:@14345.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_10 ( // @[package.scala 93:22:@14353.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_11 ( // @[package.scala 93:22:@14361.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_12 ( // @[package.scala 93:22:@14369.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_13 ( // @[package.scala 93:22:@14377.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_14 ( // @[package.scala 93:22:@14385.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_15 ( // @[package.scala 93:22:@14393.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_16 ( // @[package.scala 93:22:@14433.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@14441.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_18 ( // @[package.scala 93:22:@14449.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_19 ( // @[package.scala 93:22:@14457.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_20 ( // @[package.scala 93:22:@14465.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_21 ( // @[package.scala 93:22:@14473.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_22 ( // @[package.scala 93:22:@14481.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_23 ( // @[package.scala 93:22:@14489.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_24 ( // @[package.scala 93:22:@14529.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_25 ( // @[package.scala 93:22:@14537.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_26 ( // @[package.scala 93:22:@14545.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_27 ( // @[package.scala 93:22:@14553.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_28 ( // @[package.scala 93:22:@14561.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_29 ( // @[package.scala 93:22:@14569.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_30 ( // @[package.scala 93:22:@14577.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@14585.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_32 ( // @[package.scala 93:22:@14625.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_33 ( // @[package.scala 93:22:@14633.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_34 ( // @[package.scala 93:22:@14641.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@14649.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_36 ( // @[package.scala 93:22:@14657.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_37 ( // @[package.scala 93:22:@14665.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_38 ( // @[package.scala 93:22:@14673.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@14681.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_40 ( // @[package.scala 93:22:@14721.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_41 ( // @[package.scala 93:22:@14729.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_42 ( // @[package.scala 93:22:@14737.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@14745.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_44 ( // @[package.scala 93:22:@14753.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_45 ( // @[package.scala 93:22:@14761.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@14769.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_47 ( // @[package.scala 93:22:@14777.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_48 ( // @[package.scala 93:22:@14817.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@14825.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_50 ( // @[package.scala 93:22:@14833.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@14841.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_52 ( // @[package.scala 93:22:@14849.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_53 ( // @[package.scala 93:22:@14857.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@14865.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_55 ( // @[package.scala 93:22:@14873.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@14913.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_57 ( // @[package.scala 93:22:@14921.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@14929.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_59 ( // @[package.scala 93:22:@14937.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_60 ( // @[package.scala 93:22:@14945.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_61 ( // @[package.scala 93:22:@14953.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_62 ( // @[package.scala 93:22:@14961.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_63 ( // @[package.scala 93:22:@14969.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_64 ( // @[package.scala 93:22:@15009.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_65 ( // @[package.scala 93:22:@15017.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_66 ( // @[package.scala 93:22:@15025.4]
    .clock(RetimeWrapper_66_clock),
    .reset(RetimeWrapper_66_reset),
    .io_flow(RetimeWrapper_66_io_flow),
    .io_in(RetimeWrapper_66_io_in),
    .io_out(RetimeWrapper_66_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_67 ( // @[package.scala 93:22:@15033.4]
    .clock(RetimeWrapper_67_clock),
    .reset(RetimeWrapper_67_reset),
    .io_flow(RetimeWrapper_67_io_flow),
    .io_in(RetimeWrapper_67_io_in),
    .io_out(RetimeWrapper_67_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_68 ( // @[package.scala 93:22:@15041.4]
    .clock(RetimeWrapper_68_clock),
    .reset(RetimeWrapper_68_reset),
    .io_flow(RetimeWrapper_68_io_flow),
    .io_in(RetimeWrapper_68_io_in),
    .io_out(RetimeWrapper_68_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_69 ( // @[package.scala 93:22:@15049.4]
    .clock(RetimeWrapper_69_clock),
    .reset(RetimeWrapper_69_reset),
    .io_flow(RetimeWrapper_69_io_flow),
    .io_in(RetimeWrapper_69_io_in),
    .io_out(RetimeWrapper_69_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_70 ( // @[package.scala 93:22:@15057.4]
    .clock(RetimeWrapper_70_clock),
    .reset(RetimeWrapper_70_reset),
    .io_flow(RetimeWrapper_70_io_flow),
    .io_in(RetimeWrapper_70_io_in),
    .io_out(RetimeWrapper_70_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_71 ( // @[package.scala 93:22:@15065.4]
    .clock(RetimeWrapper_71_clock),
    .reset(RetimeWrapper_71_reset),
    .io_flow(RetimeWrapper_71_io_flow),
    .io_in(RetimeWrapper_71_io_in),
    .io_out(RetimeWrapper_71_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_72 ( // @[package.scala 93:22:@15105.4]
    .clock(RetimeWrapper_72_clock),
    .reset(RetimeWrapper_72_reset),
    .io_flow(RetimeWrapper_72_io_flow),
    .io_in(RetimeWrapper_72_io_in),
    .io_out(RetimeWrapper_72_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_73 ( // @[package.scala 93:22:@15113.4]
    .clock(RetimeWrapper_73_clock),
    .reset(RetimeWrapper_73_reset),
    .io_flow(RetimeWrapper_73_io_flow),
    .io_in(RetimeWrapper_73_io_in),
    .io_out(RetimeWrapper_73_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_74 ( // @[package.scala 93:22:@15121.4]
    .clock(RetimeWrapper_74_clock),
    .reset(RetimeWrapper_74_reset),
    .io_flow(RetimeWrapper_74_io_flow),
    .io_in(RetimeWrapper_74_io_in),
    .io_out(RetimeWrapper_74_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_75 ( // @[package.scala 93:22:@15129.4]
    .clock(RetimeWrapper_75_clock),
    .reset(RetimeWrapper_75_reset),
    .io_flow(RetimeWrapper_75_io_flow),
    .io_in(RetimeWrapper_75_io_in),
    .io_out(RetimeWrapper_75_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_76 ( // @[package.scala 93:22:@15137.4]
    .clock(RetimeWrapper_76_clock),
    .reset(RetimeWrapper_76_reset),
    .io_flow(RetimeWrapper_76_io_flow),
    .io_in(RetimeWrapper_76_io_in),
    .io_out(RetimeWrapper_76_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_77 ( // @[package.scala 93:22:@15145.4]
    .clock(RetimeWrapper_77_clock),
    .reset(RetimeWrapper_77_reset),
    .io_flow(RetimeWrapper_77_io_flow),
    .io_in(RetimeWrapper_77_io_in),
    .io_out(RetimeWrapper_77_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_78 ( // @[package.scala 93:22:@15153.4]
    .clock(RetimeWrapper_78_clock),
    .reset(RetimeWrapper_78_reset),
    .io_flow(RetimeWrapper_78_io_flow),
    .io_in(RetimeWrapper_78_io_in),
    .io_out(RetimeWrapper_78_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_79 ( // @[package.scala 93:22:@15161.4]
    .clock(RetimeWrapper_79_clock),
    .reset(RetimeWrapper_79_reset),
    .io_flow(RetimeWrapper_79_io_flow),
    .io_in(RetimeWrapper_79_io_in),
    .io_out(RetimeWrapper_79_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_80 ( // @[package.scala 93:22:@15201.4]
    .clock(RetimeWrapper_80_clock),
    .reset(RetimeWrapper_80_reset),
    .io_flow(RetimeWrapper_80_io_flow),
    .io_in(RetimeWrapper_80_io_in),
    .io_out(RetimeWrapper_80_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_81 ( // @[package.scala 93:22:@15209.4]
    .clock(RetimeWrapper_81_clock),
    .reset(RetimeWrapper_81_reset),
    .io_flow(RetimeWrapper_81_io_flow),
    .io_in(RetimeWrapper_81_io_in),
    .io_out(RetimeWrapper_81_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_82 ( // @[package.scala 93:22:@15217.4]
    .clock(RetimeWrapper_82_clock),
    .reset(RetimeWrapper_82_reset),
    .io_flow(RetimeWrapper_82_io_flow),
    .io_in(RetimeWrapper_82_io_in),
    .io_out(RetimeWrapper_82_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_83 ( // @[package.scala 93:22:@15225.4]
    .clock(RetimeWrapper_83_clock),
    .reset(RetimeWrapper_83_reset),
    .io_flow(RetimeWrapper_83_io_flow),
    .io_in(RetimeWrapper_83_io_in),
    .io_out(RetimeWrapper_83_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_84 ( // @[package.scala 93:22:@15233.4]
    .clock(RetimeWrapper_84_clock),
    .reset(RetimeWrapper_84_reset),
    .io_flow(RetimeWrapper_84_io_flow),
    .io_in(RetimeWrapper_84_io_in),
    .io_out(RetimeWrapper_84_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_85 ( // @[package.scala 93:22:@15241.4]
    .clock(RetimeWrapper_85_clock),
    .reset(RetimeWrapper_85_reset),
    .io_flow(RetimeWrapper_85_io_flow),
    .io_in(RetimeWrapper_85_io_in),
    .io_out(RetimeWrapper_85_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_86 ( // @[package.scala 93:22:@15249.4]
    .clock(RetimeWrapper_86_clock),
    .reset(RetimeWrapper_86_reset),
    .io_flow(RetimeWrapper_86_io_flow),
    .io_in(RetimeWrapper_86_io_in),
    .io_out(RetimeWrapper_86_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_87 ( // @[package.scala 93:22:@15257.4]
    .clock(RetimeWrapper_87_clock),
    .reset(RetimeWrapper_87_reset),
    .io_flow(RetimeWrapper_87_io_flow),
    .io_in(RetimeWrapper_87_io_in),
    .io_out(RetimeWrapper_87_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_88 ( // @[package.scala 93:22:@15297.4]
    .clock(RetimeWrapper_88_clock),
    .reset(RetimeWrapper_88_reset),
    .io_flow(RetimeWrapper_88_io_flow),
    .io_in(RetimeWrapper_88_io_in),
    .io_out(RetimeWrapper_88_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_89 ( // @[package.scala 93:22:@15305.4]
    .clock(RetimeWrapper_89_clock),
    .reset(RetimeWrapper_89_reset),
    .io_flow(RetimeWrapper_89_io_flow),
    .io_in(RetimeWrapper_89_io_in),
    .io_out(RetimeWrapper_89_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_90 ( // @[package.scala 93:22:@15313.4]
    .clock(RetimeWrapper_90_clock),
    .reset(RetimeWrapper_90_reset),
    .io_flow(RetimeWrapper_90_io_flow),
    .io_in(RetimeWrapper_90_io_in),
    .io_out(RetimeWrapper_90_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_91 ( // @[package.scala 93:22:@15321.4]
    .clock(RetimeWrapper_91_clock),
    .reset(RetimeWrapper_91_reset),
    .io_flow(RetimeWrapper_91_io_flow),
    .io_in(RetimeWrapper_91_io_in),
    .io_out(RetimeWrapper_91_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_92 ( // @[package.scala 93:22:@15329.4]
    .clock(RetimeWrapper_92_clock),
    .reset(RetimeWrapper_92_reset),
    .io_flow(RetimeWrapper_92_io_flow),
    .io_in(RetimeWrapper_92_io_in),
    .io_out(RetimeWrapper_92_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_93 ( // @[package.scala 93:22:@15337.4]
    .clock(RetimeWrapper_93_clock),
    .reset(RetimeWrapper_93_reset),
    .io_flow(RetimeWrapper_93_io_flow),
    .io_in(RetimeWrapper_93_io_in),
    .io_out(RetimeWrapper_93_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_94 ( // @[package.scala 93:22:@15345.4]
    .clock(RetimeWrapper_94_clock),
    .reset(RetimeWrapper_94_reset),
    .io_flow(RetimeWrapper_94_io_flow),
    .io_in(RetimeWrapper_94_io_in),
    .io_out(RetimeWrapper_94_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_95 ( // @[package.scala 93:22:@15353.4]
    .clock(RetimeWrapper_95_clock),
    .reset(RetimeWrapper_95_reset),
    .io_flow(RetimeWrapper_95_io_flow),
    .io_in(RetimeWrapper_95_io_in),
    .io_out(RetimeWrapper_95_io_out)
  );
  assign _T_444 = io_wPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13032.4]
  assign _T_446 = io_wPort_0_banks_1 == 3'h0; // @[MemPrimitives.scala 82:210:@13033.4]
  assign _T_447 = _T_444 & _T_446; // @[MemPrimitives.scala 82:228:@13034.4]
  assign _T_448 = io_wPort_0_en_0 & _T_447; // @[MemPrimitives.scala 83:102:@13035.4]
  assign _T_450 = {_T_448,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13037.4]
  assign _T_455 = io_wPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 82:210:@13044.4]
  assign _T_457 = io_wPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 82:210:@13045.4]
  assign _T_458 = _T_455 & _T_457; // @[MemPrimitives.scala 82:228:@13046.4]
  assign _T_459 = io_wPort_1_en_0 & _T_458; // @[MemPrimitives.scala 83:102:@13047.4]
  assign _T_461 = {_T_459,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13049.4]
  assign _T_468 = io_wPort_0_banks_1 == 3'h2; // @[MemPrimitives.scala 82:210:@13057.4]
  assign _T_469 = _T_444 & _T_468; // @[MemPrimitives.scala 82:228:@13058.4]
  assign _T_470 = io_wPort_0_en_0 & _T_469; // @[MemPrimitives.scala 83:102:@13059.4]
  assign _T_472 = {_T_470,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13061.4]
  assign _T_479 = io_wPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 82:210:@13069.4]
  assign _T_480 = _T_455 & _T_479; // @[MemPrimitives.scala 82:228:@13070.4]
  assign _T_481 = io_wPort_1_en_0 & _T_480; // @[MemPrimitives.scala 83:102:@13071.4]
  assign _T_483 = {_T_481,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13073.4]
  assign _T_488 = io_wPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13080.4]
  assign _T_491 = _T_488 & _T_446; // @[MemPrimitives.scala 82:228:@13082.4]
  assign _T_492 = io_wPort_0_en_0 & _T_491; // @[MemPrimitives.scala 83:102:@13083.4]
  assign _T_494 = {_T_492,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13085.4]
  assign _T_499 = io_wPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 82:210:@13092.4]
  assign _T_502 = _T_499 & _T_457; // @[MemPrimitives.scala 82:228:@13094.4]
  assign _T_503 = io_wPort_1_en_0 & _T_502; // @[MemPrimitives.scala 83:102:@13095.4]
  assign _T_505 = {_T_503,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13097.4]
  assign _T_513 = _T_488 & _T_468; // @[MemPrimitives.scala 82:228:@13106.4]
  assign _T_514 = io_wPort_0_en_0 & _T_513; // @[MemPrimitives.scala 83:102:@13107.4]
  assign _T_516 = {_T_514,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13109.4]
  assign _T_524 = _T_499 & _T_479; // @[MemPrimitives.scala 82:228:@13118.4]
  assign _T_525 = io_wPort_1_en_0 & _T_524; // @[MemPrimitives.scala 83:102:@13119.4]
  assign _T_527 = {_T_525,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13121.4]
  assign _T_532 = io_wPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13128.4]
  assign _T_535 = _T_532 & _T_446; // @[MemPrimitives.scala 82:228:@13130.4]
  assign _T_536 = io_wPort_0_en_0 & _T_535; // @[MemPrimitives.scala 83:102:@13131.4]
  assign _T_538 = {_T_536,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13133.4]
  assign _T_543 = io_wPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 82:210:@13140.4]
  assign _T_546 = _T_543 & _T_457; // @[MemPrimitives.scala 82:228:@13142.4]
  assign _T_547 = io_wPort_1_en_0 & _T_546; // @[MemPrimitives.scala 83:102:@13143.4]
  assign _T_549 = {_T_547,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13145.4]
  assign _T_557 = _T_532 & _T_468; // @[MemPrimitives.scala 82:228:@13154.4]
  assign _T_558 = io_wPort_0_en_0 & _T_557; // @[MemPrimitives.scala 83:102:@13155.4]
  assign _T_560 = {_T_558,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13157.4]
  assign _T_568 = _T_543 & _T_479; // @[MemPrimitives.scala 82:228:@13166.4]
  assign _T_569 = io_wPort_1_en_0 & _T_568; // @[MemPrimitives.scala 83:102:@13167.4]
  assign _T_571 = {_T_569,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13169.4]
  assign _T_576 = io_wPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13176.4]
  assign _T_579 = _T_576 & _T_446; // @[MemPrimitives.scala 82:228:@13178.4]
  assign _T_580 = io_wPort_0_en_0 & _T_579; // @[MemPrimitives.scala 83:102:@13179.4]
  assign _T_582 = {_T_580,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13181.4]
  assign _T_587 = io_wPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 82:210:@13188.4]
  assign _T_590 = _T_587 & _T_457; // @[MemPrimitives.scala 82:228:@13190.4]
  assign _T_591 = io_wPort_1_en_0 & _T_590; // @[MemPrimitives.scala 83:102:@13191.4]
  assign _T_593 = {_T_591,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13193.4]
  assign _T_601 = _T_576 & _T_468; // @[MemPrimitives.scala 82:228:@13202.4]
  assign _T_602 = io_wPort_0_en_0 & _T_601; // @[MemPrimitives.scala 83:102:@13203.4]
  assign _T_604 = {_T_602,io_wPort_0_data_0,io_wPort_0_ofs_0}; // @[Cat.scala 30:58:@13205.4]
  assign _T_612 = _T_587 & _T_479; // @[MemPrimitives.scala 82:228:@13214.4]
  assign _T_613 = io_wPort_1_en_0 & _T_612; // @[MemPrimitives.scala 83:102:@13215.4]
  assign _T_615 = {_T_613,io_wPort_1_data_0,io_wPort_1_ofs_0}; // @[Cat.scala 30:58:@13217.4]
  assign _T_620 = io_rPort_2_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13224.4]
  assign _T_622 = io_rPort_2_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13225.4]
  assign _T_623 = _T_620 & _T_622; // @[MemPrimitives.scala 110:228:@13226.4]
  assign _T_626 = io_rPort_4_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13228.4]
  assign _T_628 = io_rPort_4_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13229.4]
  assign _T_629 = _T_626 & _T_628; // @[MemPrimitives.scala 110:228:@13230.4]
  assign _T_632 = io_rPort_6_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13232.4]
  assign _T_634 = io_rPort_6_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13233.4]
  assign _T_635 = _T_632 & _T_634; // @[MemPrimitives.scala 110:228:@13234.4]
  assign _T_638 = io_rPort_7_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13236.4]
  assign _T_640 = io_rPort_7_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13237.4]
  assign _T_641 = _T_638 & _T_640; // @[MemPrimitives.scala 110:228:@13238.4]
  assign _T_644 = io_rPort_8_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13240.4]
  assign _T_646 = io_rPort_8_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13241.4]
  assign _T_647 = _T_644 & _T_646; // @[MemPrimitives.scala 110:228:@13242.4]
  assign _T_650 = io_rPort_10_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13244.4]
  assign _T_652 = io_rPort_10_banks_1 == 3'h0; // @[MemPrimitives.scala 110:210:@13245.4]
  assign _T_653 = _T_650 & _T_652; // @[MemPrimitives.scala 110:228:@13246.4]
  assign _T_655 = StickySelects_io_outs_0; // @[MemPrimitives.scala 126:35:@13257.4]
  assign _T_656 = StickySelects_io_outs_1; // @[MemPrimitives.scala 126:35:@13258.4]
  assign _T_657 = StickySelects_io_outs_2; // @[MemPrimitives.scala 126:35:@13259.4]
  assign _T_658 = StickySelects_io_outs_3; // @[MemPrimitives.scala 126:35:@13260.4]
  assign _T_659 = StickySelects_io_outs_4; // @[MemPrimitives.scala 126:35:@13261.4]
  assign _T_660 = StickySelects_io_outs_5; // @[MemPrimitives.scala 126:35:@13262.4]
  assign _T_662 = {_T_655,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13264.4]
  assign _T_664 = {_T_656,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13266.4]
  assign _T_666 = {_T_657,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13268.4]
  assign _T_668 = {_T_658,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13270.4]
  assign _T_670 = {_T_659,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13272.4]
  assign _T_672 = {_T_660,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13274.4]
  assign _T_673 = _T_659 ? _T_670 : _T_672; // @[Mux.scala 31:69:@13275.4]
  assign _T_674 = _T_658 ? _T_668 : _T_673; // @[Mux.scala 31:69:@13276.4]
  assign _T_675 = _T_657 ? _T_666 : _T_674; // @[Mux.scala 31:69:@13277.4]
  assign _T_676 = _T_656 ? _T_664 : _T_675; // @[Mux.scala 31:69:@13278.4]
  assign _T_677 = _T_655 ? _T_662 : _T_676; // @[Mux.scala 31:69:@13279.4]
  assign _T_682 = io_rPort_0_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13286.4]
  assign _T_684 = io_rPort_0_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13287.4]
  assign _T_685 = _T_682 & _T_684; // @[MemPrimitives.scala 110:228:@13288.4]
  assign _T_688 = io_rPort_1_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13290.4]
  assign _T_690 = io_rPort_1_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13291.4]
  assign _T_691 = _T_688 & _T_690; // @[MemPrimitives.scala 110:228:@13292.4]
  assign _T_694 = io_rPort_3_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13294.4]
  assign _T_696 = io_rPort_3_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13295.4]
  assign _T_697 = _T_694 & _T_696; // @[MemPrimitives.scala 110:228:@13296.4]
  assign _T_700 = io_rPort_5_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13298.4]
  assign _T_702 = io_rPort_5_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13299.4]
  assign _T_703 = _T_700 & _T_702; // @[MemPrimitives.scala 110:228:@13300.4]
  assign _T_706 = io_rPort_9_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13302.4]
  assign _T_708 = io_rPort_9_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13303.4]
  assign _T_709 = _T_706 & _T_708; // @[MemPrimitives.scala 110:228:@13304.4]
  assign _T_712 = io_rPort_11_banks_0 == 3'h0; // @[MemPrimitives.scala 110:210:@13306.4]
  assign _T_714 = io_rPort_11_banks_1 == 3'h1; // @[MemPrimitives.scala 110:210:@13307.4]
  assign _T_715 = _T_712 & _T_714; // @[MemPrimitives.scala 110:228:@13308.4]
  assign _T_717 = StickySelects_1_io_outs_0; // @[MemPrimitives.scala 126:35:@13319.4]
  assign _T_718 = StickySelects_1_io_outs_1; // @[MemPrimitives.scala 126:35:@13320.4]
  assign _T_719 = StickySelects_1_io_outs_2; // @[MemPrimitives.scala 126:35:@13321.4]
  assign _T_720 = StickySelects_1_io_outs_3; // @[MemPrimitives.scala 126:35:@13322.4]
  assign _T_721 = StickySelects_1_io_outs_4; // @[MemPrimitives.scala 126:35:@13323.4]
  assign _T_722 = StickySelects_1_io_outs_5; // @[MemPrimitives.scala 126:35:@13324.4]
  assign _T_724 = {_T_717,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13326.4]
  assign _T_726 = {_T_718,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13328.4]
  assign _T_728 = {_T_719,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13330.4]
  assign _T_730 = {_T_720,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13332.4]
  assign _T_732 = {_T_721,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13334.4]
  assign _T_734 = {_T_722,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13336.4]
  assign _T_735 = _T_721 ? _T_732 : _T_734; // @[Mux.scala 31:69:@13337.4]
  assign _T_736 = _T_720 ? _T_730 : _T_735; // @[Mux.scala 31:69:@13338.4]
  assign _T_737 = _T_719 ? _T_728 : _T_736; // @[Mux.scala 31:69:@13339.4]
  assign _T_738 = _T_718 ? _T_726 : _T_737; // @[Mux.scala 31:69:@13340.4]
  assign _T_739 = _T_717 ? _T_724 : _T_738; // @[Mux.scala 31:69:@13341.4]
  assign _T_746 = io_rPort_2_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13349.4]
  assign _T_747 = _T_620 & _T_746; // @[MemPrimitives.scala 110:228:@13350.4]
  assign _T_752 = io_rPort_4_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13353.4]
  assign _T_753 = _T_626 & _T_752; // @[MemPrimitives.scala 110:228:@13354.4]
  assign _T_758 = io_rPort_6_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13357.4]
  assign _T_759 = _T_632 & _T_758; // @[MemPrimitives.scala 110:228:@13358.4]
  assign _T_764 = io_rPort_7_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13361.4]
  assign _T_765 = _T_638 & _T_764; // @[MemPrimitives.scala 110:228:@13362.4]
  assign _T_770 = io_rPort_8_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13365.4]
  assign _T_771 = _T_644 & _T_770; // @[MemPrimitives.scala 110:228:@13366.4]
  assign _T_776 = io_rPort_10_banks_1 == 3'h2; // @[MemPrimitives.scala 110:210:@13369.4]
  assign _T_777 = _T_650 & _T_776; // @[MemPrimitives.scala 110:228:@13370.4]
  assign _T_779 = StickySelects_2_io_outs_0; // @[MemPrimitives.scala 126:35:@13381.4]
  assign _T_780 = StickySelects_2_io_outs_1; // @[MemPrimitives.scala 126:35:@13382.4]
  assign _T_781 = StickySelects_2_io_outs_2; // @[MemPrimitives.scala 126:35:@13383.4]
  assign _T_782 = StickySelects_2_io_outs_3; // @[MemPrimitives.scala 126:35:@13384.4]
  assign _T_783 = StickySelects_2_io_outs_4; // @[MemPrimitives.scala 126:35:@13385.4]
  assign _T_784 = StickySelects_2_io_outs_5; // @[MemPrimitives.scala 126:35:@13386.4]
  assign _T_786 = {_T_779,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13388.4]
  assign _T_788 = {_T_780,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13390.4]
  assign _T_790 = {_T_781,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13392.4]
  assign _T_792 = {_T_782,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13394.4]
  assign _T_794 = {_T_783,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13396.4]
  assign _T_796 = {_T_784,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13398.4]
  assign _T_797 = _T_783 ? _T_794 : _T_796; // @[Mux.scala 31:69:@13399.4]
  assign _T_798 = _T_782 ? _T_792 : _T_797; // @[Mux.scala 31:69:@13400.4]
  assign _T_799 = _T_781 ? _T_790 : _T_798; // @[Mux.scala 31:69:@13401.4]
  assign _T_800 = _T_780 ? _T_788 : _T_799; // @[Mux.scala 31:69:@13402.4]
  assign _T_801 = _T_779 ? _T_786 : _T_800; // @[Mux.scala 31:69:@13403.4]
  assign _T_808 = io_rPort_0_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13411.4]
  assign _T_809 = _T_682 & _T_808; // @[MemPrimitives.scala 110:228:@13412.4]
  assign _T_814 = io_rPort_1_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13415.4]
  assign _T_815 = _T_688 & _T_814; // @[MemPrimitives.scala 110:228:@13416.4]
  assign _T_820 = io_rPort_3_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13419.4]
  assign _T_821 = _T_694 & _T_820; // @[MemPrimitives.scala 110:228:@13420.4]
  assign _T_826 = io_rPort_5_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13423.4]
  assign _T_827 = _T_700 & _T_826; // @[MemPrimitives.scala 110:228:@13424.4]
  assign _T_832 = io_rPort_9_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13427.4]
  assign _T_833 = _T_706 & _T_832; // @[MemPrimitives.scala 110:228:@13428.4]
  assign _T_838 = io_rPort_11_banks_1 == 3'h3; // @[MemPrimitives.scala 110:210:@13431.4]
  assign _T_839 = _T_712 & _T_838; // @[MemPrimitives.scala 110:228:@13432.4]
  assign _T_841 = StickySelects_3_io_outs_0; // @[MemPrimitives.scala 126:35:@13443.4]
  assign _T_842 = StickySelects_3_io_outs_1; // @[MemPrimitives.scala 126:35:@13444.4]
  assign _T_843 = StickySelects_3_io_outs_2; // @[MemPrimitives.scala 126:35:@13445.4]
  assign _T_844 = StickySelects_3_io_outs_3; // @[MemPrimitives.scala 126:35:@13446.4]
  assign _T_845 = StickySelects_3_io_outs_4; // @[MemPrimitives.scala 126:35:@13447.4]
  assign _T_846 = StickySelects_3_io_outs_5; // @[MemPrimitives.scala 126:35:@13448.4]
  assign _T_848 = {_T_841,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13450.4]
  assign _T_850 = {_T_842,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13452.4]
  assign _T_852 = {_T_843,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13454.4]
  assign _T_854 = {_T_844,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13456.4]
  assign _T_856 = {_T_845,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13458.4]
  assign _T_858 = {_T_846,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13460.4]
  assign _T_859 = _T_845 ? _T_856 : _T_858; // @[Mux.scala 31:69:@13461.4]
  assign _T_860 = _T_844 ? _T_854 : _T_859; // @[Mux.scala 31:69:@13462.4]
  assign _T_861 = _T_843 ? _T_852 : _T_860; // @[Mux.scala 31:69:@13463.4]
  assign _T_862 = _T_842 ? _T_850 : _T_861; // @[Mux.scala 31:69:@13464.4]
  assign _T_863 = _T_841 ? _T_848 : _T_862; // @[Mux.scala 31:69:@13465.4]
  assign _T_868 = io_rPort_2_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13472.4]
  assign _T_871 = _T_868 & _T_622; // @[MemPrimitives.scala 110:228:@13474.4]
  assign _T_874 = io_rPort_4_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13476.4]
  assign _T_877 = _T_874 & _T_628; // @[MemPrimitives.scala 110:228:@13478.4]
  assign _T_880 = io_rPort_6_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13480.4]
  assign _T_883 = _T_880 & _T_634; // @[MemPrimitives.scala 110:228:@13482.4]
  assign _T_886 = io_rPort_7_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13484.4]
  assign _T_889 = _T_886 & _T_640; // @[MemPrimitives.scala 110:228:@13486.4]
  assign _T_892 = io_rPort_8_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13488.4]
  assign _T_895 = _T_892 & _T_646; // @[MemPrimitives.scala 110:228:@13490.4]
  assign _T_898 = io_rPort_10_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13492.4]
  assign _T_901 = _T_898 & _T_652; // @[MemPrimitives.scala 110:228:@13494.4]
  assign _T_903 = StickySelects_4_io_outs_0; // @[MemPrimitives.scala 126:35:@13505.4]
  assign _T_904 = StickySelects_4_io_outs_1; // @[MemPrimitives.scala 126:35:@13506.4]
  assign _T_905 = StickySelects_4_io_outs_2; // @[MemPrimitives.scala 126:35:@13507.4]
  assign _T_906 = StickySelects_4_io_outs_3; // @[MemPrimitives.scala 126:35:@13508.4]
  assign _T_907 = StickySelects_4_io_outs_4; // @[MemPrimitives.scala 126:35:@13509.4]
  assign _T_908 = StickySelects_4_io_outs_5; // @[MemPrimitives.scala 126:35:@13510.4]
  assign _T_910 = {_T_903,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13512.4]
  assign _T_912 = {_T_904,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13514.4]
  assign _T_914 = {_T_905,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13516.4]
  assign _T_916 = {_T_906,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13518.4]
  assign _T_918 = {_T_907,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13520.4]
  assign _T_920 = {_T_908,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13522.4]
  assign _T_921 = _T_907 ? _T_918 : _T_920; // @[Mux.scala 31:69:@13523.4]
  assign _T_922 = _T_906 ? _T_916 : _T_921; // @[Mux.scala 31:69:@13524.4]
  assign _T_923 = _T_905 ? _T_914 : _T_922; // @[Mux.scala 31:69:@13525.4]
  assign _T_924 = _T_904 ? _T_912 : _T_923; // @[Mux.scala 31:69:@13526.4]
  assign _T_925 = _T_903 ? _T_910 : _T_924; // @[Mux.scala 31:69:@13527.4]
  assign _T_930 = io_rPort_0_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13534.4]
  assign _T_933 = _T_930 & _T_684; // @[MemPrimitives.scala 110:228:@13536.4]
  assign _T_936 = io_rPort_1_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13538.4]
  assign _T_939 = _T_936 & _T_690; // @[MemPrimitives.scala 110:228:@13540.4]
  assign _T_942 = io_rPort_3_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13542.4]
  assign _T_945 = _T_942 & _T_696; // @[MemPrimitives.scala 110:228:@13544.4]
  assign _T_948 = io_rPort_5_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13546.4]
  assign _T_951 = _T_948 & _T_702; // @[MemPrimitives.scala 110:228:@13548.4]
  assign _T_954 = io_rPort_9_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13550.4]
  assign _T_957 = _T_954 & _T_708; // @[MemPrimitives.scala 110:228:@13552.4]
  assign _T_960 = io_rPort_11_banks_0 == 3'h1; // @[MemPrimitives.scala 110:210:@13554.4]
  assign _T_963 = _T_960 & _T_714; // @[MemPrimitives.scala 110:228:@13556.4]
  assign _T_965 = StickySelects_5_io_outs_0; // @[MemPrimitives.scala 126:35:@13567.4]
  assign _T_966 = StickySelects_5_io_outs_1; // @[MemPrimitives.scala 126:35:@13568.4]
  assign _T_967 = StickySelects_5_io_outs_2; // @[MemPrimitives.scala 126:35:@13569.4]
  assign _T_968 = StickySelects_5_io_outs_3; // @[MemPrimitives.scala 126:35:@13570.4]
  assign _T_969 = StickySelects_5_io_outs_4; // @[MemPrimitives.scala 126:35:@13571.4]
  assign _T_970 = StickySelects_5_io_outs_5; // @[MemPrimitives.scala 126:35:@13572.4]
  assign _T_972 = {_T_965,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13574.4]
  assign _T_974 = {_T_966,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13576.4]
  assign _T_976 = {_T_967,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13578.4]
  assign _T_978 = {_T_968,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13580.4]
  assign _T_980 = {_T_969,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13582.4]
  assign _T_982 = {_T_970,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13584.4]
  assign _T_983 = _T_969 ? _T_980 : _T_982; // @[Mux.scala 31:69:@13585.4]
  assign _T_984 = _T_968 ? _T_978 : _T_983; // @[Mux.scala 31:69:@13586.4]
  assign _T_985 = _T_967 ? _T_976 : _T_984; // @[Mux.scala 31:69:@13587.4]
  assign _T_986 = _T_966 ? _T_974 : _T_985; // @[Mux.scala 31:69:@13588.4]
  assign _T_987 = _T_965 ? _T_972 : _T_986; // @[Mux.scala 31:69:@13589.4]
  assign _T_995 = _T_868 & _T_746; // @[MemPrimitives.scala 110:228:@13598.4]
  assign _T_1001 = _T_874 & _T_752; // @[MemPrimitives.scala 110:228:@13602.4]
  assign _T_1007 = _T_880 & _T_758; // @[MemPrimitives.scala 110:228:@13606.4]
  assign _T_1013 = _T_886 & _T_764; // @[MemPrimitives.scala 110:228:@13610.4]
  assign _T_1019 = _T_892 & _T_770; // @[MemPrimitives.scala 110:228:@13614.4]
  assign _T_1025 = _T_898 & _T_776; // @[MemPrimitives.scala 110:228:@13618.4]
  assign _T_1027 = StickySelects_6_io_outs_0; // @[MemPrimitives.scala 126:35:@13629.4]
  assign _T_1028 = StickySelects_6_io_outs_1; // @[MemPrimitives.scala 126:35:@13630.4]
  assign _T_1029 = StickySelects_6_io_outs_2; // @[MemPrimitives.scala 126:35:@13631.4]
  assign _T_1030 = StickySelects_6_io_outs_3; // @[MemPrimitives.scala 126:35:@13632.4]
  assign _T_1031 = StickySelects_6_io_outs_4; // @[MemPrimitives.scala 126:35:@13633.4]
  assign _T_1032 = StickySelects_6_io_outs_5; // @[MemPrimitives.scala 126:35:@13634.4]
  assign _T_1034 = {_T_1027,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13636.4]
  assign _T_1036 = {_T_1028,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13638.4]
  assign _T_1038 = {_T_1029,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13640.4]
  assign _T_1040 = {_T_1030,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13642.4]
  assign _T_1042 = {_T_1031,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13644.4]
  assign _T_1044 = {_T_1032,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13646.4]
  assign _T_1045 = _T_1031 ? _T_1042 : _T_1044; // @[Mux.scala 31:69:@13647.4]
  assign _T_1046 = _T_1030 ? _T_1040 : _T_1045; // @[Mux.scala 31:69:@13648.4]
  assign _T_1047 = _T_1029 ? _T_1038 : _T_1046; // @[Mux.scala 31:69:@13649.4]
  assign _T_1048 = _T_1028 ? _T_1036 : _T_1047; // @[Mux.scala 31:69:@13650.4]
  assign _T_1049 = _T_1027 ? _T_1034 : _T_1048; // @[Mux.scala 31:69:@13651.4]
  assign _T_1057 = _T_930 & _T_808; // @[MemPrimitives.scala 110:228:@13660.4]
  assign _T_1063 = _T_936 & _T_814; // @[MemPrimitives.scala 110:228:@13664.4]
  assign _T_1069 = _T_942 & _T_820; // @[MemPrimitives.scala 110:228:@13668.4]
  assign _T_1075 = _T_948 & _T_826; // @[MemPrimitives.scala 110:228:@13672.4]
  assign _T_1081 = _T_954 & _T_832; // @[MemPrimitives.scala 110:228:@13676.4]
  assign _T_1087 = _T_960 & _T_838; // @[MemPrimitives.scala 110:228:@13680.4]
  assign _T_1089 = StickySelects_7_io_outs_0; // @[MemPrimitives.scala 126:35:@13691.4]
  assign _T_1090 = StickySelects_7_io_outs_1; // @[MemPrimitives.scala 126:35:@13692.4]
  assign _T_1091 = StickySelects_7_io_outs_2; // @[MemPrimitives.scala 126:35:@13693.4]
  assign _T_1092 = StickySelects_7_io_outs_3; // @[MemPrimitives.scala 126:35:@13694.4]
  assign _T_1093 = StickySelects_7_io_outs_4; // @[MemPrimitives.scala 126:35:@13695.4]
  assign _T_1094 = StickySelects_7_io_outs_5; // @[MemPrimitives.scala 126:35:@13696.4]
  assign _T_1096 = {_T_1089,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13698.4]
  assign _T_1098 = {_T_1090,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13700.4]
  assign _T_1100 = {_T_1091,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13702.4]
  assign _T_1102 = {_T_1092,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13704.4]
  assign _T_1104 = {_T_1093,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13706.4]
  assign _T_1106 = {_T_1094,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13708.4]
  assign _T_1107 = _T_1093 ? _T_1104 : _T_1106; // @[Mux.scala 31:69:@13709.4]
  assign _T_1108 = _T_1092 ? _T_1102 : _T_1107; // @[Mux.scala 31:69:@13710.4]
  assign _T_1109 = _T_1091 ? _T_1100 : _T_1108; // @[Mux.scala 31:69:@13711.4]
  assign _T_1110 = _T_1090 ? _T_1098 : _T_1109; // @[Mux.scala 31:69:@13712.4]
  assign _T_1111 = _T_1089 ? _T_1096 : _T_1110; // @[Mux.scala 31:69:@13713.4]
  assign _T_1116 = io_rPort_2_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13720.4]
  assign _T_1119 = _T_1116 & _T_622; // @[MemPrimitives.scala 110:228:@13722.4]
  assign _T_1122 = io_rPort_4_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13724.4]
  assign _T_1125 = _T_1122 & _T_628; // @[MemPrimitives.scala 110:228:@13726.4]
  assign _T_1128 = io_rPort_6_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13728.4]
  assign _T_1131 = _T_1128 & _T_634; // @[MemPrimitives.scala 110:228:@13730.4]
  assign _T_1134 = io_rPort_7_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13732.4]
  assign _T_1137 = _T_1134 & _T_640; // @[MemPrimitives.scala 110:228:@13734.4]
  assign _T_1140 = io_rPort_8_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13736.4]
  assign _T_1143 = _T_1140 & _T_646; // @[MemPrimitives.scala 110:228:@13738.4]
  assign _T_1146 = io_rPort_10_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13740.4]
  assign _T_1149 = _T_1146 & _T_652; // @[MemPrimitives.scala 110:228:@13742.4]
  assign _T_1151 = StickySelects_8_io_outs_0; // @[MemPrimitives.scala 126:35:@13753.4]
  assign _T_1152 = StickySelects_8_io_outs_1; // @[MemPrimitives.scala 126:35:@13754.4]
  assign _T_1153 = StickySelects_8_io_outs_2; // @[MemPrimitives.scala 126:35:@13755.4]
  assign _T_1154 = StickySelects_8_io_outs_3; // @[MemPrimitives.scala 126:35:@13756.4]
  assign _T_1155 = StickySelects_8_io_outs_4; // @[MemPrimitives.scala 126:35:@13757.4]
  assign _T_1156 = StickySelects_8_io_outs_5; // @[MemPrimitives.scala 126:35:@13758.4]
  assign _T_1158 = {_T_1151,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13760.4]
  assign _T_1160 = {_T_1152,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13762.4]
  assign _T_1162 = {_T_1153,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13764.4]
  assign _T_1164 = {_T_1154,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13766.4]
  assign _T_1166 = {_T_1155,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13768.4]
  assign _T_1168 = {_T_1156,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13770.4]
  assign _T_1169 = _T_1155 ? _T_1166 : _T_1168; // @[Mux.scala 31:69:@13771.4]
  assign _T_1170 = _T_1154 ? _T_1164 : _T_1169; // @[Mux.scala 31:69:@13772.4]
  assign _T_1171 = _T_1153 ? _T_1162 : _T_1170; // @[Mux.scala 31:69:@13773.4]
  assign _T_1172 = _T_1152 ? _T_1160 : _T_1171; // @[Mux.scala 31:69:@13774.4]
  assign _T_1173 = _T_1151 ? _T_1158 : _T_1172; // @[Mux.scala 31:69:@13775.4]
  assign _T_1178 = io_rPort_0_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13782.4]
  assign _T_1181 = _T_1178 & _T_684; // @[MemPrimitives.scala 110:228:@13784.4]
  assign _T_1184 = io_rPort_1_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13786.4]
  assign _T_1187 = _T_1184 & _T_690; // @[MemPrimitives.scala 110:228:@13788.4]
  assign _T_1190 = io_rPort_3_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13790.4]
  assign _T_1193 = _T_1190 & _T_696; // @[MemPrimitives.scala 110:228:@13792.4]
  assign _T_1196 = io_rPort_5_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13794.4]
  assign _T_1199 = _T_1196 & _T_702; // @[MemPrimitives.scala 110:228:@13796.4]
  assign _T_1202 = io_rPort_9_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13798.4]
  assign _T_1205 = _T_1202 & _T_708; // @[MemPrimitives.scala 110:228:@13800.4]
  assign _T_1208 = io_rPort_11_banks_0 == 3'h2; // @[MemPrimitives.scala 110:210:@13802.4]
  assign _T_1211 = _T_1208 & _T_714; // @[MemPrimitives.scala 110:228:@13804.4]
  assign _T_1213 = StickySelects_9_io_outs_0; // @[MemPrimitives.scala 126:35:@13815.4]
  assign _T_1214 = StickySelects_9_io_outs_1; // @[MemPrimitives.scala 126:35:@13816.4]
  assign _T_1215 = StickySelects_9_io_outs_2; // @[MemPrimitives.scala 126:35:@13817.4]
  assign _T_1216 = StickySelects_9_io_outs_3; // @[MemPrimitives.scala 126:35:@13818.4]
  assign _T_1217 = StickySelects_9_io_outs_4; // @[MemPrimitives.scala 126:35:@13819.4]
  assign _T_1218 = StickySelects_9_io_outs_5; // @[MemPrimitives.scala 126:35:@13820.4]
  assign _T_1220 = {_T_1213,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13822.4]
  assign _T_1222 = {_T_1214,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13824.4]
  assign _T_1224 = {_T_1215,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13826.4]
  assign _T_1226 = {_T_1216,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13828.4]
  assign _T_1228 = {_T_1217,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13830.4]
  assign _T_1230 = {_T_1218,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13832.4]
  assign _T_1231 = _T_1217 ? _T_1228 : _T_1230; // @[Mux.scala 31:69:@13833.4]
  assign _T_1232 = _T_1216 ? _T_1226 : _T_1231; // @[Mux.scala 31:69:@13834.4]
  assign _T_1233 = _T_1215 ? _T_1224 : _T_1232; // @[Mux.scala 31:69:@13835.4]
  assign _T_1234 = _T_1214 ? _T_1222 : _T_1233; // @[Mux.scala 31:69:@13836.4]
  assign _T_1235 = _T_1213 ? _T_1220 : _T_1234; // @[Mux.scala 31:69:@13837.4]
  assign _T_1243 = _T_1116 & _T_746; // @[MemPrimitives.scala 110:228:@13846.4]
  assign _T_1249 = _T_1122 & _T_752; // @[MemPrimitives.scala 110:228:@13850.4]
  assign _T_1255 = _T_1128 & _T_758; // @[MemPrimitives.scala 110:228:@13854.4]
  assign _T_1261 = _T_1134 & _T_764; // @[MemPrimitives.scala 110:228:@13858.4]
  assign _T_1267 = _T_1140 & _T_770; // @[MemPrimitives.scala 110:228:@13862.4]
  assign _T_1273 = _T_1146 & _T_776; // @[MemPrimitives.scala 110:228:@13866.4]
  assign _T_1275 = StickySelects_10_io_outs_0; // @[MemPrimitives.scala 126:35:@13877.4]
  assign _T_1276 = StickySelects_10_io_outs_1; // @[MemPrimitives.scala 126:35:@13878.4]
  assign _T_1277 = StickySelects_10_io_outs_2; // @[MemPrimitives.scala 126:35:@13879.4]
  assign _T_1278 = StickySelects_10_io_outs_3; // @[MemPrimitives.scala 126:35:@13880.4]
  assign _T_1279 = StickySelects_10_io_outs_4; // @[MemPrimitives.scala 126:35:@13881.4]
  assign _T_1280 = StickySelects_10_io_outs_5; // @[MemPrimitives.scala 126:35:@13882.4]
  assign _T_1282 = {_T_1275,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@13884.4]
  assign _T_1284 = {_T_1276,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@13886.4]
  assign _T_1286 = {_T_1277,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@13888.4]
  assign _T_1288 = {_T_1278,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@13890.4]
  assign _T_1290 = {_T_1279,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@13892.4]
  assign _T_1292 = {_T_1280,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@13894.4]
  assign _T_1293 = _T_1279 ? _T_1290 : _T_1292; // @[Mux.scala 31:69:@13895.4]
  assign _T_1294 = _T_1278 ? _T_1288 : _T_1293; // @[Mux.scala 31:69:@13896.4]
  assign _T_1295 = _T_1277 ? _T_1286 : _T_1294; // @[Mux.scala 31:69:@13897.4]
  assign _T_1296 = _T_1276 ? _T_1284 : _T_1295; // @[Mux.scala 31:69:@13898.4]
  assign _T_1297 = _T_1275 ? _T_1282 : _T_1296; // @[Mux.scala 31:69:@13899.4]
  assign _T_1305 = _T_1178 & _T_808; // @[MemPrimitives.scala 110:228:@13908.4]
  assign _T_1311 = _T_1184 & _T_814; // @[MemPrimitives.scala 110:228:@13912.4]
  assign _T_1317 = _T_1190 & _T_820; // @[MemPrimitives.scala 110:228:@13916.4]
  assign _T_1323 = _T_1196 & _T_826; // @[MemPrimitives.scala 110:228:@13920.4]
  assign _T_1329 = _T_1202 & _T_832; // @[MemPrimitives.scala 110:228:@13924.4]
  assign _T_1335 = _T_1208 & _T_838; // @[MemPrimitives.scala 110:228:@13928.4]
  assign _T_1337 = StickySelects_11_io_outs_0; // @[MemPrimitives.scala 126:35:@13939.4]
  assign _T_1338 = StickySelects_11_io_outs_1; // @[MemPrimitives.scala 126:35:@13940.4]
  assign _T_1339 = StickySelects_11_io_outs_2; // @[MemPrimitives.scala 126:35:@13941.4]
  assign _T_1340 = StickySelects_11_io_outs_3; // @[MemPrimitives.scala 126:35:@13942.4]
  assign _T_1341 = StickySelects_11_io_outs_4; // @[MemPrimitives.scala 126:35:@13943.4]
  assign _T_1342 = StickySelects_11_io_outs_5; // @[MemPrimitives.scala 126:35:@13944.4]
  assign _T_1344 = {_T_1337,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@13946.4]
  assign _T_1346 = {_T_1338,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@13948.4]
  assign _T_1348 = {_T_1339,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@13950.4]
  assign _T_1350 = {_T_1340,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@13952.4]
  assign _T_1352 = {_T_1341,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@13954.4]
  assign _T_1354 = {_T_1342,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@13956.4]
  assign _T_1355 = _T_1341 ? _T_1352 : _T_1354; // @[Mux.scala 31:69:@13957.4]
  assign _T_1356 = _T_1340 ? _T_1350 : _T_1355; // @[Mux.scala 31:69:@13958.4]
  assign _T_1357 = _T_1339 ? _T_1348 : _T_1356; // @[Mux.scala 31:69:@13959.4]
  assign _T_1358 = _T_1338 ? _T_1346 : _T_1357; // @[Mux.scala 31:69:@13960.4]
  assign _T_1359 = _T_1337 ? _T_1344 : _T_1358; // @[Mux.scala 31:69:@13961.4]
  assign _T_1364 = io_rPort_2_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13968.4]
  assign _T_1367 = _T_1364 & _T_622; // @[MemPrimitives.scala 110:228:@13970.4]
  assign _T_1370 = io_rPort_4_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13972.4]
  assign _T_1373 = _T_1370 & _T_628; // @[MemPrimitives.scala 110:228:@13974.4]
  assign _T_1376 = io_rPort_6_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13976.4]
  assign _T_1379 = _T_1376 & _T_634; // @[MemPrimitives.scala 110:228:@13978.4]
  assign _T_1382 = io_rPort_7_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13980.4]
  assign _T_1385 = _T_1382 & _T_640; // @[MemPrimitives.scala 110:228:@13982.4]
  assign _T_1388 = io_rPort_8_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13984.4]
  assign _T_1391 = _T_1388 & _T_646; // @[MemPrimitives.scala 110:228:@13986.4]
  assign _T_1394 = io_rPort_10_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@13988.4]
  assign _T_1397 = _T_1394 & _T_652; // @[MemPrimitives.scala 110:228:@13990.4]
  assign _T_1399 = StickySelects_12_io_outs_0; // @[MemPrimitives.scala 126:35:@14001.4]
  assign _T_1400 = StickySelects_12_io_outs_1; // @[MemPrimitives.scala 126:35:@14002.4]
  assign _T_1401 = StickySelects_12_io_outs_2; // @[MemPrimitives.scala 126:35:@14003.4]
  assign _T_1402 = StickySelects_12_io_outs_3; // @[MemPrimitives.scala 126:35:@14004.4]
  assign _T_1403 = StickySelects_12_io_outs_4; // @[MemPrimitives.scala 126:35:@14005.4]
  assign _T_1404 = StickySelects_12_io_outs_5; // @[MemPrimitives.scala 126:35:@14006.4]
  assign _T_1406 = {_T_1399,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14008.4]
  assign _T_1408 = {_T_1400,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14010.4]
  assign _T_1410 = {_T_1401,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14012.4]
  assign _T_1412 = {_T_1402,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14014.4]
  assign _T_1414 = {_T_1403,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14016.4]
  assign _T_1416 = {_T_1404,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@14018.4]
  assign _T_1417 = _T_1403 ? _T_1414 : _T_1416; // @[Mux.scala 31:69:@14019.4]
  assign _T_1418 = _T_1402 ? _T_1412 : _T_1417; // @[Mux.scala 31:69:@14020.4]
  assign _T_1419 = _T_1401 ? _T_1410 : _T_1418; // @[Mux.scala 31:69:@14021.4]
  assign _T_1420 = _T_1400 ? _T_1408 : _T_1419; // @[Mux.scala 31:69:@14022.4]
  assign _T_1421 = _T_1399 ? _T_1406 : _T_1420; // @[Mux.scala 31:69:@14023.4]
  assign _T_1426 = io_rPort_0_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14030.4]
  assign _T_1429 = _T_1426 & _T_684; // @[MemPrimitives.scala 110:228:@14032.4]
  assign _T_1432 = io_rPort_1_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14034.4]
  assign _T_1435 = _T_1432 & _T_690; // @[MemPrimitives.scala 110:228:@14036.4]
  assign _T_1438 = io_rPort_3_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14038.4]
  assign _T_1441 = _T_1438 & _T_696; // @[MemPrimitives.scala 110:228:@14040.4]
  assign _T_1444 = io_rPort_5_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14042.4]
  assign _T_1447 = _T_1444 & _T_702; // @[MemPrimitives.scala 110:228:@14044.4]
  assign _T_1450 = io_rPort_9_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14046.4]
  assign _T_1453 = _T_1450 & _T_708; // @[MemPrimitives.scala 110:228:@14048.4]
  assign _T_1456 = io_rPort_11_banks_0 == 3'h3; // @[MemPrimitives.scala 110:210:@14050.4]
  assign _T_1459 = _T_1456 & _T_714; // @[MemPrimitives.scala 110:228:@14052.4]
  assign _T_1461 = StickySelects_13_io_outs_0; // @[MemPrimitives.scala 126:35:@14063.4]
  assign _T_1462 = StickySelects_13_io_outs_1; // @[MemPrimitives.scala 126:35:@14064.4]
  assign _T_1463 = StickySelects_13_io_outs_2; // @[MemPrimitives.scala 126:35:@14065.4]
  assign _T_1464 = StickySelects_13_io_outs_3; // @[MemPrimitives.scala 126:35:@14066.4]
  assign _T_1465 = StickySelects_13_io_outs_4; // @[MemPrimitives.scala 126:35:@14067.4]
  assign _T_1466 = StickySelects_13_io_outs_5; // @[MemPrimitives.scala 126:35:@14068.4]
  assign _T_1468 = {_T_1461,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14070.4]
  assign _T_1470 = {_T_1462,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14072.4]
  assign _T_1472 = {_T_1463,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14074.4]
  assign _T_1474 = {_T_1464,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14076.4]
  assign _T_1476 = {_T_1465,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14078.4]
  assign _T_1478 = {_T_1466,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@14080.4]
  assign _T_1479 = _T_1465 ? _T_1476 : _T_1478; // @[Mux.scala 31:69:@14081.4]
  assign _T_1480 = _T_1464 ? _T_1474 : _T_1479; // @[Mux.scala 31:69:@14082.4]
  assign _T_1481 = _T_1463 ? _T_1472 : _T_1480; // @[Mux.scala 31:69:@14083.4]
  assign _T_1482 = _T_1462 ? _T_1470 : _T_1481; // @[Mux.scala 31:69:@14084.4]
  assign _T_1483 = _T_1461 ? _T_1468 : _T_1482; // @[Mux.scala 31:69:@14085.4]
  assign _T_1491 = _T_1364 & _T_746; // @[MemPrimitives.scala 110:228:@14094.4]
  assign _T_1497 = _T_1370 & _T_752; // @[MemPrimitives.scala 110:228:@14098.4]
  assign _T_1503 = _T_1376 & _T_758; // @[MemPrimitives.scala 110:228:@14102.4]
  assign _T_1509 = _T_1382 & _T_764; // @[MemPrimitives.scala 110:228:@14106.4]
  assign _T_1515 = _T_1388 & _T_770; // @[MemPrimitives.scala 110:228:@14110.4]
  assign _T_1521 = _T_1394 & _T_776; // @[MemPrimitives.scala 110:228:@14114.4]
  assign _T_1523 = StickySelects_14_io_outs_0; // @[MemPrimitives.scala 126:35:@14125.4]
  assign _T_1524 = StickySelects_14_io_outs_1; // @[MemPrimitives.scala 126:35:@14126.4]
  assign _T_1525 = StickySelects_14_io_outs_2; // @[MemPrimitives.scala 126:35:@14127.4]
  assign _T_1526 = StickySelects_14_io_outs_3; // @[MemPrimitives.scala 126:35:@14128.4]
  assign _T_1527 = StickySelects_14_io_outs_4; // @[MemPrimitives.scala 126:35:@14129.4]
  assign _T_1528 = StickySelects_14_io_outs_5; // @[MemPrimitives.scala 126:35:@14130.4]
  assign _T_1530 = {_T_1523,io_rPort_2_backpressure,io_rPort_2_ofs_0}; // @[Cat.scala 30:58:@14132.4]
  assign _T_1532 = {_T_1524,io_rPort_4_backpressure,io_rPort_4_ofs_0}; // @[Cat.scala 30:58:@14134.4]
  assign _T_1534 = {_T_1525,io_rPort_6_backpressure,io_rPort_6_ofs_0}; // @[Cat.scala 30:58:@14136.4]
  assign _T_1536 = {_T_1526,io_rPort_7_backpressure,io_rPort_7_ofs_0}; // @[Cat.scala 30:58:@14138.4]
  assign _T_1538 = {_T_1527,io_rPort_8_backpressure,io_rPort_8_ofs_0}; // @[Cat.scala 30:58:@14140.4]
  assign _T_1540 = {_T_1528,io_rPort_10_backpressure,io_rPort_10_ofs_0}; // @[Cat.scala 30:58:@14142.4]
  assign _T_1541 = _T_1527 ? _T_1538 : _T_1540; // @[Mux.scala 31:69:@14143.4]
  assign _T_1542 = _T_1526 ? _T_1536 : _T_1541; // @[Mux.scala 31:69:@14144.4]
  assign _T_1543 = _T_1525 ? _T_1534 : _T_1542; // @[Mux.scala 31:69:@14145.4]
  assign _T_1544 = _T_1524 ? _T_1532 : _T_1543; // @[Mux.scala 31:69:@14146.4]
  assign _T_1545 = _T_1523 ? _T_1530 : _T_1544; // @[Mux.scala 31:69:@14147.4]
  assign _T_1553 = _T_1426 & _T_808; // @[MemPrimitives.scala 110:228:@14156.4]
  assign _T_1559 = _T_1432 & _T_814; // @[MemPrimitives.scala 110:228:@14160.4]
  assign _T_1565 = _T_1438 & _T_820; // @[MemPrimitives.scala 110:228:@14164.4]
  assign _T_1571 = _T_1444 & _T_826; // @[MemPrimitives.scala 110:228:@14168.4]
  assign _T_1577 = _T_1450 & _T_832; // @[MemPrimitives.scala 110:228:@14172.4]
  assign _T_1583 = _T_1456 & _T_838; // @[MemPrimitives.scala 110:228:@14176.4]
  assign _T_1585 = StickySelects_15_io_outs_0; // @[MemPrimitives.scala 126:35:@14187.4]
  assign _T_1586 = StickySelects_15_io_outs_1; // @[MemPrimitives.scala 126:35:@14188.4]
  assign _T_1587 = StickySelects_15_io_outs_2; // @[MemPrimitives.scala 126:35:@14189.4]
  assign _T_1588 = StickySelects_15_io_outs_3; // @[MemPrimitives.scala 126:35:@14190.4]
  assign _T_1589 = StickySelects_15_io_outs_4; // @[MemPrimitives.scala 126:35:@14191.4]
  assign _T_1590 = StickySelects_15_io_outs_5; // @[MemPrimitives.scala 126:35:@14192.4]
  assign _T_1592 = {_T_1585,io_rPort_0_backpressure,io_rPort_0_ofs_0}; // @[Cat.scala 30:58:@14194.4]
  assign _T_1594 = {_T_1586,io_rPort_1_backpressure,io_rPort_1_ofs_0}; // @[Cat.scala 30:58:@14196.4]
  assign _T_1596 = {_T_1587,io_rPort_3_backpressure,io_rPort_3_ofs_0}; // @[Cat.scala 30:58:@14198.4]
  assign _T_1598 = {_T_1588,io_rPort_5_backpressure,io_rPort_5_ofs_0}; // @[Cat.scala 30:58:@14200.4]
  assign _T_1600 = {_T_1589,io_rPort_9_backpressure,io_rPort_9_ofs_0}; // @[Cat.scala 30:58:@14202.4]
  assign _T_1602 = {_T_1590,io_rPort_11_backpressure,io_rPort_11_ofs_0}; // @[Cat.scala 30:58:@14204.4]
  assign _T_1603 = _T_1589 ? _T_1600 : _T_1602; // @[Mux.scala 31:69:@14205.4]
  assign _T_1604 = _T_1588 ? _T_1598 : _T_1603; // @[Mux.scala 31:69:@14206.4]
  assign _T_1605 = _T_1587 ? _T_1596 : _T_1604; // @[Mux.scala 31:69:@14207.4]
  assign _T_1606 = _T_1586 ? _T_1594 : _T_1605; // @[Mux.scala 31:69:@14208.4]
  assign _T_1607 = _T_1585 ? _T_1592 : _T_1606; // @[Mux.scala 31:69:@14209.4]
  assign _T_1671 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@14294.4 package.scala 96:25:@14295.4]
  assign _T_1675 = _T_1671 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14304.4]
  assign _T_1668 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@14286.4 package.scala 96:25:@14287.4]
  assign _T_1676 = _T_1668 ? Mem1D_11_io_output : _T_1675; // @[Mux.scala 31:69:@14305.4]
  assign _T_1665 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@14278.4 package.scala 96:25:@14279.4]
  assign _T_1677 = _T_1665 ? Mem1D_9_io_output : _T_1676; // @[Mux.scala 31:69:@14306.4]
  assign _T_1662 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@14270.4 package.scala 96:25:@14271.4]
  assign _T_1678 = _T_1662 ? Mem1D_7_io_output : _T_1677; // @[Mux.scala 31:69:@14307.4]
  assign _T_1659 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@14262.4 package.scala 96:25:@14263.4]
  assign _T_1679 = _T_1659 ? Mem1D_5_io_output : _T_1678; // @[Mux.scala 31:69:@14308.4]
  assign _T_1656 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@14254.4 package.scala 96:25:@14255.4]
  assign _T_1680 = _T_1656 ? Mem1D_3_io_output : _T_1679; // @[Mux.scala 31:69:@14309.4]
  assign _T_1653 = RetimeWrapper_io_out; // @[package.scala 96:25:@14246.4 package.scala 96:25:@14247.4]
  assign _T_1742 = RetimeWrapper_14_io_out; // @[package.scala 96:25:@14390.4 package.scala 96:25:@14391.4]
  assign _T_1746 = _T_1742 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14400.4]
  assign _T_1739 = RetimeWrapper_13_io_out; // @[package.scala 96:25:@14382.4 package.scala 96:25:@14383.4]
  assign _T_1747 = _T_1739 ? Mem1D_11_io_output : _T_1746; // @[Mux.scala 31:69:@14401.4]
  assign _T_1736 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@14374.4 package.scala 96:25:@14375.4]
  assign _T_1748 = _T_1736 ? Mem1D_9_io_output : _T_1747; // @[Mux.scala 31:69:@14402.4]
  assign _T_1733 = RetimeWrapper_11_io_out; // @[package.scala 96:25:@14366.4 package.scala 96:25:@14367.4]
  assign _T_1749 = _T_1733 ? Mem1D_7_io_output : _T_1748; // @[Mux.scala 31:69:@14403.4]
  assign _T_1730 = RetimeWrapper_10_io_out; // @[package.scala 96:25:@14358.4 package.scala 96:25:@14359.4]
  assign _T_1750 = _T_1730 ? Mem1D_5_io_output : _T_1749; // @[Mux.scala 31:69:@14404.4]
  assign _T_1727 = RetimeWrapper_9_io_out; // @[package.scala 96:25:@14350.4 package.scala 96:25:@14351.4]
  assign _T_1751 = _T_1727 ? Mem1D_3_io_output : _T_1750; // @[Mux.scala 31:69:@14405.4]
  assign _T_1724 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@14342.4 package.scala 96:25:@14343.4]
  assign _T_1813 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@14486.4 package.scala 96:25:@14487.4]
  assign _T_1817 = _T_1813 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14496.4]
  assign _T_1810 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@14478.4 package.scala 96:25:@14479.4]
  assign _T_1818 = _T_1810 ? Mem1D_10_io_output : _T_1817; // @[Mux.scala 31:69:@14497.4]
  assign _T_1807 = RetimeWrapper_20_io_out; // @[package.scala 96:25:@14470.4 package.scala 96:25:@14471.4]
  assign _T_1819 = _T_1807 ? Mem1D_8_io_output : _T_1818; // @[Mux.scala 31:69:@14498.4]
  assign _T_1804 = RetimeWrapper_19_io_out; // @[package.scala 96:25:@14462.4 package.scala 96:25:@14463.4]
  assign _T_1820 = _T_1804 ? Mem1D_6_io_output : _T_1819; // @[Mux.scala 31:69:@14499.4]
  assign _T_1801 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@14454.4 package.scala 96:25:@14455.4]
  assign _T_1821 = _T_1801 ? Mem1D_4_io_output : _T_1820; // @[Mux.scala 31:69:@14500.4]
  assign _T_1798 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@14446.4 package.scala 96:25:@14447.4]
  assign _T_1822 = _T_1798 ? Mem1D_2_io_output : _T_1821; // @[Mux.scala 31:69:@14501.4]
  assign _T_1795 = RetimeWrapper_16_io_out; // @[package.scala 96:25:@14438.4 package.scala 96:25:@14439.4]
  assign _T_1884 = RetimeWrapper_30_io_out; // @[package.scala 96:25:@14582.4 package.scala 96:25:@14583.4]
  assign _T_1888 = _T_1884 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14592.4]
  assign _T_1881 = RetimeWrapper_29_io_out; // @[package.scala 96:25:@14574.4 package.scala 96:25:@14575.4]
  assign _T_1889 = _T_1881 ? Mem1D_11_io_output : _T_1888; // @[Mux.scala 31:69:@14593.4]
  assign _T_1878 = RetimeWrapper_28_io_out; // @[package.scala 96:25:@14566.4 package.scala 96:25:@14567.4]
  assign _T_1890 = _T_1878 ? Mem1D_9_io_output : _T_1889; // @[Mux.scala 31:69:@14594.4]
  assign _T_1875 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@14558.4 package.scala 96:25:@14559.4]
  assign _T_1891 = _T_1875 ? Mem1D_7_io_output : _T_1890; // @[Mux.scala 31:69:@14595.4]
  assign _T_1872 = RetimeWrapper_26_io_out; // @[package.scala 96:25:@14550.4 package.scala 96:25:@14551.4]
  assign _T_1892 = _T_1872 ? Mem1D_5_io_output : _T_1891; // @[Mux.scala 31:69:@14596.4]
  assign _T_1869 = RetimeWrapper_25_io_out; // @[package.scala 96:25:@14542.4 package.scala 96:25:@14543.4]
  assign _T_1893 = _T_1869 ? Mem1D_3_io_output : _T_1892; // @[Mux.scala 31:69:@14597.4]
  assign _T_1866 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@14534.4 package.scala 96:25:@14535.4]
  assign _T_1955 = RetimeWrapper_38_io_out; // @[package.scala 96:25:@14678.4 package.scala 96:25:@14679.4]
  assign _T_1959 = _T_1955 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14688.4]
  assign _T_1952 = RetimeWrapper_37_io_out; // @[package.scala 96:25:@14670.4 package.scala 96:25:@14671.4]
  assign _T_1960 = _T_1952 ? Mem1D_10_io_output : _T_1959; // @[Mux.scala 31:69:@14689.4]
  assign _T_1949 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@14662.4 package.scala 96:25:@14663.4]
  assign _T_1961 = _T_1949 ? Mem1D_8_io_output : _T_1960; // @[Mux.scala 31:69:@14690.4]
  assign _T_1946 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@14654.4 package.scala 96:25:@14655.4]
  assign _T_1962 = _T_1946 ? Mem1D_6_io_output : _T_1961; // @[Mux.scala 31:69:@14691.4]
  assign _T_1943 = RetimeWrapper_34_io_out; // @[package.scala 96:25:@14646.4 package.scala 96:25:@14647.4]
  assign _T_1963 = _T_1943 ? Mem1D_4_io_output : _T_1962; // @[Mux.scala 31:69:@14692.4]
  assign _T_1940 = RetimeWrapper_33_io_out; // @[package.scala 96:25:@14638.4 package.scala 96:25:@14639.4]
  assign _T_1964 = _T_1940 ? Mem1D_2_io_output : _T_1963; // @[Mux.scala 31:69:@14693.4]
  assign _T_1937 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@14630.4 package.scala 96:25:@14631.4]
  assign _T_2026 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@14774.4 package.scala 96:25:@14775.4]
  assign _T_2030 = _T_2026 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@14784.4]
  assign _T_2023 = RetimeWrapper_45_io_out; // @[package.scala 96:25:@14766.4 package.scala 96:25:@14767.4]
  assign _T_2031 = _T_2023 ? Mem1D_11_io_output : _T_2030; // @[Mux.scala 31:69:@14785.4]
  assign _T_2020 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@14758.4 package.scala 96:25:@14759.4]
  assign _T_2032 = _T_2020 ? Mem1D_9_io_output : _T_2031; // @[Mux.scala 31:69:@14786.4]
  assign _T_2017 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@14750.4 package.scala 96:25:@14751.4]
  assign _T_2033 = _T_2017 ? Mem1D_7_io_output : _T_2032; // @[Mux.scala 31:69:@14787.4]
  assign _T_2014 = RetimeWrapper_42_io_out; // @[package.scala 96:25:@14742.4 package.scala 96:25:@14743.4]
  assign _T_2034 = _T_2014 ? Mem1D_5_io_output : _T_2033; // @[Mux.scala 31:69:@14788.4]
  assign _T_2011 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@14734.4 package.scala 96:25:@14735.4]
  assign _T_2035 = _T_2011 ? Mem1D_3_io_output : _T_2034; // @[Mux.scala 31:69:@14789.4]
  assign _T_2008 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@14726.4 package.scala 96:25:@14727.4]
  assign _T_2097 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@14870.4 package.scala 96:25:@14871.4]
  assign _T_2101 = _T_2097 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14880.4]
  assign _T_2094 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@14862.4 package.scala 96:25:@14863.4]
  assign _T_2102 = _T_2094 ? Mem1D_10_io_output : _T_2101; // @[Mux.scala 31:69:@14881.4]
  assign _T_2091 = RetimeWrapper_52_io_out; // @[package.scala 96:25:@14854.4 package.scala 96:25:@14855.4]
  assign _T_2103 = _T_2091 ? Mem1D_8_io_output : _T_2102; // @[Mux.scala 31:69:@14882.4]
  assign _T_2088 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@14846.4 package.scala 96:25:@14847.4]
  assign _T_2104 = _T_2088 ? Mem1D_6_io_output : _T_2103; // @[Mux.scala 31:69:@14883.4]
  assign _T_2085 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@14838.4 package.scala 96:25:@14839.4]
  assign _T_2105 = _T_2085 ? Mem1D_4_io_output : _T_2104; // @[Mux.scala 31:69:@14884.4]
  assign _T_2082 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@14830.4 package.scala 96:25:@14831.4]
  assign _T_2106 = _T_2082 ? Mem1D_2_io_output : _T_2105; // @[Mux.scala 31:69:@14885.4]
  assign _T_2079 = RetimeWrapper_48_io_out; // @[package.scala 96:25:@14822.4 package.scala 96:25:@14823.4]
  assign _T_2168 = RetimeWrapper_62_io_out; // @[package.scala 96:25:@14966.4 package.scala 96:25:@14967.4]
  assign _T_2172 = _T_2168 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@14976.4]
  assign _T_2165 = RetimeWrapper_61_io_out; // @[package.scala 96:25:@14958.4 package.scala 96:25:@14959.4]
  assign _T_2173 = _T_2165 ? Mem1D_10_io_output : _T_2172; // @[Mux.scala 31:69:@14977.4]
  assign _T_2162 = RetimeWrapper_60_io_out; // @[package.scala 96:25:@14950.4 package.scala 96:25:@14951.4]
  assign _T_2174 = _T_2162 ? Mem1D_8_io_output : _T_2173; // @[Mux.scala 31:69:@14978.4]
  assign _T_2159 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@14942.4 package.scala 96:25:@14943.4]
  assign _T_2175 = _T_2159 ? Mem1D_6_io_output : _T_2174; // @[Mux.scala 31:69:@14979.4]
  assign _T_2156 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@14934.4 package.scala 96:25:@14935.4]
  assign _T_2176 = _T_2156 ? Mem1D_4_io_output : _T_2175; // @[Mux.scala 31:69:@14980.4]
  assign _T_2153 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@14926.4 package.scala 96:25:@14927.4]
  assign _T_2177 = _T_2153 ? Mem1D_2_io_output : _T_2176; // @[Mux.scala 31:69:@14981.4]
  assign _T_2150 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@14918.4 package.scala 96:25:@14919.4]
  assign _T_2239 = RetimeWrapper_70_io_out; // @[package.scala 96:25:@15062.4 package.scala 96:25:@15063.4]
  assign _T_2243 = _T_2239 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@15072.4]
  assign _T_2236 = RetimeWrapper_69_io_out; // @[package.scala 96:25:@15054.4 package.scala 96:25:@15055.4]
  assign _T_2244 = _T_2236 ? Mem1D_10_io_output : _T_2243; // @[Mux.scala 31:69:@15073.4]
  assign _T_2233 = RetimeWrapper_68_io_out; // @[package.scala 96:25:@15046.4 package.scala 96:25:@15047.4]
  assign _T_2245 = _T_2233 ? Mem1D_8_io_output : _T_2244; // @[Mux.scala 31:69:@15074.4]
  assign _T_2230 = RetimeWrapper_67_io_out; // @[package.scala 96:25:@15038.4 package.scala 96:25:@15039.4]
  assign _T_2246 = _T_2230 ? Mem1D_6_io_output : _T_2245; // @[Mux.scala 31:69:@15075.4]
  assign _T_2227 = RetimeWrapper_66_io_out; // @[package.scala 96:25:@15030.4 package.scala 96:25:@15031.4]
  assign _T_2247 = _T_2227 ? Mem1D_4_io_output : _T_2246; // @[Mux.scala 31:69:@15076.4]
  assign _T_2224 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@15022.4 package.scala 96:25:@15023.4]
  assign _T_2248 = _T_2224 ? Mem1D_2_io_output : _T_2247; // @[Mux.scala 31:69:@15077.4]
  assign _T_2221 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@15014.4 package.scala 96:25:@15015.4]
  assign _T_2310 = RetimeWrapper_78_io_out; // @[package.scala 96:25:@15158.4 package.scala 96:25:@15159.4]
  assign _T_2314 = _T_2310 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15168.4]
  assign _T_2307 = RetimeWrapper_77_io_out; // @[package.scala 96:25:@15150.4 package.scala 96:25:@15151.4]
  assign _T_2315 = _T_2307 ? Mem1D_11_io_output : _T_2314; // @[Mux.scala 31:69:@15169.4]
  assign _T_2304 = RetimeWrapper_76_io_out; // @[package.scala 96:25:@15142.4 package.scala 96:25:@15143.4]
  assign _T_2316 = _T_2304 ? Mem1D_9_io_output : _T_2315; // @[Mux.scala 31:69:@15170.4]
  assign _T_2301 = RetimeWrapper_75_io_out; // @[package.scala 96:25:@15134.4 package.scala 96:25:@15135.4]
  assign _T_2317 = _T_2301 ? Mem1D_7_io_output : _T_2316; // @[Mux.scala 31:69:@15171.4]
  assign _T_2298 = RetimeWrapper_74_io_out; // @[package.scala 96:25:@15126.4 package.scala 96:25:@15127.4]
  assign _T_2318 = _T_2298 ? Mem1D_5_io_output : _T_2317; // @[Mux.scala 31:69:@15172.4]
  assign _T_2295 = RetimeWrapper_73_io_out; // @[package.scala 96:25:@15118.4 package.scala 96:25:@15119.4]
  assign _T_2319 = _T_2295 ? Mem1D_3_io_output : _T_2318; // @[Mux.scala 31:69:@15173.4]
  assign _T_2292 = RetimeWrapper_72_io_out; // @[package.scala 96:25:@15110.4 package.scala 96:25:@15111.4]
  assign _T_2381 = RetimeWrapper_86_io_out; // @[package.scala 96:25:@15254.4 package.scala 96:25:@15255.4]
  assign _T_2385 = _T_2381 ? Mem1D_12_io_output : Mem1D_14_io_output; // @[Mux.scala 31:69:@15264.4]
  assign _T_2378 = RetimeWrapper_85_io_out; // @[package.scala 96:25:@15246.4 package.scala 96:25:@15247.4]
  assign _T_2386 = _T_2378 ? Mem1D_10_io_output : _T_2385; // @[Mux.scala 31:69:@15265.4]
  assign _T_2375 = RetimeWrapper_84_io_out; // @[package.scala 96:25:@15238.4 package.scala 96:25:@15239.4]
  assign _T_2387 = _T_2375 ? Mem1D_8_io_output : _T_2386; // @[Mux.scala 31:69:@15266.4]
  assign _T_2372 = RetimeWrapper_83_io_out; // @[package.scala 96:25:@15230.4 package.scala 96:25:@15231.4]
  assign _T_2388 = _T_2372 ? Mem1D_6_io_output : _T_2387; // @[Mux.scala 31:69:@15267.4]
  assign _T_2369 = RetimeWrapper_82_io_out; // @[package.scala 96:25:@15222.4 package.scala 96:25:@15223.4]
  assign _T_2389 = _T_2369 ? Mem1D_4_io_output : _T_2388; // @[Mux.scala 31:69:@15268.4]
  assign _T_2366 = RetimeWrapper_81_io_out; // @[package.scala 96:25:@15214.4 package.scala 96:25:@15215.4]
  assign _T_2390 = _T_2366 ? Mem1D_2_io_output : _T_2389; // @[Mux.scala 31:69:@15269.4]
  assign _T_2363 = RetimeWrapper_80_io_out; // @[package.scala 96:25:@15206.4 package.scala 96:25:@15207.4]
  assign _T_2452 = RetimeWrapper_94_io_out; // @[package.scala 96:25:@15350.4 package.scala 96:25:@15351.4]
  assign _T_2456 = _T_2452 ? Mem1D_13_io_output : Mem1D_15_io_output; // @[Mux.scala 31:69:@15360.4]
  assign _T_2449 = RetimeWrapper_93_io_out; // @[package.scala 96:25:@15342.4 package.scala 96:25:@15343.4]
  assign _T_2457 = _T_2449 ? Mem1D_11_io_output : _T_2456; // @[Mux.scala 31:69:@15361.4]
  assign _T_2446 = RetimeWrapper_92_io_out; // @[package.scala 96:25:@15334.4 package.scala 96:25:@15335.4]
  assign _T_2458 = _T_2446 ? Mem1D_9_io_output : _T_2457; // @[Mux.scala 31:69:@15362.4]
  assign _T_2443 = RetimeWrapper_91_io_out; // @[package.scala 96:25:@15326.4 package.scala 96:25:@15327.4]
  assign _T_2459 = _T_2443 ? Mem1D_7_io_output : _T_2458; // @[Mux.scala 31:69:@15363.4]
  assign _T_2440 = RetimeWrapper_90_io_out; // @[package.scala 96:25:@15318.4 package.scala 96:25:@15319.4]
  assign _T_2460 = _T_2440 ? Mem1D_5_io_output : _T_2459; // @[Mux.scala 31:69:@15364.4]
  assign _T_2437 = RetimeWrapper_89_io_out; // @[package.scala 96:25:@15310.4 package.scala 96:25:@15311.4]
  assign _T_2461 = _T_2437 ? Mem1D_3_io_output : _T_2460; // @[Mux.scala 31:69:@15365.4]
  assign _T_2434 = RetimeWrapper_88_io_out; // @[package.scala 96:25:@15302.4 package.scala 96:25:@15303.4]
  assign io_rPort_11_output_0 = _T_2434 ? Mem1D_1_io_output : _T_2461; // @[MemPrimitives.scala 152:13:@15367.4]
  assign io_rPort_10_output_0 = _T_2363 ? Mem1D_io_output : _T_2390; // @[MemPrimitives.scala 152:13:@15271.4]
  assign io_rPort_9_output_0 = _T_2292 ? Mem1D_1_io_output : _T_2319; // @[MemPrimitives.scala 152:13:@15175.4]
  assign io_rPort_8_output_0 = _T_2221 ? Mem1D_io_output : _T_2248; // @[MemPrimitives.scala 152:13:@15079.4]
  assign io_rPort_7_output_0 = _T_2150 ? Mem1D_io_output : _T_2177; // @[MemPrimitives.scala 152:13:@14983.4]
  assign io_rPort_6_output_0 = _T_2079 ? Mem1D_io_output : _T_2106; // @[MemPrimitives.scala 152:13:@14887.4]
  assign io_rPort_5_output_0 = _T_2008 ? Mem1D_1_io_output : _T_2035; // @[MemPrimitives.scala 152:13:@14791.4]
  assign io_rPort_4_output_0 = _T_1937 ? Mem1D_io_output : _T_1964; // @[MemPrimitives.scala 152:13:@14695.4]
  assign io_rPort_3_output_0 = _T_1866 ? Mem1D_1_io_output : _T_1893; // @[MemPrimitives.scala 152:13:@14599.4]
  assign io_rPort_2_output_0 = _T_1795 ? Mem1D_io_output : _T_1822; // @[MemPrimitives.scala 152:13:@14503.4]
  assign io_rPort_1_output_0 = _T_1724 ? Mem1D_1_io_output : _T_1751; // @[MemPrimitives.scala 152:13:@14407.4]
  assign io_rPort_0_output_0 = _T_1653 ? Mem1D_1_io_output : _T_1680; // @[MemPrimitives.scala 152:13:@14311.4]
  assign Mem1D_clock = clock; // @[:@12777.4]
  assign Mem1D_reset = reset; // @[:@12778.4]
  assign Mem1D_io_r_ofs_0 = _T_677[8:0]; // @[MemPrimitives.scala 131:28:@13283.4]
  assign Mem1D_io_r_backpressure = _T_677[9]; // @[MemPrimitives.scala 132:32:@13284.4]
  assign Mem1D_io_w_ofs_0 = _T_450[8:0]; // @[MemPrimitives.scala 94:28:@13041.4]
  assign Mem1D_io_w_data_0 = _T_450[40:9]; // @[MemPrimitives.scala 95:29:@13042.4]
  assign Mem1D_io_w_en_0 = _T_450[41]; // @[MemPrimitives.scala 96:27:@13043.4]
  assign Mem1D_1_clock = clock; // @[:@12793.4]
  assign Mem1D_1_reset = reset; // @[:@12794.4]
  assign Mem1D_1_io_r_ofs_0 = _T_739[8:0]; // @[MemPrimitives.scala 131:28:@13345.4]
  assign Mem1D_1_io_r_backpressure = _T_739[9]; // @[MemPrimitives.scala 132:32:@13346.4]
  assign Mem1D_1_io_w_ofs_0 = _T_461[8:0]; // @[MemPrimitives.scala 94:28:@13053.4]
  assign Mem1D_1_io_w_data_0 = _T_461[40:9]; // @[MemPrimitives.scala 95:29:@13054.4]
  assign Mem1D_1_io_w_en_0 = _T_461[41]; // @[MemPrimitives.scala 96:27:@13055.4]
  assign Mem1D_2_clock = clock; // @[:@12809.4]
  assign Mem1D_2_reset = reset; // @[:@12810.4]
  assign Mem1D_2_io_r_ofs_0 = _T_801[8:0]; // @[MemPrimitives.scala 131:28:@13407.4]
  assign Mem1D_2_io_r_backpressure = _T_801[9]; // @[MemPrimitives.scala 132:32:@13408.4]
  assign Mem1D_2_io_w_ofs_0 = _T_472[8:0]; // @[MemPrimitives.scala 94:28:@13065.4]
  assign Mem1D_2_io_w_data_0 = _T_472[40:9]; // @[MemPrimitives.scala 95:29:@13066.4]
  assign Mem1D_2_io_w_en_0 = _T_472[41]; // @[MemPrimitives.scala 96:27:@13067.4]
  assign Mem1D_3_clock = clock; // @[:@12825.4]
  assign Mem1D_3_reset = reset; // @[:@12826.4]
  assign Mem1D_3_io_r_ofs_0 = _T_863[8:0]; // @[MemPrimitives.scala 131:28:@13469.4]
  assign Mem1D_3_io_r_backpressure = _T_863[9]; // @[MemPrimitives.scala 132:32:@13470.4]
  assign Mem1D_3_io_w_ofs_0 = _T_483[8:0]; // @[MemPrimitives.scala 94:28:@13077.4]
  assign Mem1D_3_io_w_data_0 = _T_483[40:9]; // @[MemPrimitives.scala 95:29:@13078.4]
  assign Mem1D_3_io_w_en_0 = _T_483[41]; // @[MemPrimitives.scala 96:27:@13079.4]
  assign Mem1D_4_clock = clock; // @[:@12841.4]
  assign Mem1D_4_reset = reset; // @[:@12842.4]
  assign Mem1D_4_io_r_ofs_0 = _T_925[8:0]; // @[MemPrimitives.scala 131:28:@13531.4]
  assign Mem1D_4_io_r_backpressure = _T_925[9]; // @[MemPrimitives.scala 132:32:@13532.4]
  assign Mem1D_4_io_w_ofs_0 = _T_494[8:0]; // @[MemPrimitives.scala 94:28:@13089.4]
  assign Mem1D_4_io_w_data_0 = _T_494[40:9]; // @[MemPrimitives.scala 95:29:@13090.4]
  assign Mem1D_4_io_w_en_0 = _T_494[41]; // @[MemPrimitives.scala 96:27:@13091.4]
  assign Mem1D_5_clock = clock; // @[:@12857.4]
  assign Mem1D_5_reset = reset; // @[:@12858.4]
  assign Mem1D_5_io_r_ofs_0 = _T_987[8:0]; // @[MemPrimitives.scala 131:28:@13593.4]
  assign Mem1D_5_io_r_backpressure = _T_987[9]; // @[MemPrimitives.scala 132:32:@13594.4]
  assign Mem1D_5_io_w_ofs_0 = _T_505[8:0]; // @[MemPrimitives.scala 94:28:@13101.4]
  assign Mem1D_5_io_w_data_0 = _T_505[40:9]; // @[MemPrimitives.scala 95:29:@13102.4]
  assign Mem1D_5_io_w_en_0 = _T_505[41]; // @[MemPrimitives.scala 96:27:@13103.4]
  assign Mem1D_6_clock = clock; // @[:@12873.4]
  assign Mem1D_6_reset = reset; // @[:@12874.4]
  assign Mem1D_6_io_r_ofs_0 = _T_1049[8:0]; // @[MemPrimitives.scala 131:28:@13655.4]
  assign Mem1D_6_io_r_backpressure = _T_1049[9]; // @[MemPrimitives.scala 132:32:@13656.4]
  assign Mem1D_6_io_w_ofs_0 = _T_516[8:0]; // @[MemPrimitives.scala 94:28:@13113.4]
  assign Mem1D_6_io_w_data_0 = _T_516[40:9]; // @[MemPrimitives.scala 95:29:@13114.4]
  assign Mem1D_6_io_w_en_0 = _T_516[41]; // @[MemPrimitives.scala 96:27:@13115.4]
  assign Mem1D_7_clock = clock; // @[:@12889.4]
  assign Mem1D_7_reset = reset; // @[:@12890.4]
  assign Mem1D_7_io_r_ofs_0 = _T_1111[8:0]; // @[MemPrimitives.scala 131:28:@13717.4]
  assign Mem1D_7_io_r_backpressure = _T_1111[9]; // @[MemPrimitives.scala 132:32:@13718.4]
  assign Mem1D_7_io_w_ofs_0 = _T_527[8:0]; // @[MemPrimitives.scala 94:28:@13125.4]
  assign Mem1D_7_io_w_data_0 = _T_527[40:9]; // @[MemPrimitives.scala 95:29:@13126.4]
  assign Mem1D_7_io_w_en_0 = _T_527[41]; // @[MemPrimitives.scala 96:27:@13127.4]
  assign Mem1D_8_clock = clock; // @[:@12905.4]
  assign Mem1D_8_reset = reset; // @[:@12906.4]
  assign Mem1D_8_io_r_ofs_0 = _T_1173[8:0]; // @[MemPrimitives.scala 131:28:@13779.4]
  assign Mem1D_8_io_r_backpressure = _T_1173[9]; // @[MemPrimitives.scala 132:32:@13780.4]
  assign Mem1D_8_io_w_ofs_0 = _T_538[8:0]; // @[MemPrimitives.scala 94:28:@13137.4]
  assign Mem1D_8_io_w_data_0 = _T_538[40:9]; // @[MemPrimitives.scala 95:29:@13138.4]
  assign Mem1D_8_io_w_en_0 = _T_538[41]; // @[MemPrimitives.scala 96:27:@13139.4]
  assign Mem1D_9_clock = clock; // @[:@12921.4]
  assign Mem1D_9_reset = reset; // @[:@12922.4]
  assign Mem1D_9_io_r_ofs_0 = _T_1235[8:0]; // @[MemPrimitives.scala 131:28:@13841.4]
  assign Mem1D_9_io_r_backpressure = _T_1235[9]; // @[MemPrimitives.scala 132:32:@13842.4]
  assign Mem1D_9_io_w_ofs_0 = _T_549[8:0]; // @[MemPrimitives.scala 94:28:@13149.4]
  assign Mem1D_9_io_w_data_0 = _T_549[40:9]; // @[MemPrimitives.scala 95:29:@13150.4]
  assign Mem1D_9_io_w_en_0 = _T_549[41]; // @[MemPrimitives.scala 96:27:@13151.4]
  assign Mem1D_10_clock = clock; // @[:@12937.4]
  assign Mem1D_10_reset = reset; // @[:@12938.4]
  assign Mem1D_10_io_r_ofs_0 = _T_1297[8:0]; // @[MemPrimitives.scala 131:28:@13903.4]
  assign Mem1D_10_io_r_backpressure = _T_1297[9]; // @[MemPrimitives.scala 132:32:@13904.4]
  assign Mem1D_10_io_w_ofs_0 = _T_560[8:0]; // @[MemPrimitives.scala 94:28:@13161.4]
  assign Mem1D_10_io_w_data_0 = _T_560[40:9]; // @[MemPrimitives.scala 95:29:@13162.4]
  assign Mem1D_10_io_w_en_0 = _T_560[41]; // @[MemPrimitives.scala 96:27:@13163.4]
  assign Mem1D_11_clock = clock; // @[:@12953.4]
  assign Mem1D_11_reset = reset; // @[:@12954.4]
  assign Mem1D_11_io_r_ofs_0 = _T_1359[8:0]; // @[MemPrimitives.scala 131:28:@13965.4]
  assign Mem1D_11_io_r_backpressure = _T_1359[9]; // @[MemPrimitives.scala 132:32:@13966.4]
  assign Mem1D_11_io_w_ofs_0 = _T_571[8:0]; // @[MemPrimitives.scala 94:28:@13173.4]
  assign Mem1D_11_io_w_data_0 = _T_571[40:9]; // @[MemPrimitives.scala 95:29:@13174.4]
  assign Mem1D_11_io_w_en_0 = _T_571[41]; // @[MemPrimitives.scala 96:27:@13175.4]
  assign Mem1D_12_clock = clock; // @[:@12969.4]
  assign Mem1D_12_reset = reset; // @[:@12970.4]
  assign Mem1D_12_io_r_ofs_0 = _T_1421[8:0]; // @[MemPrimitives.scala 131:28:@14027.4]
  assign Mem1D_12_io_r_backpressure = _T_1421[9]; // @[MemPrimitives.scala 132:32:@14028.4]
  assign Mem1D_12_io_w_ofs_0 = _T_582[8:0]; // @[MemPrimitives.scala 94:28:@13185.4]
  assign Mem1D_12_io_w_data_0 = _T_582[40:9]; // @[MemPrimitives.scala 95:29:@13186.4]
  assign Mem1D_12_io_w_en_0 = _T_582[41]; // @[MemPrimitives.scala 96:27:@13187.4]
  assign Mem1D_13_clock = clock; // @[:@12985.4]
  assign Mem1D_13_reset = reset; // @[:@12986.4]
  assign Mem1D_13_io_r_ofs_0 = _T_1483[8:0]; // @[MemPrimitives.scala 131:28:@14089.4]
  assign Mem1D_13_io_r_backpressure = _T_1483[9]; // @[MemPrimitives.scala 132:32:@14090.4]
  assign Mem1D_13_io_w_ofs_0 = _T_593[8:0]; // @[MemPrimitives.scala 94:28:@13197.4]
  assign Mem1D_13_io_w_data_0 = _T_593[40:9]; // @[MemPrimitives.scala 95:29:@13198.4]
  assign Mem1D_13_io_w_en_0 = _T_593[41]; // @[MemPrimitives.scala 96:27:@13199.4]
  assign Mem1D_14_clock = clock; // @[:@13001.4]
  assign Mem1D_14_reset = reset; // @[:@13002.4]
  assign Mem1D_14_io_r_ofs_0 = _T_1545[8:0]; // @[MemPrimitives.scala 131:28:@14151.4]
  assign Mem1D_14_io_r_backpressure = _T_1545[9]; // @[MemPrimitives.scala 132:32:@14152.4]
  assign Mem1D_14_io_w_ofs_0 = _T_604[8:0]; // @[MemPrimitives.scala 94:28:@13209.4]
  assign Mem1D_14_io_w_data_0 = _T_604[40:9]; // @[MemPrimitives.scala 95:29:@13210.4]
  assign Mem1D_14_io_w_en_0 = _T_604[41]; // @[MemPrimitives.scala 96:27:@13211.4]
  assign Mem1D_15_clock = clock; // @[:@13017.4]
  assign Mem1D_15_reset = reset; // @[:@13018.4]
  assign Mem1D_15_io_r_ofs_0 = _T_1607[8:0]; // @[MemPrimitives.scala 131:28:@14213.4]
  assign Mem1D_15_io_r_backpressure = _T_1607[9]; // @[MemPrimitives.scala 132:32:@14214.4]
  assign Mem1D_15_io_w_ofs_0 = _T_615[8:0]; // @[MemPrimitives.scala 94:28:@13221.4]
  assign Mem1D_15_io_w_data_0 = _T_615[40:9]; // @[MemPrimitives.scala 95:29:@13222.4]
  assign Mem1D_15_io_w_en_0 = _T_615[41]; // @[MemPrimitives.scala 96:27:@13223.4]
  assign StickySelects_clock = clock; // @[:@13249.4]
  assign StickySelects_reset = reset; // @[:@13250.4]
  assign StickySelects_io_ins_0 = io_rPort_2_en_0 & _T_623; // @[MemPrimitives.scala 125:64:@13251.4]
  assign StickySelects_io_ins_1 = io_rPort_4_en_0 & _T_629; // @[MemPrimitives.scala 125:64:@13252.4]
  assign StickySelects_io_ins_2 = io_rPort_6_en_0 & _T_635; // @[MemPrimitives.scala 125:64:@13253.4]
  assign StickySelects_io_ins_3 = io_rPort_7_en_0 & _T_641; // @[MemPrimitives.scala 125:64:@13254.4]
  assign StickySelects_io_ins_4 = io_rPort_8_en_0 & _T_647; // @[MemPrimitives.scala 125:64:@13255.4]
  assign StickySelects_io_ins_5 = io_rPort_10_en_0 & _T_653; // @[MemPrimitives.scala 125:64:@13256.4]
  assign StickySelects_1_clock = clock; // @[:@13311.4]
  assign StickySelects_1_reset = reset; // @[:@13312.4]
  assign StickySelects_1_io_ins_0 = io_rPort_0_en_0 & _T_685; // @[MemPrimitives.scala 125:64:@13313.4]
  assign StickySelects_1_io_ins_1 = io_rPort_1_en_0 & _T_691; // @[MemPrimitives.scala 125:64:@13314.4]
  assign StickySelects_1_io_ins_2 = io_rPort_3_en_0 & _T_697; // @[MemPrimitives.scala 125:64:@13315.4]
  assign StickySelects_1_io_ins_3 = io_rPort_5_en_0 & _T_703; // @[MemPrimitives.scala 125:64:@13316.4]
  assign StickySelects_1_io_ins_4 = io_rPort_9_en_0 & _T_709; // @[MemPrimitives.scala 125:64:@13317.4]
  assign StickySelects_1_io_ins_5 = io_rPort_11_en_0 & _T_715; // @[MemPrimitives.scala 125:64:@13318.4]
  assign StickySelects_2_clock = clock; // @[:@13373.4]
  assign StickySelects_2_reset = reset; // @[:@13374.4]
  assign StickySelects_2_io_ins_0 = io_rPort_2_en_0 & _T_747; // @[MemPrimitives.scala 125:64:@13375.4]
  assign StickySelects_2_io_ins_1 = io_rPort_4_en_0 & _T_753; // @[MemPrimitives.scala 125:64:@13376.4]
  assign StickySelects_2_io_ins_2 = io_rPort_6_en_0 & _T_759; // @[MemPrimitives.scala 125:64:@13377.4]
  assign StickySelects_2_io_ins_3 = io_rPort_7_en_0 & _T_765; // @[MemPrimitives.scala 125:64:@13378.4]
  assign StickySelects_2_io_ins_4 = io_rPort_8_en_0 & _T_771; // @[MemPrimitives.scala 125:64:@13379.4]
  assign StickySelects_2_io_ins_5 = io_rPort_10_en_0 & _T_777; // @[MemPrimitives.scala 125:64:@13380.4]
  assign StickySelects_3_clock = clock; // @[:@13435.4]
  assign StickySelects_3_reset = reset; // @[:@13436.4]
  assign StickySelects_3_io_ins_0 = io_rPort_0_en_0 & _T_809; // @[MemPrimitives.scala 125:64:@13437.4]
  assign StickySelects_3_io_ins_1 = io_rPort_1_en_0 & _T_815; // @[MemPrimitives.scala 125:64:@13438.4]
  assign StickySelects_3_io_ins_2 = io_rPort_3_en_0 & _T_821; // @[MemPrimitives.scala 125:64:@13439.4]
  assign StickySelects_3_io_ins_3 = io_rPort_5_en_0 & _T_827; // @[MemPrimitives.scala 125:64:@13440.4]
  assign StickySelects_3_io_ins_4 = io_rPort_9_en_0 & _T_833; // @[MemPrimitives.scala 125:64:@13441.4]
  assign StickySelects_3_io_ins_5 = io_rPort_11_en_0 & _T_839; // @[MemPrimitives.scala 125:64:@13442.4]
  assign StickySelects_4_clock = clock; // @[:@13497.4]
  assign StickySelects_4_reset = reset; // @[:@13498.4]
  assign StickySelects_4_io_ins_0 = io_rPort_2_en_0 & _T_871; // @[MemPrimitives.scala 125:64:@13499.4]
  assign StickySelects_4_io_ins_1 = io_rPort_4_en_0 & _T_877; // @[MemPrimitives.scala 125:64:@13500.4]
  assign StickySelects_4_io_ins_2 = io_rPort_6_en_0 & _T_883; // @[MemPrimitives.scala 125:64:@13501.4]
  assign StickySelects_4_io_ins_3 = io_rPort_7_en_0 & _T_889; // @[MemPrimitives.scala 125:64:@13502.4]
  assign StickySelects_4_io_ins_4 = io_rPort_8_en_0 & _T_895; // @[MemPrimitives.scala 125:64:@13503.4]
  assign StickySelects_4_io_ins_5 = io_rPort_10_en_0 & _T_901; // @[MemPrimitives.scala 125:64:@13504.4]
  assign StickySelects_5_clock = clock; // @[:@13559.4]
  assign StickySelects_5_reset = reset; // @[:@13560.4]
  assign StickySelects_5_io_ins_0 = io_rPort_0_en_0 & _T_933; // @[MemPrimitives.scala 125:64:@13561.4]
  assign StickySelects_5_io_ins_1 = io_rPort_1_en_0 & _T_939; // @[MemPrimitives.scala 125:64:@13562.4]
  assign StickySelects_5_io_ins_2 = io_rPort_3_en_0 & _T_945; // @[MemPrimitives.scala 125:64:@13563.4]
  assign StickySelects_5_io_ins_3 = io_rPort_5_en_0 & _T_951; // @[MemPrimitives.scala 125:64:@13564.4]
  assign StickySelects_5_io_ins_4 = io_rPort_9_en_0 & _T_957; // @[MemPrimitives.scala 125:64:@13565.4]
  assign StickySelects_5_io_ins_5 = io_rPort_11_en_0 & _T_963; // @[MemPrimitives.scala 125:64:@13566.4]
  assign StickySelects_6_clock = clock; // @[:@13621.4]
  assign StickySelects_6_reset = reset; // @[:@13622.4]
  assign StickySelects_6_io_ins_0 = io_rPort_2_en_0 & _T_995; // @[MemPrimitives.scala 125:64:@13623.4]
  assign StickySelects_6_io_ins_1 = io_rPort_4_en_0 & _T_1001; // @[MemPrimitives.scala 125:64:@13624.4]
  assign StickySelects_6_io_ins_2 = io_rPort_6_en_0 & _T_1007; // @[MemPrimitives.scala 125:64:@13625.4]
  assign StickySelects_6_io_ins_3 = io_rPort_7_en_0 & _T_1013; // @[MemPrimitives.scala 125:64:@13626.4]
  assign StickySelects_6_io_ins_4 = io_rPort_8_en_0 & _T_1019; // @[MemPrimitives.scala 125:64:@13627.4]
  assign StickySelects_6_io_ins_5 = io_rPort_10_en_0 & _T_1025; // @[MemPrimitives.scala 125:64:@13628.4]
  assign StickySelects_7_clock = clock; // @[:@13683.4]
  assign StickySelects_7_reset = reset; // @[:@13684.4]
  assign StickySelects_7_io_ins_0 = io_rPort_0_en_0 & _T_1057; // @[MemPrimitives.scala 125:64:@13685.4]
  assign StickySelects_7_io_ins_1 = io_rPort_1_en_0 & _T_1063; // @[MemPrimitives.scala 125:64:@13686.4]
  assign StickySelects_7_io_ins_2 = io_rPort_3_en_0 & _T_1069; // @[MemPrimitives.scala 125:64:@13687.4]
  assign StickySelects_7_io_ins_3 = io_rPort_5_en_0 & _T_1075; // @[MemPrimitives.scala 125:64:@13688.4]
  assign StickySelects_7_io_ins_4 = io_rPort_9_en_0 & _T_1081; // @[MemPrimitives.scala 125:64:@13689.4]
  assign StickySelects_7_io_ins_5 = io_rPort_11_en_0 & _T_1087; // @[MemPrimitives.scala 125:64:@13690.4]
  assign StickySelects_8_clock = clock; // @[:@13745.4]
  assign StickySelects_8_reset = reset; // @[:@13746.4]
  assign StickySelects_8_io_ins_0 = io_rPort_2_en_0 & _T_1119; // @[MemPrimitives.scala 125:64:@13747.4]
  assign StickySelects_8_io_ins_1 = io_rPort_4_en_0 & _T_1125; // @[MemPrimitives.scala 125:64:@13748.4]
  assign StickySelects_8_io_ins_2 = io_rPort_6_en_0 & _T_1131; // @[MemPrimitives.scala 125:64:@13749.4]
  assign StickySelects_8_io_ins_3 = io_rPort_7_en_0 & _T_1137; // @[MemPrimitives.scala 125:64:@13750.4]
  assign StickySelects_8_io_ins_4 = io_rPort_8_en_0 & _T_1143; // @[MemPrimitives.scala 125:64:@13751.4]
  assign StickySelects_8_io_ins_5 = io_rPort_10_en_0 & _T_1149; // @[MemPrimitives.scala 125:64:@13752.4]
  assign StickySelects_9_clock = clock; // @[:@13807.4]
  assign StickySelects_9_reset = reset; // @[:@13808.4]
  assign StickySelects_9_io_ins_0 = io_rPort_0_en_0 & _T_1181; // @[MemPrimitives.scala 125:64:@13809.4]
  assign StickySelects_9_io_ins_1 = io_rPort_1_en_0 & _T_1187; // @[MemPrimitives.scala 125:64:@13810.4]
  assign StickySelects_9_io_ins_2 = io_rPort_3_en_0 & _T_1193; // @[MemPrimitives.scala 125:64:@13811.4]
  assign StickySelects_9_io_ins_3 = io_rPort_5_en_0 & _T_1199; // @[MemPrimitives.scala 125:64:@13812.4]
  assign StickySelects_9_io_ins_4 = io_rPort_9_en_0 & _T_1205; // @[MemPrimitives.scala 125:64:@13813.4]
  assign StickySelects_9_io_ins_5 = io_rPort_11_en_0 & _T_1211; // @[MemPrimitives.scala 125:64:@13814.4]
  assign StickySelects_10_clock = clock; // @[:@13869.4]
  assign StickySelects_10_reset = reset; // @[:@13870.4]
  assign StickySelects_10_io_ins_0 = io_rPort_2_en_0 & _T_1243; // @[MemPrimitives.scala 125:64:@13871.4]
  assign StickySelects_10_io_ins_1 = io_rPort_4_en_0 & _T_1249; // @[MemPrimitives.scala 125:64:@13872.4]
  assign StickySelects_10_io_ins_2 = io_rPort_6_en_0 & _T_1255; // @[MemPrimitives.scala 125:64:@13873.4]
  assign StickySelects_10_io_ins_3 = io_rPort_7_en_0 & _T_1261; // @[MemPrimitives.scala 125:64:@13874.4]
  assign StickySelects_10_io_ins_4 = io_rPort_8_en_0 & _T_1267; // @[MemPrimitives.scala 125:64:@13875.4]
  assign StickySelects_10_io_ins_5 = io_rPort_10_en_0 & _T_1273; // @[MemPrimitives.scala 125:64:@13876.4]
  assign StickySelects_11_clock = clock; // @[:@13931.4]
  assign StickySelects_11_reset = reset; // @[:@13932.4]
  assign StickySelects_11_io_ins_0 = io_rPort_0_en_0 & _T_1305; // @[MemPrimitives.scala 125:64:@13933.4]
  assign StickySelects_11_io_ins_1 = io_rPort_1_en_0 & _T_1311; // @[MemPrimitives.scala 125:64:@13934.4]
  assign StickySelects_11_io_ins_2 = io_rPort_3_en_0 & _T_1317; // @[MemPrimitives.scala 125:64:@13935.4]
  assign StickySelects_11_io_ins_3 = io_rPort_5_en_0 & _T_1323; // @[MemPrimitives.scala 125:64:@13936.4]
  assign StickySelects_11_io_ins_4 = io_rPort_9_en_0 & _T_1329; // @[MemPrimitives.scala 125:64:@13937.4]
  assign StickySelects_11_io_ins_5 = io_rPort_11_en_0 & _T_1335; // @[MemPrimitives.scala 125:64:@13938.4]
  assign StickySelects_12_clock = clock; // @[:@13993.4]
  assign StickySelects_12_reset = reset; // @[:@13994.4]
  assign StickySelects_12_io_ins_0 = io_rPort_2_en_0 & _T_1367; // @[MemPrimitives.scala 125:64:@13995.4]
  assign StickySelects_12_io_ins_1 = io_rPort_4_en_0 & _T_1373; // @[MemPrimitives.scala 125:64:@13996.4]
  assign StickySelects_12_io_ins_2 = io_rPort_6_en_0 & _T_1379; // @[MemPrimitives.scala 125:64:@13997.4]
  assign StickySelects_12_io_ins_3 = io_rPort_7_en_0 & _T_1385; // @[MemPrimitives.scala 125:64:@13998.4]
  assign StickySelects_12_io_ins_4 = io_rPort_8_en_0 & _T_1391; // @[MemPrimitives.scala 125:64:@13999.4]
  assign StickySelects_12_io_ins_5 = io_rPort_10_en_0 & _T_1397; // @[MemPrimitives.scala 125:64:@14000.4]
  assign StickySelects_13_clock = clock; // @[:@14055.4]
  assign StickySelects_13_reset = reset; // @[:@14056.4]
  assign StickySelects_13_io_ins_0 = io_rPort_0_en_0 & _T_1429; // @[MemPrimitives.scala 125:64:@14057.4]
  assign StickySelects_13_io_ins_1 = io_rPort_1_en_0 & _T_1435; // @[MemPrimitives.scala 125:64:@14058.4]
  assign StickySelects_13_io_ins_2 = io_rPort_3_en_0 & _T_1441; // @[MemPrimitives.scala 125:64:@14059.4]
  assign StickySelects_13_io_ins_3 = io_rPort_5_en_0 & _T_1447; // @[MemPrimitives.scala 125:64:@14060.4]
  assign StickySelects_13_io_ins_4 = io_rPort_9_en_0 & _T_1453; // @[MemPrimitives.scala 125:64:@14061.4]
  assign StickySelects_13_io_ins_5 = io_rPort_11_en_0 & _T_1459; // @[MemPrimitives.scala 125:64:@14062.4]
  assign StickySelects_14_clock = clock; // @[:@14117.4]
  assign StickySelects_14_reset = reset; // @[:@14118.4]
  assign StickySelects_14_io_ins_0 = io_rPort_2_en_0 & _T_1491; // @[MemPrimitives.scala 125:64:@14119.4]
  assign StickySelects_14_io_ins_1 = io_rPort_4_en_0 & _T_1497; // @[MemPrimitives.scala 125:64:@14120.4]
  assign StickySelects_14_io_ins_2 = io_rPort_6_en_0 & _T_1503; // @[MemPrimitives.scala 125:64:@14121.4]
  assign StickySelects_14_io_ins_3 = io_rPort_7_en_0 & _T_1509; // @[MemPrimitives.scala 125:64:@14122.4]
  assign StickySelects_14_io_ins_4 = io_rPort_8_en_0 & _T_1515; // @[MemPrimitives.scala 125:64:@14123.4]
  assign StickySelects_14_io_ins_5 = io_rPort_10_en_0 & _T_1521; // @[MemPrimitives.scala 125:64:@14124.4]
  assign StickySelects_15_clock = clock; // @[:@14179.4]
  assign StickySelects_15_reset = reset; // @[:@14180.4]
  assign StickySelects_15_io_ins_0 = io_rPort_0_en_0 & _T_1553; // @[MemPrimitives.scala 125:64:@14181.4]
  assign StickySelects_15_io_ins_1 = io_rPort_1_en_0 & _T_1559; // @[MemPrimitives.scala 125:64:@14182.4]
  assign StickySelects_15_io_ins_2 = io_rPort_3_en_0 & _T_1565; // @[MemPrimitives.scala 125:64:@14183.4]
  assign StickySelects_15_io_ins_3 = io_rPort_5_en_0 & _T_1571; // @[MemPrimitives.scala 125:64:@14184.4]
  assign StickySelects_15_io_ins_4 = io_rPort_9_en_0 & _T_1577; // @[MemPrimitives.scala 125:64:@14185.4]
  assign StickySelects_15_io_ins_5 = io_rPort_11_en_0 & _T_1583; // @[MemPrimitives.scala 125:64:@14186.4]
  assign RetimeWrapper_clock = clock; // @[:@14242.4]
  assign RetimeWrapper_reset = reset; // @[:@14243.4]
  assign RetimeWrapper_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14245.4]
  assign RetimeWrapper_io_in = _T_685 & io_rPort_0_en_0; // @[package.scala 94:16:@14244.4]
  assign RetimeWrapper_1_clock = clock; // @[:@14250.4]
  assign RetimeWrapper_1_reset = reset; // @[:@14251.4]
  assign RetimeWrapper_1_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14253.4]
  assign RetimeWrapper_1_io_in = _T_809 & io_rPort_0_en_0; // @[package.scala 94:16:@14252.4]
  assign RetimeWrapper_2_clock = clock; // @[:@14258.4]
  assign RetimeWrapper_2_reset = reset; // @[:@14259.4]
  assign RetimeWrapper_2_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14261.4]
  assign RetimeWrapper_2_io_in = _T_933 & io_rPort_0_en_0; // @[package.scala 94:16:@14260.4]
  assign RetimeWrapper_3_clock = clock; // @[:@14266.4]
  assign RetimeWrapper_3_reset = reset; // @[:@14267.4]
  assign RetimeWrapper_3_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14269.4]
  assign RetimeWrapper_3_io_in = _T_1057 & io_rPort_0_en_0; // @[package.scala 94:16:@14268.4]
  assign RetimeWrapper_4_clock = clock; // @[:@14274.4]
  assign RetimeWrapper_4_reset = reset; // @[:@14275.4]
  assign RetimeWrapper_4_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14277.4]
  assign RetimeWrapper_4_io_in = _T_1181 & io_rPort_0_en_0; // @[package.scala 94:16:@14276.4]
  assign RetimeWrapper_5_clock = clock; // @[:@14282.4]
  assign RetimeWrapper_5_reset = reset; // @[:@14283.4]
  assign RetimeWrapper_5_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14285.4]
  assign RetimeWrapper_5_io_in = _T_1305 & io_rPort_0_en_0; // @[package.scala 94:16:@14284.4]
  assign RetimeWrapper_6_clock = clock; // @[:@14290.4]
  assign RetimeWrapper_6_reset = reset; // @[:@14291.4]
  assign RetimeWrapper_6_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14293.4]
  assign RetimeWrapper_6_io_in = _T_1429 & io_rPort_0_en_0; // @[package.scala 94:16:@14292.4]
  assign RetimeWrapper_7_clock = clock; // @[:@14298.4]
  assign RetimeWrapper_7_reset = reset; // @[:@14299.4]
  assign RetimeWrapper_7_io_flow = io_rPort_0_backpressure; // @[package.scala 95:18:@14301.4]
  assign RetimeWrapper_7_io_in = _T_1553 & io_rPort_0_en_0; // @[package.scala 94:16:@14300.4]
  assign RetimeWrapper_8_clock = clock; // @[:@14338.4]
  assign RetimeWrapper_8_reset = reset; // @[:@14339.4]
  assign RetimeWrapper_8_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14341.4]
  assign RetimeWrapper_8_io_in = _T_691 & io_rPort_1_en_0; // @[package.scala 94:16:@14340.4]
  assign RetimeWrapper_9_clock = clock; // @[:@14346.4]
  assign RetimeWrapper_9_reset = reset; // @[:@14347.4]
  assign RetimeWrapper_9_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14349.4]
  assign RetimeWrapper_9_io_in = _T_815 & io_rPort_1_en_0; // @[package.scala 94:16:@14348.4]
  assign RetimeWrapper_10_clock = clock; // @[:@14354.4]
  assign RetimeWrapper_10_reset = reset; // @[:@14355.4]
  assign RetimeWrapper_10_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14357.4]
  assign RetimeWrapper_10_io_in = _T_939 & io_rPort_1_en_0; // @[package.scala 94:16:@14356.4]
  assign RetimeWrapper_11_clock = clock; // @[:@14362.4]
  assign RetimeWrapper_11_reset = reset; // @[:@14363.4]
  assign RetimeWrapper_11_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14365.4]
  assign RetimeWrapper_11_io_in = _T_1063 & io_rPort_1_en_0; // @[package.scala 94:16:@14364.4]
  assign RetimeWrapper_12_clock = clock; // @[:@14370.4]
  assign RetimeWrapper_12_reset = reset; // @[:@14371.4]
  assign RetimeWrapper_12_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14373.4]
  assign RetimeWrapper_12_io_in = _T_1187 & io_rPort_1_en_0; // @[package.scala 94:16:@14372.4]
  assign RetimeWrapper_13_clock = clock; // @[:@14378.4]
  assign RetimeWrapper_13_reset = reset; // @[:@14379.4]
  assign RetimeWrapper_13_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14381.4]
  assign RetimeWrapper_13_io_in = _T_1311 & io_rPort_1_en_0; // @[package.scala 94:16:@14380.4]
  assign RetimeWrapper_14_clock = clock; // @[:@14386.4]
  assign RetimeWrapper_14_reset = reset; // @[:@14387.4]
  assign RetimeWrapper_14_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14389.4]
  assign RetimeWrapper_14_io_in = _T_1435 & io_rPort_1_en_0; // @[package.scala 94:16:@14388.4]
  assign RetimeWrapper_15_clock = clock; // @[:@14394.4]
  assign RetimeWrapper_15_reset = reset; // @[:@14395.4]
  assign RetimeWrapper_15_io_flow = io_rPort_1_backpressure; // @[package.scala 95:18:@14397.4]
  assign RetimeWrapper_15_io_in = _T_1559 & io_rPort_1_en_0; // @[package.scala 94:16:@14396.4]
  assign RetimeWrapper_16_clock = clock; // @[:@14434.4]
  assign RetimeWrapper_16_reset = reset; // @[:@14435.4]
  assign RetimeWrapper_16_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14437.4]
  assign RetimeWrapper_16_io_in = _T_623 & io_rPort_2_en_0; // @[package.scala 94:16:@14436.4]
  assign RetimeWrapper_17_clock = clock; // @[:@14442.4]
  assign RetimeWrapper_17_reset = reset; // @[:@14443.4]
  assign RetimeWrapper_17_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14445.4]
  assign RetimeWrapper_17_io_in = _T_747 & io_rPort_2_en_0; // @[package.scala 94:16:@14444.4]
  assign RetimeWrapper_18_clock = clock; // @[:@14450.4]
  assign RetimeWrapper_18_reset = reset; // @[:@14451.4]
  assign RetimeWrapper_18_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14453.4]
  assign RetimeWrapper_18_io_in = _T_871 & io_rPort_2_en_0; // @[package.scala 94:16:@14452.4]
  assign RetimeWrapper_19_clock = clock; // @[:@14458.4]
  assign RetimeWrapper_19_reset = reset; // @[:@14459.4]
  assign RetimeWrapper_19_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14461.4]
  assign RetimeWrapper_19_io_in = _T_995 & io_rPort_2_en_0; // @[package.scala 94:16:@14460.4]
  assign RetimeWrapper_20_clock = clock; // @[:@14466.4]
  assign RetimeWrapper_20_reset = reset; // @[:@14467.4]
  assign RetimeWrapper_20_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14469.4]
  assign RetimeWrapper_20_io_in = _T_1119 & io_rPort_2_en_0; // @[package.scala 94:16:@14468.4]
  assign RetimeWrapper_21_clock = clock; // @[:@14474.4]
  assign RetimeWrapper_21_reset = reset; // @[:@14475.4]
  assign RetimeWrapper_21_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14477.4]
  assign RetimeWrapper_21_io_in = _T_1243 & io_rPort_2_en_0; // @[package.scala 94:16:@14476.4]
  assign RetimeWrapper_22_clock = clock; // @[:@14482.4]
  assign RetimeWrapper_22_reset = reset; // @[:@14483.4]
  assign RetimeWrapper_22_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14485.4]
  assign RetimeWrapper_22_io_in = _T_1367 & io_rPort_2_en_0; // @[package.scala 94:16:@14484.4]
  assign RetimeWrapper_23_clock = clock; // @[:@14490.4]
  assign RetimeWrapper_23_reset = reset; // @[:@14491.4]
  assign RetimeWrapper_23_io_flow = io_rPort_2_backpressure; // @[package.scala 95:18:@14493.4]
  assign RetimeWrapper_23_io_in = _T_1491 & io_rPort_2_en_0; // @[package.scala 94:16:@14492.4]
  assign RetimeWrapper_24_clock = clock; // @[:@14530.4]
  assign RetimeWrapper_24_reset = reset; // @[:@14531.4]
  assign RetimeWrapper_24_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14533.4]
  assign RetimeWrapper_24_io_in = _T_697 & io_rPort_3_en_0; // @[package.scala 94:16:@14532.4]
  assign RetimeWrapper_25_clock = clock; // @[:@14538.4]
  assign RetimeWrapper_25_reset = reset; // @[:@14539.4]
  assign RetimeWrapper_25_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14541.4]
  assign RetimeWrapper_25_io_in = _T_821 & io_rPort_3_en_0; // @[package.scala 94:16:@14540.4]
  assign RetimeWrapper_26_clock = clock; // @[:@14546.4]
  assign RetimeWrapper_26_reset = reset; // @[:@14547.4]
  assign RetimeWrapper_26_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14549.4]
  assign RetimeWrapper_26_io_in = _T_945 & io_rPort_3_en_0; // @[package.scala 94:16:@14548.4]
  assign RetimeWrapper_27_clock = clock; // @[:@14554.4]
  assign RetimeWrapper_27_reset = reset; // @[:@14555.4]
  assign RetimeWrapper_27_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14557.4]
  assign RetimeWrapper_27_io_in = _T_1069 & io_rPort_3_en_0; // @[package.scala 94:16:@14556.4]
  assign RetimeWrapper_28_clock = clock; // @[:@14562.4]
  assign RetimeWrapper_28_reset = reset; // @[:@14563.4]
  assign RetimeWrapper_28_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14565.4]
  assign RetimeWrapper_28_io_in = _T_1193 & io_rPort_3_en_0; // @[package.scala 94:16:@14564.4]
  assign RetimeWrapper_29_clock = clock; // @[:@14570.4]
  assign RetimeWrapper_29_reset = reset; // @[:@14571.4]
  assign RetimeWrapper_29_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14573.4]
  assign RetimeWrapper_29_io_in = _T_1317 & io_rPort_3_en_0; // @[package.scala 94:16:@14572.4]
  assign RetimeWrapper_30_clock = clock; // @[:@14578.4]
  assign RetimeWrapper_30_reset = reset; // @[:@14579.4]
  assign RetimeWrapper_30_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14581.4]
  assign RetimeWrapper_30_io_in = _T_1441 & io_rPort_3_en_0; // @[package.scala 94:16:@14580.4]
  assign RetimeWrapper_31_clock = clock; // @[:@14586.4]
  assign RetimeWrapper_31_reset = reset; // @[:@14587.4]
  assign RetimeWrapper_31_io_flow = io_rPort_3_backpressure; // @[package.scala 95:18:@14589.4]
  assign RetimeWrapper_31_io_in = _T_1565 & io_rPort_3_en_0; // @[package.scala 94:16:@14588.4]
  assign RetimeWrapper_32_clock = clock; // @[:@14626.4]
  assign RetimeWrapper_32_reset = reset; // @[:@14627.4]
  assign RetimeWrapper_32_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14629.4]
  assign RetimeWrapper_32_io_in = _T_629 & io_rPort_4_en_0; // @[package.scala 94:16:@14628.4]
  assign RetimeWrapper_33_clock = clock; // @[:@14634.4]
  assign RetimeWrapper_33_reset = reset; // @[:@14635.4]
  assign RetimeWrapper_33_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14637.4]
  assign RetimeWrapper_33_io_in = _T_753 & io_rPort_4_en_0; // @[package.scala 94:16:@14636.4]
  assign RetimeWrapper_34_clock = clock; // @[:@14642.4]
  assign RetimeWrapper_34_reset = reset; // @[:@14643.4]
  assign RetimeWrapper_34_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14645.4]
  assign RetimeWrapper_34_io_in = _T_877 & io_rPort_4_en_0; // @[package.scala 94:16:@14644.4]
  assign RetimeWrapper_35_clock = clock; // @[:@14650.4]
  assign RetimeWrapper_35_reset = reset; // @[:@14651.4]
  assign RetimeWrapper_35_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14653.4]
  assign RetimeWrapper_35_io_in = _T_1001 & io_rPort_4_en_0; // @[package.scala 94:16:@14652.4]
  assign RetimeWrapper_36_clock = clock; // @[:@14658.4]
  assign RetimeWrapper_36_reset = reset; // @[:@14659.4]
  assign RetimeWrapper_36_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14661.4]
  assign RetimeWrapper_36_io_in = _T_1125 & io_rPort_4_en_0; // @[package.scala 94:16:@14660.4]
  assign RetimeWrapper_37_clock = clock; // @[:@14666.4]
  assign RetimeWrapper_37_reset = reset; // @[:@14667.4]
  assign RetimeWrapper_37_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14669.4]
  assign RetimeWrapper_37_io_in = _T_1249 & io_rPort_4_en_0; // @[package.scala 94:16:@14668.4]
  assign RetimeWrapper_38_clock = clock; // @[:@14674.4]
  assign RetimeWrapper_38_reset = reset; // @[:@14675.4]
  assign RetimeWrapper_38_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14677.4]
  assign RetimeWrapper_38_io_in = _T_1373 & io_rPort_4_en_0; // @[package.scala 94:16:@14676.4]
  assign RetimeWrapper_39_clock = clock; // @[:@14682.4]
  assign RetimeWrapper_39_reset = reset; // @[:@14683.4]
  assign RetimeWrapper_39_io_flow = io_rPort_4_backpressure; // @[package.scala 95:18:@14685.4]
  assign RetimeWrapper_39_io_in = _T_1497 & io_rPort_4_en_0; // @[package.scala 94:16:@14684.4]
  assign RetimeWrapper_40_clock = clock; // @[:@14722.4]
  assign RetimeWrapper_40_reset = reset; // @[:@14723.4]
  assign RetimeWrapper_40_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14725.4]
  assign RetimeWrapper_40_io_in = _T_703 & io_rPort_5_en_0; // @[package.scala 94:16:@14724.4]
  assign RetimeWrapper_41_clock = clock; // @[:@14730.4]
  assign RetimeWrapper_41_reset = reset; // @[:@14731.4]
  assign RetimeWrapper_41_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14733.4]
  assign RetimeWrapper_41_io_in = _T_827 & io_rPort_5_en_0; // @[package.scala 94:16:@14732.4]
  assign RetimeWrapper_42_clock = clock; // @[:@14738.4]
  assign RetimeWrapper_42_reset = reset; // @[:@14739.4]
  assign RetimeWrapper_42_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14741.4]
  assign RetimeWrapper_42_io_in = _T_951 & io_rPort_5_en_0; // @[package.scala 94:16:@14740.4]
  assign RetimeWrapper_43_clock = clock; // @[:@14746.4]
  assign RetimeWrapper_43_reset = reset; // @[:@14747.4]
  assign RetimeWrapper_43_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14749.4]
  assign RetimeWrapper_43_io_in = _T_1075 & io_rPort_5_en_0; // @[package.scala 94:16:@14748.4]
  assign RetimeWrapper_44_clock = clock; // @[:@14754.4]
  assign RetimeWrapper_44_reset = reset; // @[:@14755.4]
  assign RetimeWrapper_44_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14757.4]
  assign RetimeWrapper_44_io_in = _T_1199 & io_rPort_5_en_0; // @[package.scala 94:16:@14756.4]
  assign RetimeWrapper_45_clock = clock; // @[:@14762.4]
  assign RetimeWrapper_45_reset = reset; // @[:@14763.4]
  assign RetimeWrapper_45_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14765.4]
  assign RetimeWrapper_45_io_in = _T_1323 & io_rPort_5_en_0; // @[package.scala 94:16:@14764.4]
  assign RetimeWrapper_46_clock = clock; // @[:@14770.4]
  assign RetimeWrapper_46_reset = reset; // @[:@14771.4]
  assign RetimeWrapper_46_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14773.4]
  assign RetimeWrapper_46_io_in = _T_1447 & io_rPort_5_en_0; // @[package.scala 94:16:@14772.4]
  assign RetimeWrapper_47_clock = clock; // @[:@14778.4]
  assign RetimeWrapper_47_reset = reset; // @[:@14779.4]
  assign RetimeWrapper_47_io_flow = io_rPort_5_backpressure; // @[package.scala 95:18:@14781.4]
  assign RetimeWrapper_47_io_in = _T_1571 & io_rPort_5_en_0; // @[package.scala 94:16:@14780.4]
  assign RetimeWrapper_48_clock = clock; // @[:@14818.4]
  assign RetimeWrapper_48_reset = reset; // @[:@14819.4]
  assign RetimeWrapper_48_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14821.4]
  assign RetimeWrapper_48_io_in = _T_635 & io_rPort_6_en_0; // @[package.scala 94:16:@14820.4]
  assign RetimeWrapper_49_clock = clock; // @[:@14826.4]
  assign RetimeWrapper_49_reset = reset; // @[:@14827.4]
  assign RetimeWrapper_49_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14829.4]
  assign RetimeWrapper_49_io_in = _T_759 & io_rPort_6_en_0; // @[package.scala 94:16:@14828.4]
  assign RetimeWrapper_50_clock = clock; // @[:@14834.4]
  assign RetimeWrapper_50_reset = reset; // @[:@14835.4]
  assign RetimeWrapper_50_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14837.4]
  assign RetimeWrapper_50_io_in = _T_883 & io_rPort_6_en_0; // @[package.scala 94:16:@14836.4]
  assign RetimeWrapper_51_clock = clock; // @[:@14842.4]
  assign RetimeWrapper_51_reset = reset; // @[:@14843.4]
  assign RetimeWrapper_51_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14845.4]
  assign RetimeWrapper_51_io_in = _T_1007 & io_rPort_6_en_0; // @[package.scala 94:16:@14844.4]
  assign RetimeWrapper_52_clock = clock; // @[:@14850.4]
  assign RetimeWrapper_52_reset = reset; // @[:@14851.4]
  assign RetimeWrapper_52_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14853.4]
  assign RetimeWrapper_52_io_in = _T_1131 & io_rPort_6_en_0; // @[package.scala 94:16:@14852.4]
  assign RetimeWrapper_53_clock = clock; // @[:@14858.4]
  assign RetimeWrapper_53_reset = reset; // @[:@14859.4]
  assign RetimeWrapper_53_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14861.4]
  assign RetimeWrapper_53_io_in = _T_1255 & io_rPort_6_en_0; // @[package.scala 94:16:@14860.4]
  assign RetimeWrapper_54_clock = clock; // @[:@14866.4]
  assign RetimeWrapper_54_reset = reset; // @[:@14867.4]
  assign RetimeWrapper_54_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14869.4]
  assign RetimeWrapper_54_io_in = _T_1379 & io_rPort_6_en_0; // @[package.scala 94:16:@14868.4]
  assign RetimeWrapper_55_clock = clock; // @[:@14874.4]
  assign RetimeWrapper_55_reset = reset; // @[:@14875.4]
  assign RetimeWrapper_55_io_flow = io_rPort_6_backpressure; // @[package.scala 95:18:@14877.4]
  assign RetimeWrapper_55_io_in = _T_1503 & io_rPort_6_en_0; // @[package.scala 94:16:@14876.4]
  assign RetimeWrapper_56_clock = clock; // @[:@14914.4]
  assign RetimeWrapper_56_reset = reset; // @[:@14915.4]
  assign RetimeWrapper_56_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14917.4]
  assign RetimeWrapper_56_io_in = _T_641 & io_rPort_7_en_0; // @[package.scala 94:16:@14916.4]
  assign RetimeWrapper_57_clock = clock; // @[:@14922.4]
  assign RetimeWrapper_57_reset = reset; // @[:@14923.4]
  assign RetimeWrapper_57_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14925.4]
  assign RetimeWrapper_57_io_in = _T_765 & io_rPort_7_en_0; // @[package.scala 94:16:@14924.4]
  assign RetimeWrapper_58_clock = clock; // @[:@14930.4]
  assign RetimeWrapper_58_reset = reset; // @[:@14931.4]
  assign RetimeWrapper_58_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14933.4]
  assign RetimeWrapper_58_io_in = _T_889 & io_rPort_7_en_0; // @[package.scala 94:16:@14932.4]
  assign RetimeWrapper_59_clock = clock; // @[:@14938.4]
  assign RetimeWrapper_59_reset = reset; // @[:@14939.4]
  assign RetimeWrapper_59_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14941.4]
  assign RetimeWrapper_59_io_in = _T_1013 & io_rPort_7_en_0; // @[package.scala 94:16:@14940.4]
  assign RetimeWrapper_60_clock = clock; // @[:@14946.4]
  assign RetimeWrapper_60_reset = reset; // @[:@14947.4]
  assign RetimeWrapper_60_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14949.4]
  assign RetimeWrapper_60_io_in = _T_1137 & io_rPort_7_en_0; // @[package.scala 94:16:@14948.4]
  assign RetimeWrapper_61_clock = clock; // @[:@14954.4]
  assign RetimeWrapper_61_reset = reset; // @[:@14955.4]
  assign RetimeWrapper_61_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14957.4]
  assign RetimeWrapper_61_io_in = _T_1261 & io_rPort_7_en_0; // @[package.scala 94:16:@14956.4]
  assign RetimeWrapper_62_clock = clock; // @[:@14962.4]
  assign RetimeWrapper_62_reset = reset; // @[:@14963.4]
  assign RetimeWrapper_62_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14965.4]
  assign RetimeWrapper_62_io_in = _T_1385 & io_rPort_7_en_0; // @[package.scala 94:16:@14964.4]
  assign RetimeWrapper_63_clock = clock; // @[:@14970.4]
  assign RetimeWrapper_63_reset = reset; // @[:@14971.4]
  assign RetimeWrapper_63_io_flow = io_rPort_7_backpressure; // @[package.scala 95:18:@14973.4]
  assign RetimeWrapper_63_io_in = _T_1509 & io_rPort_7_en_0; // @[package.scala 94:16:@14972.4]
  assign RetimeWrapper_64_clock = clock; // @[:@15010.4]
  assign RetimeWrapper_64_reset = reset; // @[:@15011.4]
  assign RetimeWrapper_64_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15013.4]
  assign RetimeWrapper_64_io_in = _T_647 & io_rPort_8_en_0; // @[package.scala 94:16:@15012.4]
  assign RetimeWrapper_65_clock = clock; // @[:@15018.4]
  assign RetimeWrapper_65_reset = reset; // @[:@15019.4]
  assign RetimeWrapper_65_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15021.4]
  assign RetimeWrapper_65_io_in = _T_771 & io_rPort_8_en_0; // @[package.scala 94:16:@15020.4]
  assign RetimeWrapper_66_clock = clock; // @[:@15026.4]
  assign RetimeWrapper_66_reset = reset; // @[:@15027.4]
  assign RetimeWrapper_66_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15029.4]
  assign RetimeWrapper_66_io_in = _T_895 & io_rPort_8_en_0; // @[package.scala 94:16:@15028.4]
  assign RetimeWrapper_67_clock = clock; // @[:@15034.4]
  assign RetimeWrapper_67_reset = reset; // @[:@15035.4]
  assign RetimeWrapper_67_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15037.4]
  assign RetimeWrapper_67_io_in = _T_1019 & io_rPort_8_en_0; // @[package.scala 94:16:@15036.4]
  assign RetimeWrapper_68_clock = clock; // @[:@15042.4]
  assign RetimeWrapper_68_reset = reset; // @[:@15043.4]
  assign RetimeWrapper_68_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15045.4]
  assign RetimeWrapper_68_io_in = _T_1143 & io_rPort_8_en_0; // @[package.scala 94:16:@15044.4]
  assign RetimeWrapper_69_clock = clock; // @[:@15050.4]
  assign RetimeWrapper_69_reset = reset; // @[:@15051.4]
  assign RetimeWrapper_69_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15053.4]
  assign RetimeWrapper_69_io_in = _T_1267 & io_rPort_8_en_0; // @[package.scala 94:16:@15052.4]
  assign RetimeWrapper_70_clock = clock; // @[:@15058.4]
  assign RetimeWrapper_70_reset = reset; // @[:@15059.4]
  assign RetimeWrapper_70_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15061.4]
  assign RetimeWrapper_70_io_in = _T_1391 & io_rPort_8_en_0; // @[package.scala 94:16:@15060.4]
  assign RetimeWrapper_71_clock = clock; // @[:@15066.4]
  assign RetimeWrapper_71_reset = reset; // @[:@15067.4]
  assign RetimeWrapper_71_io_flow = io_rPort_8_backpressure; // @[package.scala 95:18:@15069.4]
  assign RetimeWrapper_71_io_in = _T_1515 & io_rPort_8_en_0; // @[package.scala 94:16:@15068.4]
  assign RetimeWrapper_72_clock = clock; // @[:@15106.4]
  assign RetimeWrapper_72_reset = reset; // @[:@15107.4]
  assign RetimeWrapper_72_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15109.4]
  assign RetimeWrapper_72_io_in = _T_709 & io_rPort_9_en_0; // @[package.scala 94:16:@15108.4]
  assign RetimeWrapper_73_clock = clock; // @[:@15114.4]
  assign RetimeWrapper_73_reset = reset; // @[:@15115.4]
  assign RetimeWrapper_73_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15117.4]
  assign RetimeWrapper_73_io_in = _T_833 & io_rPort_9_en_0; // @[package.scala 94:16:@15116.4]
  assign RetimeWrapper_74_clock = clock; // @[:@15122.4]
  assign RetimeWrapper_74_reset = reset; // @[:@15123.4]
  assign RetimeWrapper_74_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15125.4]
  assign RetimeWrapper_74_io_in = _T_957 & io_rPort_9_en_0; // @[package.scala 94:16:@15124.4]
  assign RetimeWrapper_75_clock = clock; // @[:@15130.4]
  assign RetimeWrapper_75_reset = reset; // @[:@15131.4]
  assign RetimeWrapper_75_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15133.4]
  assign RetimeWrapper_75_io_in = _T_1081 & io_rPort_9_en_0; // @[package.scala 94:16:@15132.4]
  assign RetimeWrapper_76_clock = clock; // @[:@15138.4]
  assign RetimeWrapper_76_reset = reset; // @[:@15139.4]
  assign RetimeWrapper_76_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15141.4]
  assign RetimeWrapper_76_io_in = _T_1205 & io_rPort_9_en_0; // @[package.scala 94:16:@15140.4]
  assign RetimeWrapper_77_clock = clock; // @[:@15146.4]
  assign RetimeWrapper_77_reset = reset; // @[:@15147.4]
  assign RetimeWrapper_77_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15149.4]
  assign RetimeWrapper_77_io_in = _T_1329 & io_rPort_9_en_0; // @[package.scala 94:16:@15148.4]
  assign RetimeWrapper_78_clock = clock; // @[:@15154.4]
  assign RetimeWrapper_78_reset = reset; // @[:@15155.4]
  assign RetimeWrapper_78_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15157.4]
  assign RetimeWrapper_78_io_in = _T_1453 & io_rPort_9_en_0; // @[package.scala 94:16:@15156.4]
  assign RetimeWrapper_79_clock = clock; // @[:@15162.4]
  assign RetimeWrapper_79_reset = reset; // @[:@15163.4]
  assign RetimeWrapper_79_io_flow = io_rPort_9_backpressure; // @[package.scala 95:18:@15165.4]
  assign RetimeWrapper_79_io_in = _T_1577 & io_rPort_9_en_0; // @[package.scala 94:16:@15164.4]
  assign RetimeWrapper_80_clock = clock; // @[:@15202.4]
  assign RetimeWrapper_80_reset = reset; // @[:@15203.4]
  assign RetimeWrapper_80_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15205.4]
  assign RetimeWrapper_80_io_in = _T_653 & io_rPort_10_en_0; // @[package.scala 94:16:@15204.4]
  assign RetimeWrapper_81_clock = clock; // @[:@15210.4]
  assign RetimeWrapper_81_reset = reset; // @[:@15211.4]
  assign RetimeWrapper_81_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15213.4]
  assign RetimeWrapper_81_io_in = _T_777 & io_rPort_10_en_0; // @[package.scala 94:16:@15212.4]
  assign RetimeWrapper_82_clock = clock; // @[:@15218.4]
  assign RetimeWrapper_82_reset = reset; // @[:@15219.4]
  assign RetimeWrapper_82_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15221.4]
  assign RetimeWrapper_82_io_in = _T_901 & io_rPort_10_en_0; // @[package.scala 94:16:@15220.4]
  assign RetimeWrapper_83_clock = clock; // @[:@15226.4]
  assign RetimeWrapper_83_reset = reset; // @[:@15227.4]
  assign RetimeWrapper_83_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15229.4]
  assign RetimeWrapper_83_io_in = _T_1025 & io_rPort_10_en_0; // @[package.scala 94:16:@15228.4]
  assign RetimeWrapper_84_clock = clock; // @[:@15234.4]
  assign RetimeWrapper_84_reset = reset; // @[:@15235.4]
  assign RetimeWrapper_84_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15237.4]
  assign RetimeWrapper_84_io_in = _T_1149 & io_rPort_10_en_0; // @[package.scala 94:16:@15236.4]
  assign RetimeWrapper_85_clock = clock; // @[:@15242.4]
  assign RetimeWrapper_85_reset = reset; // @[:@15243.4]
  assign RetimeWrapper_85_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15245.4]
  assign RetimeWrapper_85_io_in = _T_1273 & io_rPort_10_en_0; // @[package.scala 94:16:@15244.4]
  assign RetimeWrapper_86_clock = clock; // @[:@15250.4]
  assign RetimeWrapper_86_reset = reset; // @[:@15251.4]
  assign RetimeWrapper_86_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15253.4]
  assign RetimeWrapper_86_io_in = _T_1397 & io_rPort_10_en_0; // @[package.scala 94:16:@15252.4]
  assign RetimeWrapper_87_clock = clock; // @[:@15258.4]
  assign RetimeWrapper_87_reset = reset; // @[:@15259.4]
  assign RetimeWrapper_87_io_flow = io_rPort_10_backpressure; // @[package.scala 95:18:@15261.4]
  assign RetimeWrapper_87_io_in = _T_1521 & io_rPort_10_en_0; // @[package.scala 94:16:@15260.4]
  assign RetimeWrapper_88_clock = clock; // @[:@15298.4]
  assign RetimeWrapper_88_reset = reset; // @[:@15299.4]
  assign RetimeWrapper_88_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15301.4]
  assign RetimeWrapper_88_io_in = _T_715 & io_rPort_11_en_0; // @[package.scala 94:16:@15300.4]
  assign RetimeWrapper_89_clock = clock; // @[:@15306.4]
  assign RetimeWrapper_89_reset = reset; // @[:@15307.4]
  assign RetimeWrapper_89_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15309.4]
  assign RetimeWrapper_89_io_in = _T_839 & io_rPort_11_en_0; // @[package.scala 94:16:@15308.4]
  assign RetimeWrapper_90_clock = clock; // @[:@15314.4]
  assign RetimeWrapper_90_reset = reset; // @[:@15315.4]
  assign RetimeWrapper_90_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15317.4]
  assign RetimeWrapper_90_io_in = _T_963 & io_rPort_11_en_0; // @[package.scala 94:16:@15316.4]
  assign RetimeWrapper_91_clock = clock; // @[:@15322.4]
  assign RetimeWrapper_91_reset = reset; // @[:@15323.4]
  assign RetimeWrapper_91_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15325.4]
  assign RetimeWrapper_91_io_in = _T_1087 & io_rPort_11_en_0; // @[package.scala 94:16:@15324.4]
  assign RetimeWrapper_92_clock = clock; // @[:@15330.4]
  assign RetimeWrapper_92_reset = reset; // @[:@15331.4]
  assign RetimeWrapper_92_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15333.4]
  assign RetimeWrapper_92_io_in = _T_1211 & io_rPort_11_en_0; // @[package.scala 94:16:@15332.4]
  assign RetimeWrapper_93_clock = clock; // @[:@15338.4]
  assign RetimeWrapper_93_reset = reset; // @[:@15339.4]
  assign RetimeWrapper_93_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15341.4]
  assign RetimeWrapper_93_io_in = _T_1335 & io_rPort_11_en_0; // @[package.scala 94:16:@15340.4]
  assign RetimeWrapper_94_clock = clock; // @[:@15346.4]
  assign RetimeWrapper_94_reset = reset; // @[:@15347.4]
  assign RetimeWrapper_94_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15349.4]
  assign RetimeWrapper_94_io_in = _T_1459 & io_rPort_11_en_0; // @[package.scala 94:16:@15348.4]
  assign RetimeWrapper_95_clock = clock; // @[:@15354.4]
  assign RetimeWrapper_95_reset = reset; // @[:@15355.4]
  assign RetimeWrapper_95_io_flow = io_rPort_11_backpressure; // @[package.scala 95:18:@15357.4]
  assign RetimeWrapper_95_io_in = _T_1583 & io_rPort_11_en_0; // @[package.scala 94:16:@15356.4]
endmodule
module RetimeWrapper_168( // @[:@15772.2]
  input         clock, // @[:@15773.4]
  input         reset, // @[:@15774.4]
  input         io_flow, // @[:@15775.4]
  input  [31:0] io_in, // @[:@15775.4]
  output [31:0] io_out // @[:@15775.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15777.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@15777.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15790.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15789.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15788.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15787.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15786.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15784.4]
endmodule
module RetimeWrapper_169( // @[:@15804.2]
  input         clock, // @[:@15805.4]
  input         reset, // @[:@15806.4]
  input         io_flow, // @[:@15807.4]
  input  [31:0] io_in, // @[:@15807.4]
  output [31:0] io_out // @[:@15807.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15809.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(2)) sr ( // @[RetimeShiftRegister.scala 15:20:@15809.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15822.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15821.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@15820.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15819.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15818.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15816.4]
endmodule
module RetimeWrapper_172( // @[:@15900.2]
  input   clock, // @[:@15901.4]
  input   reset, // @[:@15902.4]
  input   io_flow, // @[:@15903.4]
  input   io_in, // @[:@15903.4]
  output  io_out // @[:@15903.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@15905.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@15905.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@15905.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@15905.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@15905.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@15905.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@15905.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@15918.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@15917.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@15916.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@15915.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@15914.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@15912.4]
endmodule
module RetimeWrapper_181( // @[:@16482.2]
  input         clock, // @[:@16483.4]
  input         reset, // @[:@16484.4]
  input         io_flow, // @[:@16485.4]
  input  [31:0] io_in, // @[:@16485.4]
  output [31:0] io_out // @[:@16485.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16487.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(6)) sr ( // @[RetimeShiftRegister.scala 15:20:@16487.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16500.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16499.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16498.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16497.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16496.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16494.4]
endmodule
module RetimeWrapper_184( // @[:@16578.2]
  input         clock, // @[:@16579.4]
  input         reset, // @[:@16580.4]
  input         io_flow, // @[:@16581.4]
  input  [31:0] io_in, // @[:@16581.4]
  output [31:0] io_out // @[:@16581.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16583.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@16583.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16596.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16595.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16594.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16593.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16592.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16590.4]
endmodule
module RetimeWrapper_186( // @[:@16642.2]
  input   clock, // @[:@16643.4]
  input   reset, // @[:@16644.4]
  input   io_flow, // @[:@16645.4]
  input   io_in, // @[:@16645.4]
  output  io_out // @[:@16645.4]
);
  wire  sr_out; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_in; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_init; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16647.4]
  RetimeShiftRegister #(.WIDTH(1), .STAGES(9)) sr ( // @[RetimeShiftRegister.scala 15:20:@16647.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16660.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16659.4]
  assign sr_init = 1'h0; // @[RetimeShiftRegister.scala 19:16:@16658.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16657.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16656.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16654.4]
endmodule
module RetimeWrapper_187( // @[:@16674.2]
  input         clock, // @[:@16675.4]
  input         reset, // @[:@16676.4]
  input         io_flow, // @[:@16677.4]
  input  [31:0] io_in, // @[:@16677.4]
  output [31:0] io_out // @[:@16677.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16679.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(8)) sr ( // @[RetimeShiftRegister.scala 15:20:@16679.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16692.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16691.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16690.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16689.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16688.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16686.4]
endmodule
module RetimeWrapper_188( // @[:@16706.2]
  input         clock, // @[:@16707.4]
  input         reset, // @[:@16708.4]
  input         io_flow, // @[:@16709.4]
  input  [31:0] io_in, // @[:@16709.4]
  output [31:0] io_out // @[:@16709.4]
);
  wire [31:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@16711.4]
  wire [31:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@16711.4]
  wire [31:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@16711.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@16711.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@16711.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@16711.4]
  RetimeShiftRegister #(.WIDTH(32), .STAGES(7)) sr ( // @[RetimeShiftRegister.scala 15:20:@16711.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@16724.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@16723.4]
  assign sr_init = 32'h0; // @[RetimeShiftRegister.scala 19:16:@16722.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@16721.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@16720.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@16718.4]
endmodule
module Multiplier( // @[:@20852.2]
  input         clock, // @[:@20853.4]
  input         io_flow, // @[:@20855.4]
  input  [31:0] io_a, // @[:@20855.4]
  input  [31:0] io_b, // @[:@20855.4]
  output [31:0] io_out // @[:@20855.4]
);
  wire [31:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  wire [31:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  wire [31:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@20857.4]
  mul_32_32_32_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@20857.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@20867.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@20865.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@20864.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@20866.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@20863.4]
endmodule
module x357( // @[:@20887.2]
  input         clock, // @[:@20888.4]
  input  [31:0] io_a, // @[:@20890.4]
  input  [31:0] io_b, // @[:@20890.4]
  input         io_flow, // @[:@20890.4]
  output [31:0] io_result // @[:@20890.4]
);
  wire  x357_clock; // @[BigIPZynq.scala 63:21:@20897.4]
  wire  x357_io_flow; // @[BigIPZynq.scala 63:21:@20897.4]
  wire [31:0] x357_io_a; // @[BigIPZynq.scala 63:21:@20897.4]
  wire [31:0] x357_io_b; // @[BigIPZynq.scala 63:21:@20897.4]
  wire [31:0] x357_io_out; // @[BigIPZynq.scala 63:21:@20897.4]
  wire [31:0] fix2fixBox_io_a; // @[Math.scala 253:30:@20906.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@20906.4]
  Multiplier x357 ( // @[BigIPZynq.scala 63:21:@20897.4]
    .clock(x357_clock),
    .io_flow(x357_io_flow),
    .io_a(x357_io_a),
    .io_b(x357_io_b),
    .io_out(x357_io_out)
  );
  fix2fixBox fix2fixBox ( // @[Math.scala 253:30:@20906.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@20914.4]
  assign x357_clock = clock; // @[:@20898.4]
  assign x357_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@20902.4]
  assign x357_io_a = io_a; // @[BigIPZynq.scala 64:14:@20900.4]
  assign x357_io_b = io_b; // @[BigIPZynq.scala 65:14:@20901.4]
  assign fix2fixBox_io_a = x357_io_out; // @[Math.scala 254:23:@20909.4]
endmodule
module fix2fixBox_93( // @[:@21508.2]
  input  [31:0] io_a, // @[:@21511.4]
  output [32:0] io_b // @[:@21511.4]
);
  assign io_b = {1'h0,io_a}; // @[Converter.scala 95:38:@21525.4]
endmodule
module __56( // @[:@21527.2]
  input  [31:0] io_b, // @[:@21530.4]
  output [32:0] io_result // @[:@21530.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@21535.4]
  wire [32:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@21535.4]
  fix2fixBox_93 fix2fixBox ( // @[BigIPZynq.scala 219:30:@21535.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@21543.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@21538.4]
endmodule
module x366_x3( // @[:@21639.2]
  input         clock, // @[:@21640.4]
  input         reset, // @[:@21641.4]
  input  [31:0] io_a, // @[:@21642.4]
  input  [31:0] io_b, // @[:@21642.4]
  input         io_flow, // @[:@21642.4]
  output [31:0] io_result // @[:@21642.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@21650.4]
  wire [32:0] __io_result; // @[Math.scala 720:24:@21650.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@21657.4]
  wire [32:0] __1_io_result; // @[Math.scala 720:24:@21657.4]
  wire  fix2fixBox_clock; // @[Math.scala 141:30:@21667.4]
  wire  fix2fixBox_reset; // @[Math.scala 141:30:@21667.4]
  wire [32:0] fix2fixBox_io_a; // @[Math.scala 141:30:@21667.4]
  wire  fix2fixBox_io_flow; // @[Math.scala 141:30:@21667.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 141:30:@21667.4]
  wire [32:0] a_upcast_number; // @[Math.scala 723:22:@21655.4 Math.scala 724:14:@21656.4]
  wire [32:0] b_upcast_number; // @[Math.scala 723:22:@21662.4 Math.scala 724:14:@21663.4]
  wire [33:0] _T_21; // @[Math.scala 136:37:@21664.4]
  __56 _ ( // @[Math.scala 720:24:@21650.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  __56 __1 ( // @[Math.scala 720:24:@21657.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  fix2fixBox_4 fix2fixBox ( // @[Math.scala 141:30:@21667.4]
    .clock(fix2fixBox_clock),
    .reset(fix2fixBox_reset),
    .io_a(fix2fixBox_io_a),
    .io_flow(fix2fixBox_io_flow),
    .io_b(fix2fixBox_io_b)
  );
  assign a_upcast_number = __io_result; // @[Math.scala 723:22:@21655.4 Math.scala 724:14:@21656.4]
  assign b_upcast_number = __1_io_result; // @[Math.scala 723:22:@21662.4 Math.scala 724:14:@21663.4]
  assign _T_21 = a_upcast_number + b_upcast_number; // @[Math.scala 136:37:@21664.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 147:17:@21675.4]
  assign __io_b = io_a; // @[Math.scala 721:17:@21653.4]
  assign __1_io_b = io_b; // @[Math.scala 721:17:@21660.4]
  assign fix2fixBox_clock = clock; // @[:@21668.4]
  assign fix2fixBox_reset = reset; // @[:@21669.4]
  assign fix2fixBox_io_a = a_upcast_number + b_upcast_number; // @[Math.scala 142:23:@21670.4]
  assign fix2fixBox_io_flow = io_flow; // @[Math.scala 145:26:@21673.4]
endmodule
module fix2fixBox_117( // @[:@22892.2]
  input  [31:0] io_a, // @[:@22895.4]
  output [31:0] io_b // @[:@22895.4]
);
  wire [24:0] new_dec; // @[Converter.scala 63:26:@22905.4]
  assign new_dec = io_a[24:0]; // @[Converter.scala 63:26:@22905.4]
  assign io_b = {new_dec,7'h0}; // @[Converter.scala 94:38:@22908.4]
endmodule
module x374( // @[:@22910.2]
  input  [31:0] io_b, // @[:@22913.4]
  output [31:0] io_result // @[:@22913.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@22918.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@22918.4]
  fix2fixBox_117 fix2fixBox ( // @[BigIPZynq.scala 219:30:@22918.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@22926.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@22921.4]
endmodule
module Multiplier_9( // @[:@22938.2]
  input         clock, // @[:@22939.4]
  input         io_flow, // @[:@22941.4]
  input  [38:0] io_a, // @[:@22941.4]
  input  [38:0] io_b, // @[:@22941.4]
  output [38:0] io_out // @[:@22941.4]
);
  wire [38:0] m_P; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  wire [38:0] m_B; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  wire [38:0] m_A; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  wire  m_CE; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  wire  m_CLK; // @[ZynqBlackBoxes.scala 104:19:@22943.4]
  mul_39_39_39_6_Unsigned_Use_Mults m ( // @[ZynqBlackBoxes.scala 104:19:@22943.4]
    .P(m_P),
    .B(m_B),
    .A(m_A),
    .CE(m_CE),
    .CLK(m_CLK)
  );
  assign io_out = m_P; // @[ZynqBlackBoxes.scala 109:12:@22953.4]
  assign m_B = io_b; // @[ZynqBlackBoxes.scala 107:12:@22951.4]
  assign m_A = io_a; // @[ZynqBlackBoxes.scala 106:12:@22950.4]
  assign m_CE = io_flow; // @[ZynqBlackBoxes.scala 108:13:@22952.4]
  assign m_CLK = clock; // @[ZynqBlackBoxes.scala 105:14:@22949.4]
endmodule
module fix2fixBox_118( // @[:@22955.2]
  input  [38:0] io_a, // @[:@22958.4]
  output [31:0] io_b // @[:@22958.4]
);
  wire [6:0] tmp_frac; // @[Converter.scala 38:42:@22966.4]
  wire [24:0] new_dec; // @[Converter.scala 88:34:@22969.4]
  assign tmp_frac = io_a[13:7]; // @[Converter.scala 38:42:@22966.4]
  assign new_dec = io_a[38:14]; // @[Converter.scala 88:34:@22969.4]
  assign io_b = {new_dec,tmp_frac}; // @[Converter.scala 94:38:@22972.4]
endmodule
module x375_mul( // @[:@22974.2]
  input         clock, // @[:@22975.4]
  input  [31:0] io_a, // @[:@22977.4]
  input         io_flow, // @[:@22977.4]
  output [31:0] io_result // @[:@22977.4]
);
  wire  x375_mul_clock; // @[BigIPZynq.scala 63:21:@22992.4]
  wire  x375_mul_io_flow; // @[BigIPZynq.scala 63:21:@22992.4]
  wire [38:0] x375_mul_io_a; // @[BigIPZynq.scala 63:21:@22992.4]
  wire [38:0] x375_mul_io_b; // @[BigIPZynq.scala 63:21:@22992.4]
  wire [38:0] x375_mul_io_out; // @[BigIPZynq.scala 63:21:@22992.4]
  wire [38:0] fix2fixBox_io_a; // @[Math.scala 253:30:@23000.4]
  wire [31:0] fix2fixBox_io_b; // @[Math.scala 253:30:@23000.4]
  wire  _T_16; // @[FixedPoint.scala 50:25:@22984.4]
  wire [6:0] _T_20; // @[Bitwise.scala 72:12:@22986.4]
  Multiplier_9 x375_mul ( // @[BigIPZynq.scala 63:21:@22992.4]
    .clock(x375_mul_clock),
    .io_flow(x375_mul_io_flow),
    .io_a(x375_mul_io_a),
    .io_b(x375_mul_io_b),
    .io_out(x375_mul_io_out)
  );
  fix2fixBox_118 fix2fixBox ( // @[Math.scala 253:30:@23000.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign _T_16 = io_a[31]; // @[FixedPoint.scala 50:25:@22984.4]
  assign _T_20 = _T_16 ? 7'h7f : 7'h0; // @[Bitwise.scala 72:12:@22986.4]
  assign io_result = fix2fixBox_io_b; // @[Math.scala 259:17:@23008.4]
  assign x375_mul_clock = clock; // @[:@22993.4]
  assign x375_mul_io_flow = io_flow; // @[BigIPZynq.scala 66:17:@22997.4]
  assign x375_mul_io_a = {_T_20,io_a}; // @[BigIPZynq.scala 64:14:@22995.4]
  assign x375_mul_io_b = 39'h8; // @[BigIPZynq.scala 65:14:@22996.4]
  assign fix2fixBox_io_a = x375_mul_io_out; // @[Math.scala 254:23:@23003.4]
endmodule
module fix2fixBox_119( // @[:@23010.2]
  input  [31:0] io_a, // @[:@23013.4]
  output [31:0] io_b // @[:@23013.4]
);
  wire [24:0] _T_25; // @[Converter.scala 84:75:@23025.4]
  assign _T_25 = io_a[31:7]; // @[Converter.scala 84:75:@23025.4]
  assign io_b = {7'h0,_T_25}; // @[Converter.scala 95:38:@23028.4]
endmodule
module x376( // @[:@23030.2]
  input  [31:0] io_b, // @[:@23033.4]
  output [31:0] io_result // @[:@23033.4]
);
  wire [31:0] fix2fixBox_io_a; // @[BigIPZynq.scala 219:30:@23038.4]
  wire [31:0] fix2fixBox_io_b; // @[BigIPZynq.scala 219:30:@23038.4]
  fix2fixBox_119 fix2fixBox ( // @[BigIPZynq.scala 219:30:@23038.4]
    .io_a(fix2fixBox_io_a),
    .io_b(fix2fixBox_io_b)
  );
  assign io_result = fix2fixBox_io_b; // @[Math.scala 717:17:@23046.4]
  assign fix2fixBox_io_a = io_b; // @[BigIPZynq.scala 220:23:@23041.4]
endmodule
module RetimeWrapper_262( // @[:@25266.2]
  input         clock, // @[:@25267.4]
  input         reset, // @[:@25268.4]
  input         io_flow, // @[:@25269.4]
  input  [63:0] io_in, // @[:@25269.4]
  output [63:0] io_out // @[:@25269.4]
);
  wire [63:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@25271.4]
  wire [63:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@25271.4]
  wire [63:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@25271.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@25271.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@25271.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@25271.4]
  RetimeShiftRegister #(.WIDTH(64), .STAGES(3)) sr ( // @[RetimeShiftRegister.scala 15:20:@25271.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@25284.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@25283.4]
  assign sr_init = 64'h0; // @[RetimeShiftRegister.scala 19:16:@25282.4]
  assign sr_flow = io_flow; // @[RetimeShiftRegister.scala 18:16:@25281.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@25280.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@25278.4]
endmodule
module x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1( // @[:@25382.2]
  input          clock, // @[:@25383.4]
  input          reset, // @[:@25384.4]
  output         io_in_x221_TREADY, // @[:@25385.4]
  input  [255:0] io_in_x221_TDATA, // @[:@25385.4]
  input  [7:0]   io_in_x221_TID, // @[:@25385.4]
  input  [7:0]   io_in_x221_TDEST, // @[:@25385.4]
  output         io_in_x222_TVALID, // @[:@25385.4]
  input          io_in_x222_TREADY, // @[:@25385.4]
  output [255:0] io_in_x222_TDATA, // @[:@25385.4]
  input          io_sigsIn_backpressure, // @[:@25385.4]
  input          io_sigsIn_datapathEn, // @[:@25385.4]
  input          io_sigsIn_break, // @[:@25385.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_1, // @[:@25385.4]
  input  [31:0]  io_sigsIn_cchainOutputs_0_counts_0, // @[:@25385.4]
  input          io_sigsIn_cchainOutputs_0_oobs_0, // @[:@25385.4]
  input          io_sigsIn_cchainOutputs_0_oobs_1, // @[:@25385.4]
  input          io_rr // @[:@25385.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@25399.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@25399.4]
  wire [31:0] __1_io_b; // @[Math.scala 720:24:@25411.4]
  wire [31:0] __1_io_result; // @[Math.scala 720:24:@25411.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@25434.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@25434.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@25434.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@25434.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@25434.4]
  wire  x258_lb_0_clock; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_reset; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_11_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_11_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_11_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_11_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_11_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_11_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_10_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_10_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_10_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_10_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_10_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_10_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_9_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_9_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_9_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_9_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_9_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_9_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_8_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_8_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_8_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_8_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_8_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_8_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_7_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_7_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_7_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_7_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_7_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_7_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_6_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_6_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_6_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_6_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_6_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_6_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_5_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_5_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_5_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_5_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_5_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_5_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_4_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_4_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_4_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_4_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_4_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_4_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_3_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_3_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_3_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_3_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_3_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_3_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_2_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_2_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_2_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_2_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_2_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_2_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_1_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_1_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_1_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_1_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_1_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_1_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_0_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_rPort_0_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_rPort_0_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_0_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_rPort_0_backpressure; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_rPort_0_output_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_wPort_1_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_wPort_1_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_wPort_1_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_wPort_1_data_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_wPort_1_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_wPort_0_banks_1; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [2:0] x258_lb_0_io_wPort_0_banks_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [8:0] x258_lb_0_io_wPort_0_ofs_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire [31:0] x258_lb_0_io_wPort_0_data_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x258_lb_0_io_wPort_0_en_0; // @[m_x258_lb_0.scala 39:17:@25444.4]
  wire  x464_sub_1_clock; // @[Math.scala 191:24:@25607.4]
  wire  x464_sub_1_reset; // @[Math.scala 191:24:@25607.4]
  wire [31:0] x464_sub_1_io_a; // @[Math.scala 191:24:@25607.4]
  wire [31:0] x464_sub_1_io_b; // @[Math.scala 191:24:@25607.4]
  wire  x464_sub_1_io_flow; // @[Math.scala 191:24:@25607.4]
  wire [31:0] x464_sub_1_io_result; // @[Math.scala 191:24:@25607.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@25634.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@25634.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@25634.4]
  wire [31:0] RetimeWrapper_1_io_in; // @[package.scala 93:22:@25634.4]
  wire [31:0] RetimeWrapper_1_io_out; // @[package.scala 93:22:@25634.4]
  wire  x267_sum_1_clock; // @[Math.scala 150:24:@25643.4]
  wire  x267_sum_1_reset; // @[Math.scala 150:24:@25643.4]
  wire [31:0] x267_sum_1_io_a; // @[Math.scala 150:24:@25643.4]
  wire [31:0] x267_sum_1_io_b; // @[Math.scala 150:24:@25643.4]
  wire  x267_sum_1_io_flow; // @[Math.scala 150:24:@25643.4]
  wire [31:0] x267_sum_1_io_result; // @[Math.scala 150:24:@25643.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@25653.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@25653.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@25653.4]
  wire [31:0] RetimeWrapper_2_io_in; // @[package.scala 93:22:@25653.4]
  wire [31:0] RetimeWrapper_2_io_out; // @[package.scala 93:22:@25653.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@25662.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@25662.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@25662.4]
  wire [31:0] RetimeWrapper_3_io_in; // @[package.scala 93:22:@25662.4]
  wire [31:0] RetimeWrapper_3_io_out; // @[package.scala 93:22:@25662.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@25671.4]
  wire [31:0] RetimeWrapper_4_io_in; // @[package.scala 93:22:@25671.4]
  wire [31:0] RetimeWrapper_4_io_out; // @[package.scala 93:22:@25671.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@25680.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@25680.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@25680.4]
  wire [31:0] RetimeWrapper_5_io_in; // @[package.scala 93:22:@25680.4]
  wire [31:0] RetimeWrapper_5_io_out; // @[package.scala 93:22:@25680.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@25689.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@25689.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@25689.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@25689.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@25689.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@25698.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@25709.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@25709.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@25709.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@25709.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@25709.4]
  wire  x269_rdcol_1_clock; // @[Math.scala 150:24:@25732.4]
  wire  x269_rdcol_1_reset; // @[Math.scala 150:24:@25732.4]
  wire [31:0] x269_rdcol_1_io_a; // @[Math.scala 150:24:@25732.4]
  wire [31:0] x269_rdcol_1_io_b; // @[Math.scala 150:24:@25732.4]
  wire  x269_rdcol_1_io_flow; // @[Math.scala 150:24:@25732.4]
  wire [31:0] x269_rdcol_1_io_result; // @[Math.scala 150:24:@25732.4]
  wire  x273_sum_1_clock; // @[Math.scala 150:24:@25772.4]
  wire  x273_sum_1_reset; // @[Math.scala 150:24:@25772.4]
  wire [31:0] x273_sum_1_io_a; // @[Math.scala 150:24:@25772.4]
  wire [31:0] x273_sum_1_io_b; // @[Math.scala 150:24:@25772.4]
  wire  x273_sum_1_io_flow; // @[Math.scala 150:24:@25772.4]
  wire [31:0] x273_sum_1_io_result; // @[Math.scala 150:24:@25772.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@25782.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@25782.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@25782.4]
  wire [31:0] RetimeWrapper_9_io_in; // @[package.scala 93:22:@25782.4]
  wire [31:0] RetimeWrapper_9_io_out; // @[package.scala 93:22:@25782.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@25791.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@25791.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@25791.4]
  wire [31:0] RetimeWrapper_10_io_in; // @[package.scala 93:22:@25791.4]
  wire [31:0] RetimeWrapper_10_io_out; // @[package.scala 93:22:@25791.4]
  wire  RetimeWrapper_11_clock; // @[package.scala 93:22:@25800.4]
  wire  RetimeWrapper_11_reset; // @[package.scala 93:22:@25800.4]
  wire  RetimeWrapper_11_io_flow; // @[package.scala 93:22:@25800.4]
  wire [31:0] RetimeWrapper_11_io_in; // @[package.scala 93:22:@25800.4]
  wire [31:0] RetimeWrapper_11_io_out; // @[package.scala 93:22:@25800.4]
  wire  RetimeWrapper_12_clock; // @[package.scala 93:22:@25811.4]
  wire  RetimeWrapper_12_reset; // @[package.scala 93:22:@25811.4]
  wire  RetimeWrapper_12_io_flow; // @[package.scala 93:22:@25811.4]
  wire  RetimeWrapper_12_io_in; // @[package.scala 93:22:@25811.4]
  wire  RetimeWrapper_12_io_out; // @[package.scala 93:22:@25811.4]
  wire  RetimeWrapper_13_clock; // @[package.scala 93:22:@25832.4]
  wire  RetimeWrapper_13_reset; // @[package.scala 93:22:@25832.4]
  wire  RetimeWrapper_13_io_flow; // @[package.scala 93:22:@25832.4]
  wire [31:0] RetimeWrapper_13_io_in; // @[package.scala 93:22:@25832.4]
  wire [31:0] RetimeWrapper_13_io_out; // @[package.scala 93:22:@25832.4]
  wire  RetimeWrapper_14_clock; // @[package.scala 93:22:@25848.4]
  wire  RetimeWrapper_14_reset; // @[package.scala 93:22:@25848.4]
  wire  RetimeWrapper_14_io_flow; // @[package.scala 93:22:@25848.4]
  wire [31:0] RetimeWrapper_14_io_in; // @[package.scala 93:22:@25848.4]
  wire [31:0] RetimeWrapper_14_io_out; // @[package.scala 93:22:@25848.4]
  wire  RetimeWrapper_15_clock; // @[package.scala 93:22:@25864.4]
  wire  RetimeWrapper_15_reset; // @[package.scala 93:22:@25864.4]
  wire  RetimeWrapper_15_io_flow; // @[package.scala 93:22:@25864.4]
  wire  RetimeWrapper_15_io_in; // @[package.scala 93:22:@25864.4]
  wire  RetimeWrapper_15_io_out; // @[package.scala 93:22:@25864.4]
  wire  RetimeWrapper_16_clock; // @[package.scala 93:22:@25879.4]
  wire  RetimeWrapper_16_reset; // @[package.scala 93:22:@25879.4]
  wire  RetimeWrapper_16_io_flow; // @[package.scala 93:22:@25879.4]
  wire [31:0] RetimeWrapper_16_io_in; // @[package.scala 93:22:@25879.4]
  wire [31:0] RetimeWrapper_16_io_out; // @[package.scala 93:22:@25879.4]
  wire  RetimeWrapper_17_clock; // @[package.scala 93:22:@25888.4]
  wire  RetimeWrapper_17_reset; // @[package.scala 93:22:@25888.4]
  wire  RetimeWrapper_17_io_flow; // @[package.scala 93:22:@25888.4]
  wire  RetimeWrapper_17_io_in; // @[package.scala 93:22:@25888.4]
  wire  RetimeWrapper_17_io_out; // @[package.scala 93:22:@25888.4]
  wire  RetimeWrapper_18_clock; // @[package.scala 93:22:@25897.4]
  wire  RetimeWrapper_18_reset; // @[package.scala 93:22:@25897.4]
  wire  RetimeWrapper_18_io_flow; // @[package.scala 93:22:@25897.4]
  wire  RetimeWrapper_18_io_in; // @[package.scala 93:22:@25897.4]
  wire  RetimeWrapper_18_io_out; // @[package.scala 93:22:@25897.4]
  wire  RetimeWrapper_19_clock; // @[package.scala 93:22:@25906.4]
  wire  RetimeWrapper_19_reset; // @[package.scala 93:22:@25906.4]
  wire  RetimeWrapper_19_io_flow; // @[package.scala 93:22:@25906.4]
  wire [31:0] RetimeWrapper_19_io_in; // @[package.scala 93:22:@25906.4]
  wire [31:0] RetimeWrapper_19_io_out; // @[package.scala 93:22:@25906.4]
  wire  RetimeWrapper_20_clock; // @[package.scala 93:22:@25915.4]
  wire  RetimeWrapper_20_reset; // @[package.scala 93:22:@25915.4]
  wire  RetimeWrapper_20_io_flow; // @[package.scala 93:22:@25915.4]
  wire [31:0] RetimeWrapper_20_io_in; // @[package.scala 93:22:@25915.4]
  wire [31:0] RetimeWrapper_20_io_out; // @[package.scala 93:22:@25915.4]
  wire  RetimeWrapper_21_clock; // @[package.scala 93:22:@25924.4]
  wire  RetimeWrapper_21_reset; // @[package.scala 93:22:@25924.4]
  wire  RetimeWrapper_21_io_flow; // @[package.scala 93:22:@25924.4]
  wire  RetimeWrapper_21_io_in; // @[package.scala 93:22:@25924.4]
  wire  RetimeWrapper_21_io_out; // @[package.scala 93:22:@25924.4]
  wire  RetimeWrapper_22_clock; // @[package.scala 93:22:@25936.4]
  wire  RetimeWrapper_22_reset; // @[package.scala 93:22:@25936.4]
  wire  RetimeWrapper_22_io_flow; // @[package.scala 93:22:@25936.4]
  wire  RetimeWrapper_22_io_in; // @[package.scala 93:22:@25936.4]
  wire  RetimeWrapper_22_io_out; // @[package.scala 93:22:@25936.4]
  wire  RetimeWrapper_23_clock; // @[package.scala 93:22:@25957.4]
  wire  RetimeWrapper_23_reset; // @[package.scala 93:22:@25957.4]
  wire  RetimeWrapper_23_io_flow; // @[package.scala 93:22:@25957.4]
  wire [31:0] RetimeWrapper_23_io_in; // @[package.scala 93:22:@25957.4]
  wire [31:0] RetimeWrapper_23_io_out; // @[package.scala 93:22:@25957.4]
  wire  RetimeWrapper_24_clock; // @[package.scala 93:22:@25981.4]
  wire  RetimeWrapper_24_reset; // @[package.scala 93:22:@25981.4]
  wire  RetimeWrapper_24_io_flow; // @[package.scala 93:22:@25981.4]
  wire  RetimeWrapper_24_io_in; // @[package.scala 93:22:@25981.4]
  wire  RetimeWrapper_24_io_out; // @[package.scala 93:22:@25981.4]
  wire  RetimeWrapper_25_clock; // @[package.scala 93:22:@25990.4]
  wire  RetimeWrapper_25_reset; // @[package.scala 93:22:@25990.4]
  wire  RetimeWrapper_25_io_flow; // @[package.scala 93:22:@25990.4]
  wire [31:0] RetimeWrapper_25_io_in; // @[package.scala 93:22:@25990.4]
  wire [31:0] RetimeWrapper_25_io_out; // @[package.scala 93:22:@25990.4]
  wire  RetimeWrapper_26_clock; // @[package.scala 93:22:@25999.4]
  wire  RetimeWrapper_26_reset; // @[package.scala 93:22:@25999.4]
  wire  RetimeWrapper_26_io_flow; // @[package.scala 93:22:@25999.4]
  wire [31:0] RetimeWrapper_26_io_in; // @[package.scala 93:22:@25999.4]
  wire [31:0] RetimeWrapper_26_io_out; // @[package.scala 93:22:@25999.4]
  wire  RetimeWrapper_27_clock; // @[package.scala 93:22:@26011.4]
  wire  RetimeWrapper_27_reset; // @[package.scala 93:22:@26011.4]
  wire  RetimeWrapper_27_io_flow; // @[package.scala 93:22:@26011.4]
  wire  RetimeWrapper_27_io_in; // @[package.scala 93:22:@26011.4]
  wire  RetimeWrapper_27_io_out; // @[package.scala 93:22:@26011.4]
  wire  x287_rdcol_1_clock; // @[Math.scala 150:24:@26034.4]
  wire  x287_rdcol_1_reset; // @[Math.scala 150:24:@26034.4]
  wire [31:0] x287_rdcol_1_io_a; // @[Math.scala 150:24:@26034.4]
  wire [31:0] x287_rdcol_1_io_b; // @[Math.scala 150:24:@26034.4]
  wire  x287_rdcol_1_io_flow; // @[Math.scala 150:24:@26034.4]
  wire [31:0] x287_rdcol_1_io_result; // @[Math.scala 150:24:@26034.4]
  wire  RetimeWrapper_28_clock; // @[package.scala 93:22:@26085.4]
  wire  RetimeWrapper_28_reset; // @[package.scala 93:22:@26085.4]
  wire  RetimeWrapper_28_io_flow; // @[package.scala 93:22:@26085.4]
  wire [31:0] RetimeWrapper_28_io_in; // @[package.scala 93:22:@26085.4]
  wire [31:0] RetimeWrapper_28_io_out; // @[package.scala 93:22:@26085.4]
  wire  x293_sum_1_clock; // @[Math.scala 150:24:@26094.4]
  wire  x293_sum_1_reset; // @[Math.scala 150:24:@26094.4]
  wire [31:0] x293_sum_1_io_a; // @[Math.scala 150:24:@26094.4]
  wire [31:0] x293_sum_1_io_b; // @[Math.scala 150:24:@26094.4]
  wire  x293_sum_1_io_flow; // @[Math.scala 150:24:@26094.4]
  wire [31:0] x293_sum_1_io_result; // @[Math.scala 150:24:@26094.4]
  wire  RetimeWrapper_29_clock; // @[package.scala 93:22:@26104.4]
  wire  RetimeWrapper_29_reset; // @[package.scala 93:22:@26104.4]
  wire  RetimeWrapper_29_io_flow; // @[package.scala 93:22:@26104.4]
  wire [31:0] RetimeWrapper_29_io_in; // @[package.scala 93:22:@26104.4]
  wire [31:0] RetimeWrapper_29_io_out; // @[package.scala 93:22:@26104.4]
  wire  RetimeWrapper_30_clock; // @[package.scala 93:22:@26113.4]
  wire  RetimeWrapper_30_reset; // @[package.scala 93:22:@26113.4]
  wire  RetimeWrapper_30_io_flow; // @[package.scala 93:22:@26113.4]
  wire [31:0] RetimeWrapper_30_io_in; // @[package.scala 93:22:@26113.4]
  wire [31:0] RetimeWrapper_30_io_out; // @[package.scala 93:22:@26113.4]
  wire  RetimeWrapper_31_clock; // @[package.scala 93:22:@26122.4]
  wire  RetimeWrapper_31_reset; // @[package.scala 93:22:@26122.4]
  wire  RetimeWrapper_31_io_flow; // @[package.scala 93:22:@26122.4]
  wire  RetimeWrapper_31_io_in; // @[package.scala 93:22:@26122.4]
  wire  RetimeWrapper_31_io_out; // @[package.scala 93:22:@26122.4]
  wire  RetimeWrapper_32_clock; // @[package.scala 93:22:@26134.4]
  wire  RetimeWrapper_32_reset; // @[package.scala 93:22:@26134.4]
  wire  RetimeWrapper_32_io_flow; // @[package.scala 93:22:@26134.4]
  wire  RetimeWrapper_32_io_in; // @[package.scala 93:22:@26134.4]
  wire  RetimeWrapper_32_io_out; // @[package.scala 93:22:@26134.4]
  wire  x296_rdcol_1_clock; // @[Math.scala 150:24:@26157.4]
  wire  x296_rdcol_1_reset; // @[Math.scala 150:24:@26157.4]
  wire [31:0] x296_rdcol_1_io_a; // @[Math.scala 150:24:@26157.4]
  wire [31:0] x296_rdcol_1_io_b; // @[Math.scala 150:24:@26157.4]
  wire  x296_rdcol_1_io_flow; // @[Math.scala 150:24:@26157.4]
  wire [31:0] x296_rdcol_1_io_result; // @[Math.scala 150:24:@26157.4]
  wire  x302_sum_1_clock; // @[Math.scala 150:24:@26208.4]
  wire  x302_sum_1_reset; // @[Math.scala 150:24:@26208.4]
  wire [31:0] x302_sum_1_io_a; // @[Math.scala 150:24:@26208.4]
  wire [31:0] x302_sum_1_io_b; // @[Math.scala 150:24:@26208.4]
  wire  x302_sum_1_io_flow; // @[Math.scala 150:24:@26208.4]
  wire [31:0] x302_sum_1_io_result; // @[Math.scala 150:24:@26208.4]
  wire  RetimeWrapper_33_clock; // @[package.scala 93:22:@26218.4]
  wire  RetimeWrapper_33_reset; // @[package.scala 93:22:@26218.4]
  wire  RetimeWrapper_33_io_flow; // @[package.scala 93:22:@26218.4]
  wire [31:0] RetimeWrapper_33_io_in; // @[package.scala 93:22:@26218.4]
  wire [31:0] RetimeWrapper_33_io_out; // @[package.scala 93:22:@26218.4]
  wire  RetimeWrapper_34_clock; // @[package.scala 93:22:@26227.4]
  wire  RetimeWrapper_34_reset; // @[package.scala 93:22:@26227.4]
  wire  RetimeWrapper_34_io_flow; // @[package.scala 93:22:@26227.4]
  wire [31:0] RetimeWrapper_34_io_in; // @[package.scala 93:22:@26227.4]
  wire [31:0] RetimeWrapper_34_io_out; // @[package.scala 93:22:@26227.4]
  wire  RetimeWrapper_35_clock; // @[package.scala 93:22:@26236.4]
  wire  RetimeWrapper_35_reset; // @[package.scala 93:22:@26236.4]
  wire  RetimeWrapper_35_io_flow; // @[package.scala 93:22:@26236.4]
  wire  RetimeWrapper_35_io_in; // @[package.scala 93:22:@26236.4]
  wire  RetimeWrapper_35_io_out; // @[package.scala 93:22:@26236.4]
  wire  RetimeWrapper_36_clock; // @[package.scala 93:22:@26248.4]
  wire  RetimeWrapper_36_reset; // @[package.scala 93:22:@26248.4]
  wire  RetimeWrapper_36_io_flow; // @[package.scala 93:22:@26248.4]
  wire  RetimeWrapper_36_io_in; // @[package.scala 93:22:@26248.4]
  wire  RetimeWrapper_36_io_out; // @[package.scala 93:22:@26248.4]
  wire  x305_rdrow_1_clock; // @[Math.scala 191:24:@26271.4]
  wire  x305_rdrow_1_reset; // @[Math.scala 191:24:@26271.4]
  wire [31:0] x305_rdrow_1_io_a; // @[Math.scala 191:24:@26271.4]
  wire [31:0] x305_rdrow_1_io_b; // @[Math.scala 191:24:@26271.4]
  wire  x305_rdrow_1_io_flow; // @[Math.scala 191:24:@26271.4]
  wire [31:0] x305_rdrow_1_io_result; // @[Math.scala 191:24:@26271.4]
  wire  x472_sub_1_clock; // @[Math.scala 191:24:@26343.4]
  wire  x472_sub_1_reset; // @[Math.scala 191:24:@26343.4]
  wire [31:0] x472_sub_1_io_a; // @[Math.scala 191:24:@26343.4]
  wire [31:0] x472_sub_1_io_b; // @[Math.scala 191:24:@26343.4]
  wire  x472_sub_1_io_flow; // @[Math.scala 191:24:@26343.4]
  wire [31:0] x472_sub_1_io_result; // @[Math.scala 191:24:@26343.4]
  wire  RetimeWrapper_37_clock; // @[package.scala 93:22:@26353.4]
  wire  RetimeWrapper_37_reset; // @[package.scala 93:22:@26353.4]
  wire  RetimeWrapper_37_io_flow; // @[package.scala 93:22:@26353.4]
  wire [31:0] RetimeWrapper_37_io_in; // @[package.scala 93:22:@26353.4]
  wire [31:0] RetimeWrapper_37_io_out; // @[package.scala 93:22:@26353.4]
  wire  x313_sum_1_clock; // @[Math.scala 150:24:@26362.4]
  wire  x313_sum_1_reset; // @[Math.scala 150:24:@26362.4]
  wire [31:0] x313_sum_1_io_a; // @[Math.scala 150:24:@26362.4]
  wire [31:0] x313_sum_1_io_b; // @[Math.scala 150:24:@26362.4]
  wire  x313_sum_1_io_flow; // @[Math.scala 150:24:@26362.4]
  wire [31:0] x313_sum_1_io_result; // @[Math.scala 150:24:@26362.4]
  wire  RetimeWrapper_38_clock; // @[package.scala 93:22:@26372.4]
  wire  RetimeWrapper_38_reset; // @[package.scala 93:22:@26372.4]
  wire  RetimeWrapper_38_io_flow; // @[package.scala 93:22:@26372.4]
  wire [31:0] RetimeWrapper_38_io_in; // @[package.scala 93:22:@26372.4]
  wire [31:0] RetimeWrapper_38_io_out; // @[package.scala 93:22:@26372.4]
  wire  RetimeWrapper_39_clock; // @[package.scala 93:22:@26381.4]
  wire  RetimeWrapper_39_reset; // @[package.scala 93:22:@26381.4]
  wire  RetimeWrapper_39_io_flow; // @[package.scala 93:22:@26381.4]
  wire  RetimeWrapper_39_io_in; // @[package.scala 93:22:@26381.4]
  wire  RetimeWrapper_39_io_out; // @[package.scala 93:22:@26381.4]
  wire  RetimeWrapper_40_clock; // @[package.scala 93:22:@26393.4]
  wire  RetimeWrapper_40_reset; // @[package.scala 93:22:@26393.4]
  wire  RetimeWrapper_40_io_flow; // @[package.scala 93:22:@26393.4]
  wire  RetimeWrapper_40_io_in; // @[package.scala 93:22:@26393.4]
  wire  RetimeWrapper_40_io_out; // @[package.scala 93:22:@26393.4]
  wire  RetimeWrapper_41_clock; // @[package.scala 93:22:@26414.4]
  wire  RetimeWrapper_41_reset; // @[package.scala 93:22:@26414.4]
  wire  RetimeWrapper_41_io_flow; // @[package.scala 93:22:@26414.4]
  wire  RetimeWrapper_41_io_in; // @[package.scala 93:22:@26414.4]
  wire  RetimeWrapper_41_io_out; // @[package.scala 93:22:@26414.4]
  wire  RetimeWrapper_42_clock; // @[package.scala 93:22:@26429.4]
  wire  RetimeWrapper_42_reset; // @[package.scala 93:22:@26429.4]
  wire  RetimeWrapper_42_io_flow; // @[package.scala 93:22:@26429.4]
  wire [31:0] RetimeWrapper_42_io_in; // @[package.scala 93:22:@26429.4]
  wire [31:0] RetimeWrapper_42_io_out; // @[package.scala 93:22:@26429.4]
  wire  x318_sum_1_clock; // @[Math.scala 150:24:@26440.4]
  wire  x318_sum_1_reset; // @[Math.scala 150:24:@26440.4]
  wire [31:0] x318_sum_1_io_a; // @[Math.scala 150:24:@26440.4]
  wire [31:0] x318_sum_1_io_b; // @[Math.scala 150:24:@26440.4]
  wire  x318_sum_1_io_flow; // @[Math.scala 150:24:@26440.4]
  wire [31:0] x318_sum_1_io_result; // @[Math.scala 150:24:@26440.4]
  wire  RetimeWrapper_43_clock; // @[package.scala 93:22:@26450.4]
  wire  RetimeWrapper_43_reset; // @[package.scala 93:22:@26450.4]
  wire  RetimeWrapper_43_io_flow; // @[package.scala 93:22:@26450.4]
  wire  RetimeWrapper_43_io_in; // @[package.scala 93:22:@26450.4]
  wire  RetimeWrapper_43_io_out; // @[package.scala 93:22:@26450.4]
  wire  RetimeWrapper_44_clock; // @[package.scala 93:22:@26462.4]
  wire  RetimeWrapper_44_reset; // @[package.scala 93:22:@26462.4]
  wire  RetimeWrapper_44_io_flow; // @[package.scala 93:22:@26462.4]
  wire  RetimeWrapper_44_io_in; // @[package.scala 93:22:@26462.4]
  wire  RetimeWrapper_44_io_out; // @[package.scala 93:22:@26462.4]
  wire  RetimeWrapper_45_clock; // @[package.scala 93:22:@26489.4]
  wire  RetimeWrapper_45_reset; // @[package.scala 93:22:@26489.4]
  wire  RetimeWrapper_45_io_flow; // @[package.scala 93:22:@26489.4]
  wire [31:0] RetimeWrapper_45_io_in; // @[package.scala 93:22:@26489.4]
  wire [31:0] RetimeWrapper_45_io_out; // @[package.scala 93:22:@26489.4]
  wire  x323_sum_1_clock; // @[Math.scala 150:24:@26498.4]
  wire  x323_sum_1_reset; // @[Math.scala 150:24:@26498.4]
  wire [31:0] x323_sum_1_io_a; // @[Math.scala 150:24:@26498.4]
  wire [31:0] x323_sum_1_io_b; // @[Math.scala 150:24:@26498.4]
  wire  x323_sum_1_io_flow; // @[Math.scala 150:24:@26498.4]
  wire [31:0] x323_sum_1_io_result; // @[Math.scala 150:24:@26498.4]
  wire  RetimeWrapper_46_clock; // @[package.scala 93:22:@26508.4]
  wire  RetimeWrapper_46_reset; // @[package.scala 93:22:@26508.4]
  wire  RetimeWrapper_46_io_flow; // @[package.scala 93:22:@26508.4]
  wire  RetimeWrapper_46_io_in; // @[package.scala 93:22:@26508.4]
  wire  RetimeWrapper_46_io_out; // @[package.scala 93:22:@26508.4]
  wire  RetimeWrapper_47_clock; // @[package.scala 93:22:@26520.4]
  wire  RetimeWrapper_47_reset; // @[package.scala 93:22:@26520.4]
  wire  RetimeWrapper_47_io_flow; // @[package.scala 93:22:@26520.4]
  wire  RetimeWrapper_47_io_in; // @[package.scala 93:22:@26520.4]
  wire  RetimeWrapper_47_io_out; // @[package.scala 93:22:@26520.4]
  wire  RetimeWrapper_48_clock; // @[package.scala 93:22:@26547.4]
  wire  RetimeWrapper_48_reset; // @[package.scala 93:22:@26547.4]
  wire  RetimeWrapper_48_io_flow; // @[package.scala 93:22:@26547.4]
  wire [31:0] RetimeWrapper_48_io_in; // @[package.scala 93:22:@26547.4]
  wire [31:0] RetimeWrapper_48_io_out; // @[package.scala 93:22:@26547.4]
  wire  x328_sum_1_clock; // @[Math.scala 150:24:@26556.4]
  wire  x328_sum_1_reset; // @[Math.scala 150:24:@26556.4]
  wire [31:0] x328_sum_1_io_a; // @[Math.scala 150:24:@26556.4]
  wire [31:0] x328_sum_1_io_b; // @[Math.scala 150:24:@26556.4]
  wire  x328_sum_1_io_flow; // @[Math.scala 150:24:@26556.4]
  wire [31:0] x328_sum_1_io_result; // @[Math.scala 150:24:@26556.4]
  wire  RetimeWrapper_49_clock; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_49_reset; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_49_io_flow; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_49_io_in; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_49_io_out; // @[package.scala 93:22:@26566.4]
  wire  RetimeWrapper_50_clock; // @[package.scala 93:22:@26578.4]
  wire  RetimeWrapper_50_reset; // @[package.scala 93:22:@26578.4]
  wire  RetimeWrapper_50_io_flow; // @[package.scala 93:22:@26578.4]
  wire  RetimeWrapper_50_io_in; // @[package.scala 93:22:@26578.4]
  wire  RetimeWrapper_50_io_out; // @[package.scala 93:22:@26578.4]
  wire  x331_rdrow_1_clock; // @[Math.scala 191:24:@26601.4]
  wire  x331_rdrow_1_reset; // @[Math.scala 191:24:@26601.4]
  wire [31:0] x331_rdrow_1_io_a; // @[Math.scala 191:24:@26601.4]
  wire [31:0] x331_rdrow_1_io_b; // @[Math.scala 191:24:@26601.4]
  wire  x331_rdrow_1_io_flow; // @[Math.scala 191:24:@26601.4]
  wire [31:0] x331_rdrow_1_io_result; // @[Math.scala 191:24:@26601.4]
  wire  x477_sub_1_clock; // @[Math.scala 191:24:@26673.4]
  wire  x477_sub_1_reset; // @[Math.scala 191:24:@26673.4]
  wire [31:0] x477_sub_1_io_a; // @[Math.scala 191:24:@26673.4]
  wire [31:0] x477_sub_1_io_b; // @[Math.scala 191:24:@26673.4]
  wire  x477_sub_1_io_flow; // @[Math.scala 191:24:@26673.4]
  wire [31:0] x477_sub_1_io_result; // @[Math.scala 191:24:@26673.4]
  wire  x339_sum_1_clock; // @[Math.scala 150:24:@26683.4]
  wire  x339_sum_1_reset; // @[Math.scala 150:24:@26683.4]
  wire [31:0] x339_sum_1_io_a; // @[Math.scala 150:24:@26683.4]
  wire [31:0] x339_sum_1_io_b; // @[Math.scala 150:24:@26683.4]
  wire  x339_sum_1_io_flow; // @[Math.scala 150:24:@26683.4]
  wire [31:0] x339_sum_1_io_result; // @[Math.scala 150:24:@26683.4]
  wire  RetimeWrapper_51_clock; // @[package.scala 93:22:@26693.4]
  wire  RetimeWrapper_51_reset; // @[package.scala 93:22:@26693.4]
  wire  RetimeWrapper_51_io_flow; // @[package.scala 93:22:@26693.4]
  wire  RetimeWrapper_51_io_in; // @[package.scala 93:22:@26693.4]
  wire  RetimeWrapper_51_io_out; // @[package.scala 93:22:@26693.4]
  wire  RetimeWrapper_52_clock; // @[package.scala 93:22:@26702.4]
  wire  RetimeWrapper_52_reset; // @[package.scala 93:22:@26702.4]
  wire  RetimeWrapper_52_io_flow; // @[package.scala 93:22:@26702.4]
  wire [31:0] RetimeWrapper_52_io_in; // @[package.scala 93:22:@26702.4]
  wire [31:0] RetimeWrapper_52_io_out; // @[package.scala 93:22:@26702.4]
  wire  RetimeWrapper_53_clock; // @[package.scala 93:22:@26714.4]
  wire  RetimeWrapper_53_reset; // @[package.scala 93:22:@26714.4]
  wire  RetimeWrapper_53_io_flow; // @[package.scala 93:22:@26714.4]
  wire  RetimeWrapper_53_io_in; // @[package.scala 93:22:@26714.4]
  wire  RetimeWrapper_53_io_out; // @[package.scala 93:22:@26714.4]
  wire  x344_sum_1_clock; // @[Math.scala 150:24:@26741.4]
  wire  x344_sum_1_reset; // @[Math.scala 150:24:@26741.4]
  wire [31:0] x344_sum_1_io_a; // @[Math.scala 150:24:@26741.4]
  wire [31:0] x344_sum_1_io_b; // @[Math.scala 150:24:@26741.4]
  wire  x344_sum_1_io_flow; // @[Math.scala 150:24:@26741.4]
  wire [31:0] x344_sum_1_io_result; // @[Math.scala 150:24:@26741.4]
  wire  RetimeWrapper_54_clock; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_54_reset; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_54_io_flow; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_54_io_in; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_54_io_out; // @[package.scala 93:22:@26751.4]
  wire  RetimeWrapper_55_clock; // @[package.scala 93:22:@26763.4]
  wire  RetimeWrapper_55_reset; // @[package.scala 93:22:@26763.4]
  wire  RetimeWrapper_55_io_flow; // @[package.scala 93:22:@26763.4]
  wire  RetimeWrapper_55_io_in; // @[package.scala 93:22:@26763.4]
  wire  RetimeWrapper_55_io_out; // @[package.scala 93:22:@26763.4]
  wire  x349_sum_1_clock; // @[Math.scala 150:24:@26790.4]
  wire  x349_sum_1_reset; // @[Math.scala 150:24:@26790.4]
  wire [31:0] x349_sum_1_io_a; // @[Math.scala 150:24:@26790.4]
  wire [31:0] x349_sum_1_io_b; // @[Math.scala 150:24:@26790.4]
  wire  x349_sum_1_io_flow; // @[Math.scala 150:24:@26790.4]
  wire [31:0] x349_sum_1_io_result; // @[Math.scala 150:24:@26790.4]
  wire  RetimeWrapper_56_clock; // @[package.scala 93:22:@26800.4]
  wire  RetimeWrapper_56_reset; // @[package.scala 93:22:@26800.4]
  wire  RetimeWrapper_56_io_flow; // @[package.scala 93:22:@26800.4]
  wire  RetimeWrapper_56_io_in; // @[package.scala 93:22:@26800.4]
  wire  RetimeWrapper_56_io_out; // @[package.scala 93:22:@26800.4]
  wire  RetimeWrapper_57_clock; // @[package.scala 93:22:@26812.4]
  wire  RetimeWrapper_57_reset; // @[package.scala 93:22:@26812.4]
  wire  RetimeWrapper_57_io_flow; // @[package.scala 93:22:@26812.4]
  wire  RetimeWrapper_57_io_in; // @[package.scala 93:22:@26812.4]
  wire  RetimeWrapper_57_io_out; // @[package.scala 93:22:@26812.4]
  wire  x354_sum_1_clock; // @[Math.scala 150:24:@26841.4]
  wire  x354_sum_1_reset; // @[Math.scala 150:24:@26841.4]
  wire [31:0] x354_sum_1_io_a; // @[Math.scala 150:24:@26841.4]
  wire [31:0] x354_sum_1_io_b; // @[Math.scala 150:24:@26841.4]
  wire  x354_sum_1_io_flow; // @[Math.scala 150:24:@26841.4]
  wire [31:0] x354_sum_1_io_result; // @[Math.scala 150:24:@26841.4]
  wire  RetimeWrapper_58_clock; // @[package.scala 93:22:@26851.4]
  wire  RetimeWrapper_58_reset; // @[package.scala 93:22:@26851.4]
  wire  RetimeWrapper_58_io_flow; // @[package.scala 93:22:@26851.4]
  wire  RetimeWrapper_58_io_in; // @[package.scala 93:22:@26851.4]
  wire  RetimeWrapper_58_io_out; // @[package.scala 93:22:@26851.4]
  wire  RetimeWrapper_59_clock; // @[package.scala 93:22:@26863.4]
  wire  RetimeWrapper_59_reset; // @[package.scala 93:22:@26863.4]
  wire  RetimeWrapper_59_io_flow; // @[package.scala 93:22:@26863.4]
  wire  RetimeWrapper_59_io_in; // @[package.scala 93:22:@26863.4]
  wire  RetimeWrapper_59_io_out; // @[package.scala 93:22:@26863.4]
  wire  x357_1_clock; // @[Math.scala 262:24:@26886.4]
  wire [31:0] x357_1_io_a; // @[Math.scala 262:24:@26886.4]
  wire [31:0] x357_1_io_b; // @[Math.scala 262:24:@26886.4]
  wire  x357_1_io_flow; // @[Math.scala 262:24:@26886.4]
  wire [31:0] x357_1_io_result; // @[Math.scala 262:24:@26886.4]
  wire  x358_1_clock; // @[Math.scala 262:24:@26898.4]
  wire [31:0] x358_1_io_a; // @[Math.scala 262:24:@26898.4]
  wire [31:0] x358_1_io_b; // @[Math.scala 262:24:@26898.4]
  wire  x358_1_io_flow; // @[Math.scala 262:24:@26898.4]
  wire [31:0] x358_1_io_result; // @[Math.scala 262:24:@26898.4]
  wire  x359_1_clock; // @[Math.scala 262:24:@26910.4]
  wire [31:0] x359_1_io_a; // @[Math.scala 262:24:@26910.4]
  wire [31:0] x359_1_io_b; // @[Math.scala 262:24:@26910.4]
  wire  x359_1_io_flow; // @[Math.scala 262:24:@26910.4]
  wire [31:0] x359_1_io_result; // @[Math.scala 262:24:@26910.4]
  wire  x360_1_clock; // @[Math.scala 262:24:@26922.4]
  wire [31:0] x360_1_io_a; // @[Math.scala 262:24:@26922.4]
  wire [31:0] x360_1_io_b; // @[Math.scala 262:24:@26922.4]
  wire  x360_1_io_flow; // @[Math.scala 262:24:@26922.4]
  wire [31:0] x360_1_io_result; // @[Math.scala 262:24:@26922.4]
  wire  x361_1_clock; // @[Math.scala 262:24:@26934.4]
  wire [31:0] x361_1_io_a; // @[Math.scala 262:24:@26934.4]
  wire [31:0] x361_1_io_b; // @[Math.scala 262:24:@26934.4]
  wire  x361_1_io_flow; // @[Math.scala 262:24:@26934.4]
  wire [31:0] x361_1_io_result; // @[Math.scala 262:24:@26934.4]
  wire  x362_1_clock; // @[Math.scala 262:24:@26946.4]
  wire [31:0] x362_1_io_a; // @[Math.scala 262:24:@26946.4]
  wire [31:0] x362_1_io_b; // @[Math.scala 262:24:@26946.4]
  wire  x362_1_io_flow; // @[Math.scala 262:24:@26946.4]
  wire [31:0] x362_1_io_result; // @[Math.scala 262:24:@26946.4]
  wire  x363_1_clock; // @[Math.scala 262:24:@26958.4]
  wire [31:0] x363_1_io_a; // @[Math.scala 262:24:@26958.4]
  wire [31:0] x363_1_io_b; // @[Math.scala 262:24:@26958.4]
  wire  x363_1_io_flow; // @[Math.scala 262:24:@26958.4]
  wire [31:0] x363_1_io_result; // @[Math.scala 262:24:@26958.4]
  wire  x364_1_clock; // @[Math.scala 262:24:@26970.4]
  wire [31:0] x364_1_io_a; // @[Math.scala 262:24:@26970.4]
  wire [31:0] x364_1_io_b; // @[Math.scala 262:24:@26970.4]
  wire  x364_1_io_flow; // @[Math.scala 262:24:@26970.4]
  wire [31:0] x364_1_io_result; // @[Math.scala 262:24:@26970.4]
  wire  x365_1_clock; // @[Math.scala 262:24:@26982.4]
  wire [31:0] x365_1_io_a; // @[Math.scala 262:24:@26982.4]
  wire [31:0] x365_1_io_b; // @[Math.scala 262:24:@26982.4]
  wire  x365_1_io_flow; // @[Math.scala 262:24:@26982.4]
  wire [31:0] x365_1_io_result; // @[Math.scala 262:24:@26982.4]
  wire  x366_x3_1_clock; // @[Math.scala 150:24:@26992.4]
  wire  x366_x3_1_reset; // @[Math.scala 150:24:@26992.4]
  wire [31:0] x366_x3_1_io_a; // @[Math.scala 150:24:@26992.4]
  wire [31:0] x366_x3_1_io_b; // @[Math.scala 150:24:@26992.4]
  wire  x366_x3_1_io_flow; // @[Math.scala 150:24:@26992.4]
  wire [31:0] x366_x3_1_io_result; // @[Math.scala 150:24:@26992.4]
  wire  x367_x4_1_clock; // @[Math.scala 150:24:@27002.4]
  wire  x367_x4_1_reset; // @[Math.scala 150:24:@27002.4]
  wire [31:0] x367_x4_1_io_a; // @[Math.scala 150:24:@27002.4]
  wire [31:0] x367_x4_1_io_b; // @[Math.scala 150:24:@27002.4]
  wire  x367_x4_1_io_flow; // @[Math.scala 150:24:@27002.4]
  wire [31:0] x367_x4_1_io_result; // @[Math.scala 150:24:@27002.4]
  wire  x368_x3_1_clock; // @[Math.scala 150:24:@27012.4]
  wire  x368_x3_1_reset; // @[Math.scala 150:24:@27012.4]
  wire [31:0] x368_x3_1_io_a; // @[Math.scala 150:24:@27012.4]
  wire [31:0] x368_x3_1_io_b; // @[Math.scala 150:24:@27012.4]
  wire  x368_x3_1_io_flow; // @[Math.scala 150:24:@27012.4]
  wire [31:0] x368_x3_1_io_result; // @[Math.scala 150:24:@27012.4]
  wire  x369_x4_1_clock; // @[Math.scala 150:24:@27022.4]
  wire  x369_x4_1_reset; // @[Math.scala 150:24:@27022.4]
  wire [31:0] x369_x4_1_io_a; // @[Math.scala 150:24:@27022.4]
  wire [31:0] x369_x4_1_io_b; // @[Math.scala 150:24:@27022.4]
  wire  x369_x4_1_io_flow; // @[Math.scala 150:24:@27022.4]
  wire [31:0] x369_x4_1_io_result; // @[Math.scala 150:24:@27022.4]
  wire  x370_x3_1_clock; // @[Math.scala 150:24:@27032.4]
  wire  x370_x3_1_reset; // @[Math.scala 150:24:@27032.4]
  wire [31:0] x370_x3_1_io_a; // @[Math.scala 150:24:@27032.4]
  wire [31:0] x370_x3_1_io_b; // @[Math.scala 150:24:@27032.4]
  wire  x370_x3_1_io_flow; // @[Math.scala 150:24:@27032.4]
  wire [31:0] x370_x3_1_io_result; // @[Math.scala 150:24:@27032.4]
  wire  x371_x4_1_clock; // @[Math.scala 150:24:@27042.4]
  wire  x371_x4_1_reset; // @[Math.scala 150:24:@27042.4]
  wire [31:0] x371_x4_1_io_a; // @[Math.scala 150:24:@27042.4]
  wire [31:0] x371_x4_1_io_b; // @[Math.scala 150:24:@27042.4]
  wire  x371_x4_1_io_flow; // @[Math.scala 150:24:@27042.4]
  wire [31:0] x371_x4_1_io_result; // @[Math.scala 150:24:@27042.4]
  wire  x372_x3_1_clock; // @[Math.scala 150:24:@27052.4]
  wire  x372_x3_1_reset; // @[Math.scala 150:24:@27052.4]
  wire [31:0] x372_x3_1_io_a; // @[Math.scala 150:24:@27052.4]
  wire [31:0] x372_x3_1_io_b; // @[Math.scala 150:24:@27052.4]
  wire  x372_x3_1_io_flow; // @[Math.scala 150:24:@27052.4]
  wire [31:0] x372_x3_1_io_result; // @[Math.scala 150:24:@27052.4]
  wire  RetimeWrapper_60_clock; // @[package.scala 93:22:@27062.4]
  wire  RetimeWrapper_60_reset; // @[package.scala 93:22:@27062.4]
  wire  RetimeWrapper_60_io_flow; // @[package.scala 93:22:@27062.4]
  wire [31:0] RetimeWrapper_60_io_in; // @[package.scala 93:22:@27062.4]
  wire [31:0] RetimeWrapper_60_io_out; // @[package.scala 93:22:@27062.4]
  wire  x373_sum_1_clock; // @[Math.scala 150:24:@27071.4]
  wire  x373_sum_1_reset; // @[Math.scala 150:24:@27071.4]
  wire [31:0] x373_sum_1_io_a; // @[Math.scala 150:24:@27071.4]
  wire [31:0] x373_sum_1_io_b; // @[Math.scala 150:24:@27071.4]
  wire  x373_sum_1_io_flow; // @[Math.scala 150:24:@27071.4]
  wire [31:0] x373_sum_1_io_result; // @[Math.scala 150:24:@27071.4]
  wire [31:0] x374_1_io_b; // @[Math.scala 720:24:@27081.4]
  wire [31:0] x374_1_io_result; // @[Math.scala 720:24:@27081.4]
  wire  x375_mul_1_clock; // @[Math.scala 262:24:@27092.4]
  wire [31:0] x375_mul_1_io_a; // @[Math.scala 262:24:@27092.4]
  wire  x375_mul_1_io_flow; // @[Math.scala 262:24:@27092.4]
  wire [31:0] x375_mul_1_io_result; // @[Math.scala 262:24:@27092.4]
  wire [31:0] x376_1_io_b; // @[Math.scala 720:24:@27102.4]
  wire [31:0] x376_1_io_result; // @[Math.scala 720:24:@27102.4]
  wire  x377_1_clock; // @[Math.scala 262:24:@27113.4]
  wire [31:0] x377_1_io_a; // @[Math.scala 262:24:@27113.4]
  wire [31:0] x377_1_io_b; // @[Math.scala 262:24:@27113.4]
  wire  x377_1_io_flow; // @[Math.scala 262:24:@27113.4]
  wire [31:0] x377_1_io_result; // @[Math.scala 262:24:@27113.4]
  wire  x378_1_clock; // @[Math.scala 262:24:@27125.4]
  wire [31:0] x378_1_io_a; // @[Math.scala 262:24:@27125.4]
  wire [31:0] x378_1_io_b; // @[Math.scala 262:24:@27125.4]
  wire  x378_1_io_flow; // @[Math.scala 262:24:@27125.4]
  wire [31:0] x378_1_io_result; // @[Math.scala 262:24:@27125.4]
  wire  x379_1_clock; // @[Math.scala 262:24:@27137.4]
  wire [31:0] x379_1_io_a; // @[Math.scala 262:24:@27137.4]
  wire [31:0] x379_1_io_b; // @[Math.scala 262:24:@27137.4]
  wire  x379_1_io_flow; // @[Math.scala 262:24:@27137.4]
  wire [31:0] x379_1_io_result; // @[Math.scala 262:24:@27137.4]
  wire  x380_1_clock; // @[Math.scala 262:24:@27149.4]
  wire [31:0] x380_1_io_a; // @[Math.scala 262:24:@27149.4]
  wire [31:0] x380_1_io_b; // @[Math.scala 262:24:@27149.4]
  wire  x380_1_io_flow; // @[Math.scala 262:24:@27149.4]
  wire [31:0] x380_1_io_result; // @[Math.scala 262:24:@27149.4]
  wire  x381_1_clock; // @[Math.scala 262:24:@27161.4]
  wire [31:0] x381_1_io_a; // @[Math.scala 262:24:@27161.4]
  wire [31:0] x381_1_io_b; // @[Math.scala 262:24:@27161.4]
  wire  x381_1_io_flow; // @[Math.scala 262:24:@27161.4]
  wire [31:0] x381_1_io_result; // @[Math.scala 262:24:@27161.4]
  wire  x382_1_clock; // @[Math.scala 262:24:@27173.4]
  wire [31:0] x382_1_io_a; // @[Math.scala 262:24:@27173.4]
  wire [31:0] x382_1_io_b; // @[Math.scala 262:24:@27173.4]
  wire  x382_1_io_flow; // @[Math.scala 262:24:@27173.4]
  wire [31:0] x382_1_io_result; // @[Math.scala 262:24:@27173.4]
  wire  x383_1_clock; // @[Math.scala 262:24:@27185.4]
  wire [31:0] x383_1_io_a; // @[Math.scala 262:24:@27185.4]
  wire [31:0] x383_1_io_b; // @[Math.scala 262:24:@27185.4]
  wire  x383_1_io_flow; // @[Math.scala 262:24:@27185.4]
  wire [31:0] x383_1_io_result; // @[Math.scala 262:24:@27185.4]
  wire  x384_1_clock; // @[Math.scala 262:24:@27197.4]
  wire [31:0] x384_1_io_a; // @[Math.scala 262:24:@27197.4]
  wire [31:0] x384_1_io_b; // @[Math.scala 262:24:@27197.4]
  wire  x384_1_io_flow; // @[Math.scala 262:24:@27197.4]
  wire [31:0] x384_1_io_result; // @[Math.scala 262:24:@27197.4]
  wire  x385_1_clock; // @[Math.scala 262:24:@27209.4]
  wire [31:0] x385_1_io_a; // @[Math.scala 262:24:@27209.4]
  wire [31:0] x385_1_io_b; // @[Math.scala 262:24:@27209.4]
  wire  x385_1_io_flow; // @[Math.scala 262:24:@27209.4]
  wire [31:0] x385_1_io_result; // @[Math.scala 262:24:@27209.4]
  wire  x386_x3_1_clock; // @[Math.scala 150:24:@27219.4]
  wire  x386_x3_1_reset; // @[Math.scala 150:24:@27219.4]
  wire [31:0] x386_x3_1_io_a; // @[Math.scala 150:24:@27219.4]
  wire [31:0] x386_x3_1_io_b; // @[Math.scala 150:24:@27219.4]
  wire  x386_x3_1_io_flow; // @[Math.scala 150:24:@27219.4]
  wire [31:0] x386_x3_1_io_result; // @[Math.scala 150:24:@27219.4]
  wire  x387_x4_1_clock; // @[Math.scala 150:24:@27229.4]
  wire  x387_x4_1_reset; // @[Math.scala 150:24:@27229.4]
  wire [31:0] x387_x4_1_io_a; // @[Math.scala 150:24:@27229.4]
  wire [31:0] x387_x4_1_io_b; // @[Math.scala 150:24:@27229.4]
  wire  x387_x4_1_io_flow; // @[Math.scala 150:24:@27229.4]
  wire [31:0] x387_x4_1_io_result; // @[Math.scala 150:24:@27229.4]
  wire  x388_x3_1_clock; // @[Math.scala 150:24:@27239.4]
  wire  x388_x3_1_reset; // @[Math.scala 150:24:@27239.4]
  wire [31:0] x388_x3_1_io_a; // @[Math.scala 150:24:@27239.4]
  wire [31:0] x388_x3_1_io_b; // @[Math.scala 150:24:@27239.4]
  wire  x388_x3_1_io_flow; // @[Math.scala 150:24:@27239.4]
  wire [31:0] x388_x3_1_io_result; // @[Math.scala 150:24:@27239.4]
  wire  x389_x4_1_clock; // @[Math.scala 150:24:@27249.4]
  wire  x389_x4_1_reset; // @[Math.scala 150:24:@27249.4]
  wire [31:0] x389_x4_1_io_a; // @[Math.scala 150:24:@27249.4]
  wire [31:0] x389_x4_1_io_b; // @[Math.scala 150:24:@27249.4]
  wire  x389_x4_1_io_flow; // @[Math.scala 150:24:@27249.4]
  wire [31:0] x389_x4_1_io_result; // @[Math.scala 150:24:@27249.4]
  wire  x390_x3_1_clock; // @[Math.scala 150:24:@27259.4]
  wire  x390_x3_1_reset; // @[Math.scala 150:24:@27259.4]
  wire [31:0] x390_x3_1_io_a; // @[Math.scala 150:24:@27259.4]
  wire [31:0] x390_x3_1_io_b; // @[Math.scala 150:24:@27259.4]
  wire  x390_x3_1_io_flow; // @[Math.scala 150:24:@27259.4]
  wire [31:0] x390_x3_1_io_result; // @[Math.scala 150:24:@27259.4]
  wire  x391_x4_1_clock; // @[Math.scala 150:24:@27269.4]
  wire  x391_x4_1_reset; // @[Math.scala 150:24:@27269.4]
  wire [31:0] x391_x4_1_io_a; // @[Math.scala 150:24:@27269.4]
  wire [31:0] x391_x4_1_io_b; // @[Math.scala 150:24:@27269.4]
  wire  x391_x4_1_io_flow; // @[Math.scala 150:24:@27269.4]
  wire [31:0] x391_x4_1_io_result; // @[Math.scala 150:24:@27269.4]
  wire  x392_x3_1_clock; // @[Math.scala 150:24:@27279.4]
  wire  x392_x3_1_reset; // @[Math.scala 150:24:@27279.4]
  wire [31:0] x392_x3_1_io_a; // @[Math.scala 150:24:@27279.4]
  wire [31:0] x392_x3_1_io_b; // @[Math.scala 150:24:@27279.4]
  wire  x392_x3_1_io_flow; // @[Math.scala 150:24:@27279.4]
  wire [31:0] x392_x3_1_io_result; // @[Math.scala 150:24:@27279.4]
  wire  RetimeWrapper_61_clock; // @[package.scala 93:22:@27289.4]
  wire  RetimeWrapper_61_reset; // @[package.scala 93:22:@27289.4]
  wire  RetimeWrapper_61_io_flow; // @[package.scala 93:22:@27289.4]
  wire [31:0] RetimeWrapper_61_io_in; // @[package.scala 93:22:@27289.4]
  wire [31:0] RetimeWrapper_61_io_out; // @[package.scala 93:22:@27289.4]
  wire  x393_sum_1_clock; // @[Math.scala 150:24:@27298.4]
  wire  x393_sum_1_reset; // @[Math.scala 150:24:@27298.4]
  wire [31:0] x393_sum_1_io_a; // @[Math.scala 150:24:@27298.4]
  wire [31:0] x393_sum_1_io_b; // @[Math.scala 150:24:@27298.4]
  wire  x393_sum_1_io_flow; // @[Math.scala 150:24:@27298.4]
  wire [31:0] x393_sum_1_io_result; // @[Math.scala 150:24:@27298.4]
  wire [31:0] x394_1_io_b; // @[Math.scala 720:24:@27308.4]
  wire [31:0] x394_1_io_result; // @[Math.scala 720:24:@27308.4]
  wire  x395_mul_1_clock; // @[Math.scala 262:24:@27319.4]
  wire [31:0] x395_mul_1_io_a; // @[Math.scala 262:24:@27319.4]
  wire  x395_mul_1_io_flow; // @[Math.scala 262:24:@27319.4]
  wire [31:0] x395_mul_1_io_result; // @[Math.scala 262:24:@27319.4]
  wire [31:0] x396_1_io_b; // @[Math.scala 720:24:@27329.4]
  wire [31:0] x396_1_io_result; // @[Math.scala 720:24:@27329.4]
  wire  RetimeWrapper_62_clock; // @[package.scala 93:22:@27344.4]
  wire  RetimeWrapper_62_reset; // @[package.scala 93:22:@27344.4]
  wire  RetimeWrapper_62_io_flow; // @[package.scala 93:22:@27344.4]
  wire [63:0] RetimeWrapper_62_io_in; // @[package.scala 93:22:@27344.4]
  wire [63:0] RetimeWrapper_62_io_out; // @[package.scala 93:22:@27344.4]
  wire  RetimeWrapper_63_clock; // @[package.scala 93:22:@27353.4]
  wire  RetimeWrapper_63_reset; // @[package.scala 93:22:@27353.4]
  wire  RetimeWrapper_63_io_flow; // @[package.scala 93:22:@27353.4]
  wire  RetimeWrapper_63_io_in; // @[package.scala 93:22:@27353.4]
  wire  RetimeWrapper_63_io_out; // @[package.scala 93:22:@27353.4]
  wire  RetimeWrapper_64_clock; // @[package.scala 93:22:@27362.4]
  wire  RetimeWrapper_64_reset; // @[package.scala 93:22:@27362.4]
  wire  RetimeWrapper_64_io_flow; // @[package.scala 93:22:@27362.4]
  wire  RetimeWrapper_64_io_in; // @[package.scala 93:22:@27362.4]
  wire  RetimeWrapper_64_io_out; // @[package.scala 93:22:@27362.4]
  wire  RetimeWrapper_65_clock; // @[package.scala 93:22:@27371.4]
  wire  RetimeWrapper_65_reset; // @[package.scala 93:22:@27371.4]
  wire  RetimeWrapper_65_io_flow; // @[package.scala 93:22:@27371.4]
  wire  RetimeWrapper_65_io_in; // @[package.scala 93:22:@27371.4]
  wire  RetimeWrapper_65_io_out; // @[package.scala 93:22:@27371.4]
  wire  b254; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 62:18:@25419.4]
  wire  b255; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 63:18:@25420.4]
  wire  _T_205; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 67:30:@25422.4]
  wire  _T_206; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 67:37:@25423.4]
  wire  _T_210; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 69:76:@25428.4]
  wire  _T_211; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 69:62:@25429.4]
  wire  _T_213; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 69:101:@25430.4]
  wire [63:0] x483_x256_D1_0_number; // @[package.scala 96:25:@25439.4 package.scala 96:25:@25440.4]
  wire [31:0] b252_number; // @[Math.scala 723:22:@25404.4 Math.scala 724:14:@25405.4]
  wire [31:0] _T_243; // @[Math.scala 406:49:@25548.4]
  wire [31:0] _T_245; // @[Math.scala 406:56:@25550.4]
  wire [31:0] _T_246; // @[Math.scala 406:56:@25551.4]
  wire [31:0] x459_number; // @[implicits.scala 133:21:@25552.4]
  wire [31:0] _T_256; // @[Math.scala 406:49:@25561.4]
  wire [31:0] _T_258; // @[Math.scala 406:56:@25563.4]
  wire [31:0] _T_259; // @[Math.scala 406:56:@25564.4]
  wire [31:0] b253_number; // @[Math.scala 723:22:@25416.4 Math.scala 724:14:@25417.4]
  wire [31:0] _T_268; // @[Math.scala 406:49:@25572.4]
  wire [31:0] _T_270; // @[Math.scala 406:56:@25574.4]
  wire [31:0] _T_271; // @[Math.scala 406:56:@25575.4]
  wire  _T_275; // @[FixedPoint.scala 50:25:@25581.4]
  wire [1:0] _T_279; // @[Bitwise.scala 72:12:@25583.4]
  wire [29:0] _T_280; // @[FixedPoint.scala 18:52:@25584.4]
  wire  _T_286; // @[Math.scala 451:55:@25586.4]
  wire [1:0] _T_287; // @[FixedPoint.scala 18:52:@25587.4]
  wire  _T_293; // @[Math.scala 451:110:@25589.4]
  wire  _T_294; // @[Math.scala 451:94:@25590.4]
  wire [31:0] _T_296; // @[Cat.scala 30:58:@25592.4]
  wire [31:0] x264_1_number; // @[Math.scala 454:20:@25593.4]
  wire [40:0] _GEN_0; // @[Math.scala 461:32:@25598.4]
  wire [40:0] _T_301; // @[Math.scala 461:32:@25598.4]
  wire [36:0] _GEN_1; // @[Math.scala 461:32:@25603.4]
  wire [36:0] _T_304; // @[Math.scala 461:32:@25603.4]
  wire  _T_310; // @[FixedPoint.scala 50:25:@25618.4]
  wire [1:0] _T_314; // @[Bitwise.scala 72:12:@25620.4]
  wire [29:0] _T_315; // @[FixedPoint.scala 18:52:@25621.4]
  wire  _T_321; // @[Math.scala 451:55:@25623.4]
  wire [1:0] _T_322; // @[FixedPoint.scala 18:52:@25624.4]
  wire  _T_328; // @[Math.scala 451:110:@25626.4]
  wire  _T_329; // @[Math.scala 451:94:@25627.4]
  wire [31:0] _T_331; // @[Cat.scala 30:58:@25629.4]
  wire  _T_359; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:101:@25706.4]
  wire  _T_363; // @[package.scala 96:25:@25714.4 package.scala 96:25:@25715.4]
  wire  _T_365; // @[implicits.scala 55:10:@25716.4]
  wire  _T_366; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:118:@25717.4]
  wire  _T_368; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:206:@25719.4]
  wire  _T_369; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:225:@25720.4]
  wire  x490_b254_D3; // @[package.scala 96:25:@25703.4 package.scala 96:25:@25704.4]
  wire  _T_370; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:251:@25721.4]
  wire  x489_b255_D3; // @[package.scala 96:25:@25694.4 package.scala 96:25:@25695.4]
  wire [31:0] x269_rdcol_number; // @[Math.scala 154:22:@25738.4 Math.scala 155:14:@25739.4]
  wire [31:0] _T_387; // @[Math.scala 406:49:@25747.4]
  wire [31:0] _T_389; // @[Math.scala 406:56:@25749.4]
  wire [31:0] _T_390; // @[Math.scala 406:56:@25750.4]
  wire  _T_394; // @[FixedPoint.scala 50:25:@25756.4]
  wire [1:0] _T_398; // @[Bitwise.scala 72:12:@25758.4]
  wire [29:0] _T_399; // @[FixedPoint.scala 18:52:@25759.4]
  wire  _T_405; // @[Math.scala 451:55:@25761.4]
  wire [1:0] _T_406; // @[FixedPoint.scala 18:52:@25762.4]
  wire  _T_412; // @[Math.scala 451:110:@25764.4]
  wire  _T_413; // @[Math.scala 451:94:@25765.4]
  wire [31:0] _T_415; // @[Cat.scala 30:58:@25767.4]
  wire  _T_435; // @[package.scala 96:25:@25816.4 package.scala 96:25:@25817.4]
  wire  _T_437; // @[implicits.scala 55:10:@25818.4]
  wire  _T_438; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 138:118:@25819.4]
  wire  _T_440; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 138:206:@25821.4]
  wire  _T_441; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 138:225:@25822.4]
  wire  _T_442; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 138:251:@25823.4]
  wire [31:0] x494_b252_D6_number; // @[package.scala 96:25:@25837.4 package.scala 96:25:@25838.4]
  wire [31:0] _T_452; // @[Math.scala 476:37:@25843.4]
  wire  x276; // @[Math.scala 476:44:@25845.4]
  wire [31:0] x495_x269_rdcol_D6_number; // @[package.scala 96:25:@25853.4 package.scala 96:25:@25854.4]
  wire [31:0] _T_463; // @[Math.scala 476:37:@25859.4]
  wire  x277; // @[Math.scala 476:44:@25861.4]
  wire  x496_x276_D1; // @[package.scala 96:25:@25869.4 package.scala 96:25:@25870.4]
  wire  x278; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 151:24:@25873.4]
  wire  _T_502; // @[package.scala 96:25:@25941.4 package.scala 96:25:@25942.4]
  wire  _T_504; // @[implicits.scala 55:10:@25943.4]
  wire  _T_505; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 170:146:@25944.4]
  wire  x498_x279_D2; // @[package.scala 96:25:@25893.4 package.scala 96:25:@25894.4]
  wire  _T_506; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 170:234:@25945.4]
  wire  x502_b254_D9; // @[package.scala 96:25:@25929.4 package.scala 96:25:@25930.4]
  wire  _T_507; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 170:242:@25946.4]
  wire  x499_b255_D9; // @[package.scala 96:25:@25902.4 package.scala 96:25:@25903.4]
  wire [31:0] x503_b253_D6_number; // @[package.scala 96:25:@25962.4 package.scala 96:25:@25963.4]
  wire [31:0] _T_520; // @[Math.scala 476:37:@25970.4]
  wire  x282; // @[Math.scala 476:44:@25972.4]
  wire  x283; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 186:59:@25975.4]
  wire  _T_547; // @[package.scala 96:25:@26016.4 package.scala 96:25:@26017.4]
  wire  _T_549; // @[implicits.scala 55:10:@26018.4]
  wire  _T_550; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 199:194:@26019.4]
  wire  x504_x284_D3; // @[package.scala 96:25:@25986.4 package.scala 96:25:@25987.4]
  wire  _T_551; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 199:282:@26020.4]
  wire  _T_552; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 199:290:@26021.4]
  wire [31:0] x287_rdcol_number; // @[Math.scala 154:22:@26040.4 Math.scala 155:14:@26041.4]
  wire [31:0] _T_567; // @[Math.scala 476:37:@26046.4]
  wire  x288; // @[Math.scala 476:44:@26048.4]
  wire  x289; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 207:59:@26051.4]
  wire [31:0] _T_583; // @[Math.scala 406:56:@26062.4]
  wire [31:0] _T_584; // @[Math.scala 406:56:@26063.4]
  wire  _T_588; // @[FixedPoint.scala 50:25:@26069.4]
  wire [1:0] _T_592; // @[Bitwise.scala 72:12:@26071.4]
  wire [29:0] _T_593; // @[FixedPoint.scala 18:52:@26072.4]
  wire  _T_599; // @[Math.scala 451:55:@26074.4]
  wire [1:0] _T_600; // @[FixedPoint.scala 18:52:@26075.4]
  wire  _T_606; // @[Math.scala 451:110:@26077.4]
  wire  _T_607; // @[Math.scala 451:94:@26078.4]
  wire [31:0] _T_609; // @[Cat.scala 30:58:@26080.4]
  wire  _T_638; // @[package.scala 96:25:@26139.4 package.scala 96:25:@26140.4]
  wire  _T_640; // @[implicits.scala 55:10:@26141.4]
  wire  _T_641; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 228:194:@26142.4]
  wire  x510_x290_D2; // @[package.scala 96:25:@26127.4 package.scala 96:25:@26128.4]
  wire  _T_642; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 228:282:@26143.4]
  wire  _T_643; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 228:290:@26144.4]
  wire [31:0] x296_rdcol_number; // @[Math.scala 154:22:@26163.4 Math.scala 155:14:@26164.4]
  wire [31:0] _T_658; // @[Math.scala 476:37:@26169.4]
  wire  x297; // @[Math.scala 476:44:@26171.4]
  wire  x298; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 236:59:@26174.4]
  wire [31:0] _T_674; // @[Math.scala 406:56:@26185.4]
  wire [31:0] _T_675; // @[Math.scala 406:56:@26186.4]
  wire  _T_679; // @[FixedPoint.scala 50:25:@26192.4]
  wire [1:0] _T_683; // @[Bitwise.scala 72:12:@26194.4]
  wire [29:0] _T_684; // @[FixedPoint.scala 18:52:@26195.4]
  wire  _T_690; // @[Math.scala 451:55:@26197.4]
  wire [1:0] _T_691; // @[FixedPoint.scala 18:52:@26198.4]
  wire  _T_697; // @[Math.scala 451:110:@26200.4]
  wire  _T_698; // @[Math.scala 451:94:@26201.4]
  wire [31:0] _T_700; // @[Cat.scala 30:58:@26203.4]
  wire  _T_726; // @[package.scala 96:25:@26253.4 package.scala 96:25:@26254.4]
  wire  _T_728; // @[implicits.scala 55:10:@26255.4]
  wire  _T_729; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 255:194:@26256.4]
  wire  x513_x299_D2; // @[package.scala 96:25:@26241.4 package.scala 96:25:@26242.4]
  wire  _T_730; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 255:282:@26257.4]
  wire  _T_731; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 255:290:@26258.4]
  wire [31:0] x305_rdrow_number; // @[Math.scala 195:22:@26277.4 Math.scala 196:14:@26278.4]
  wire [31:0] _T_748; // @[Math.scala 406:49:@26284.4]
  wire [31:0] _T_750; // @[Math.scala 406:56:@26286.4]
  wire [31:0] _T_751; // @[Math.scala 406:56:@26287.4]
  wire [31:0] x468_number; // @[implicits.scala 133:21:@26288.4]
  wire  x307; // @[Math.scala 476:44:@26296.4]
  wire  x308; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 265:24:@26299.4]
  wire [31:0] _T_772; // @[Math.scala 406:49:@26308.4]
  wire [31:0] _T_774; // @[Math.scala 406:56:@26310.4]
  wire [31:0] _T_775; // @[Math.scala 406:56:@26311.4]
  wire  _T_779; // @[FixedPoint.scala 50:25:@26317.4]
  wire [1:0] _T_783; // @[Bitwise.scala 72:12:@26319.4]
  wire [29:0] _T_784; // @[FixedPoint.scala 18:52:@26320.4]
  wire  _T_790; // @[Math.scala 451:55:@26322.4]
  wire [1:0] _T_791; // @[FixedPoint.scala 18:52:@26323.4]
  wire  _T_797; // @[Math.scala 451:110:@26325.4]
  wire  _T_798; // @[Math.scala 451:94:@26326.4]
  wire [31:0] _T_800; // @[Cat.scala 30:58:@26328.4]
  wire [31:0] x311_1_number; // @[Math.scala 454:20:@26329.4]
  wire [40:0] _GEN_2; // @[Math.scala 461:32:@26334.4]
  wire [40:0] _T_805; // @[Math.scala 461:32:@26334.4]
  wire [36:0] _GEN_3; // @[Math.scala 461:32:@26339.4]
  wire [36:0] _T_808; // @[Math.scala 461:32:@26339.4]
  wire  _T_835; // @[package.scala 96:25:@26398.4 package.scala 96:25:@26399.4]
  wire  _T_837; // @[implicits.scala 55:10:@26400.4]
  wire  _T_838; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 290:194:@26401.4]
  wire  x516_x309_D2; // @[package.scala 96:25:@26386.4 package.scala 96:25:@26387.4]
  wire  _T_839; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 290:282:@26402.4]
  wire  _T_840; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 290:290:@26403.4]
  wire  x517_x282_D1; // @[package.scala 96:25:@26419.4 package.scala 96:25:@26420.4]
  wire  x316; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 302:59:@26423.4]
  wire  _T_872; // @[package.scala 96:25:@26467.4 package.scala 96:25:@26468.4]
  wire  _T_874; // @[implicits.scala 55:10:@26469.4]
  wire  _T_875; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 317:194:@26470.4]
  wire  x519_x317_D2; // @[package.scala 96:25:@26455.4 package.scala 96:25:@26456.4]
  wire  _T_876; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 317:282:@26471.4]
  wire  _T_877; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 317:290:@26472.4]
  wire  x321; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 321:59:@26483.4]
  wire  _T_904; // @[package.scala 96:25:@26525.4 package.scala 96:25:@26526.4]
  wire  _T_906; // @[implicits.scala 55:10:@26527.4]
  wire  _T_907; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 334:194:@26528.4]
  wire  x521_x322_D2; // @[package.scala 96:25:@26513.4 package.scala 96:25:@26514.4]
  wire  _T_908; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 334:282:@26529.4]
  wire  _T_909; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 334:290:@26530.4]
  wire  x326; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 338:59:@26541.4]
  wire  _T_936; // @[package.scala 96:25:@26583.4 package.scala 96:25:@26584.4]
  wire  _T_938; // @[implicits.scala 55:10:@26585.4]
  wire  _T_939; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 351:194:@26586.4]
  wire  x523_x327_D2; // @[package.scala 96:25:@26571.4 package.scala 96:25:@26572.4]
  wire  _T_940; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 351:282:@26587.4]
  wire  _T_941; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 351:290:@26588.4]
  wire [31:0] x331_rdrow_number; // @[Math.scala 195:22:@26607.4 Math.scala 196:14:@26608.4]
  wire [31:0] _T_958; // @[Math.scala 406:49:@26614.4]
  wire [31:0] _T_960; // @[Math.scala 406:56:@26616.4]
  wire [31:0] _T_961; // @[Math.scala 406:56:@26617.4]
  wire [31:0] x473_number; // @[implicits.scala 133:21:@26618.4]
  wire  x333; // @[Math.scala 476:44:@26626.4]
  wire  x334; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 361:24:@26629.4]
  wire [31:0] _T_982; // @[Math.scala 406:49:@26638.4]
  wire [31:0] _T_984; // @[Math.scala 406:56:@26640.4]
  wire [31:0] _T_985; // @[Math.scala 406:56:@26641.4]
  wire  _T_989; // @[FixedPoint.scala 50:25:@26647.4]
  wire [1:0] _T_993; // @[Bitwise.scala 72:12:@26649.4]
  wire [29:0] _T_994; // @[FixedPoint.scala 18:52:@26650.4]
  wire  _T_1000; // @[Math.scala 451:55:@26652.4]
  wire [1:0] _T_1001; // @[FixedPoint.scala 18:52:@26653.4]
  wire  _T_1007; // @[Math.scala 451:110:@26655.4]
  wire  _T_1008; // @[Math.scala 451:94:@26656.4]
  wire [31:0] _T_1010; // @[Cat.scala 30:58:@26658.4]
  wire [31:0] x337_1_number; // @[Math.scala 454:20:@26659.4]
  wire [40:0] _GEN_4; // @[Math.scala 461:32:@26664.4]
  wire [40:0] _T_1015; // @[Math.scala 461:32:@26664.4]
  wire [36:0] _GEN_5; // @[Math.scala 461:32:@26669.4]
  wire [36:0] _T_1018; // @[Math.scala 461:32:@26669.4]
  wire  _T_1042; // @[package.scala 96:25:@26719.4 package.scala 96:25:@26720.4]
  wire  _T_1044; // @[implicits.scala 55:10:@26721.4]
  wire  _T_1045; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 384:194:@26722.4]
  wire  x524_x335_D2; // @[package.scala 96:25:@26698.4 package.scala 96:25:@26699.4]
  wire  _T_1046; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 384:282:@26723.4]
  wire  _T_1047; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 384:290:@26724.4]
  wire  x342; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 388:24:@26735.4]
  wire  _T_1071; // @[package.scala 96:25:@26768.4 package.scala 96:25:@26769.4]
  wire  _T_1073; // @[implicits.scala 55:10:@26770.4]
  wire  _T_1074; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 399:194:@26771.4]
  wire  x526_x343_D2; // @[package.scala 96:25:@26756.4 package.scala 96:25:@26757.4]
  wire  _T_1075; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 399:282:@26772.4]
  wire  _T_1076; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 399:290:@26773.4]
  wire  x347; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 403:24:@26784.4]
  wire  _T_1100; // @[package.scala 96:25:@26817.4 package.scala 96:25:@26818.4]
  wire  _T_1102; // @[implicits.scala 55:10:@26819.4]
  wire  _T_1103; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 414:194:@26820.4]
  wire  x527_x348_D2; // @[package.scala 96:25:@26805.4 package.scala 96:25:@26806.4]
  wire  _T_1104; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 414:282:@26821.4]
  wire  _T_1105; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 414:290:@26822.4]
  wire  x352; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 424:59:@26833.4]
  wire  _T_1131; // @[package.scala 96:25:@26868.4 package.scala 96:25:@26869.4]
  wire  _T_1133; // @[implicits.scala 55:10:@26870.4]
  wire  _T_1134; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 437:194:@26871.4]
  wire  x528_x353_D2; // @[package.scala 96:25:@26856.4 package.scala 96:25:@26857.4]
  wire  _T_1135; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 437:282:@26872.4]
  wire  _T_1136; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 437:290:@26873.4]
  wire [31:0] x376_number; // @[Math.scala 723:22:@27107.4 Math.scala 724:14:@27108.4]
  wire [31:0] x396_number; // @[Math.scala 723:22:@27334.4 Math.scala 724:14:@27335.4]
  wire  _T_1366; // @[package.scala 96:25:@27376.4 package.scala 96:25:@27377.4]
  wire  _T_1368; // @[implicits.scala 55:10:@27378.4]
  wire  x531_b254_D30; // @[package.scala 96:25:@27358.4 package.scala 96:25:@27359.4]
  wire  _T_1369; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 539:117:@27379.4]
  wire  x532_b255_D30; // @[package.scala 96:25:@27367.4 package.scala 96:25:@27368.4]
  wire  _T_1370; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 539:123:@27380.4]
  wire [31:0] x485_x460_D3_number; // @[package.scala 96:25:@25658.4 package.scala 96:25:@25659.4]
  wire [31:0] x487_x461_D3_number; // @[package.scala 96:25:@25676.4 package.scala 96:25:@25677.4]
  wire [31:0] x488_x267_sum_D1_number; // @[package.scala 96:25:@25685.4 package.scala 96:25:@25686.4]
  wire [31:0] x492_x465_D2_number; // @[package.scala 96:25:@25796.4 package.scala 96:25:@25797.4]
  wire [31:0] x493_x273_sum_D1_number; // @[package.scala 96:25:@25805.4 package.scala 96:25:@25806.4]
  wire [31:0] x497_x460_D9_number; // @[package.scala 96:25:@25884.4 package.scala 96:25:@25885.4]
  wire [31:0] x500_x465_D8_number; // @[package.scala 96:25:@25911.4 package.scala 96:25:@25912.4]
  wire [31:0] x501_x273_sum_D7_number; // @[package.scala 96:25:@25920.4 package.scala 96:25:@25921.4]
  wire [31:0] x505_x461_D9_number; // @[package.scala 96:25:@25995.4 package.scala 96:25:@25996.4]
  wire [31:0] x506_x267_sum_D7_number; // @[package.scala 96:25:@26004.4 package.scala 96:25:@26005.4]
  wire [31:0] x508_x293_sum_D1_number; // @[package.scala 96:25:@26109.4 package.scala 96:25:@26110.4]
  wire [31:0] x509_x466_D2_number; // @[package.scala 96:25:@26118.4 package.scala 96:25:@26119.4]
  wire [31:0] x511_x302_sum_D1_number; // @[package.scala 96:25:@26223.4 package.scala 96:25:@26224.4]
  wire [31:0] x512_x467_D2_number; // @[package.scala 96:25:@26232.4 package.scala 96:25:@26233.4]
  wire [31:0] x313_sum_number; // @[Math.scala 154:22:@26368.4 Math.scala 155:14:@26369.4]
  wire [31:0] x515_x469_D2_number; // @[package.scala 96:25:@26377.4 package.scala 96:25:@26378.4]
  wire [31:0] x318_sum_number; // @[Math.scala 154:22:@26446.4 Math.scala 155:14:@26447.4]
  wire [31:0] x323_sum_number; // @[Math.scala 154:22:@26504.4 Math.scala 155:14:@26505.4]
  wire [31:0] x328_sum_number; // @[Math.scala 154:22:@26562.4 Math.scala 155:14:@26563.4]
  wire [31:0] x339_sum_number; // @[Math.scala 154:22:@26689.4 Math.scala 155:14:@26690.4]
  wire [31:0] x525_x474_D2_number; // @[package.scala 96:25:@26707.4 package.scala 96:25:@26708.4]
  wire [31:0] x344_sum_number; // @[Math.scala 154:22:@26747.4 Math.scala 155:14:@26748.4]
  wire [31:0] x349_sum_number; // @[Math.scala 154:22:@26796.4 Math.scala 155:14:@26797.4]
  wire [31:0] x354_sum_number; // @[Math.scala 154:22:@26847.4 Math.scala 155:14:@26848.4]
  _ _ ( // @[Math.scala 720:24:@25399.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  _ __1 ( // @[Math.scala 720:24:@25411.4]
    .io_b(__1_io_b),
    .io_result(__1_io_result)
  );
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@25434.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  x258_lb_0 x258_lb_0 ( // @[m_x258_lb_0.scala 39:17:@25444.4]
    .clock(x258_lb_0_clock),
    .reset(x258_lb_0_reset),
    .io_rPort_11_banks_1(x258_lb_0_io_rPort_11_banks_1),
    .io_rPort_11_banks_0(x258_lb_0_io_rPort_11_banks_0),
    .io_rPort_11_ofs_0(x258_lb_0_io_rPort_11_ofs_0),
    .io_rPort_11_en_0(x258_lb_0_io_rPort_11_en_0),
    .io_rPort_11_backpressure(x258_lb_0_io_rPort_11_backpressure),
    .io_rPort_11_output_0(x258_lb_0_io_rPort_11_output_0),
    .io_rPort_10_banks_1(x258_lb_0_io_rPort_10_banks_1),
    .io_rPort_10_banks_0(x258_lb_0_io_rPort_10_banks_0),
    .io_rPort_10_ofs_0(x258_lb_0_io_rPort_10_ofs_0),
    .io_rPort_10_en_0(x258_lb_0_io_rPort_10_en_0),
    .io_rPort_10_backpressure(x258_lb_0_io_rPort_10_backpressure),
    .io_rPort_10_output_0(x258_lb_0_io_rPort_10_output_0),
    .io_rPort_9_banks_1(x258_lb_0_io_rPort_9_banks_1),
    .io_rPort_9_banks_0(x258_lb_0_io_rPort_9_banks_0),
    .io_rPort_9_ofs_0(x258_lb_0_io_rPort_9_ofs_0),
    .io_rPort_9_en_0(x258_lb_0_io_rPort_9_en_0),
    .io_rPort_9_backpressure(x258_lb_0_io_rPort_9_backpressure),
    .io_rPort_9_output_0(x258_lb_0_io_rPort_9_output_0),
    .io_rPort_8_banks_1(x258_lb_0_io_rPort_8_banks_1),
    .io_rPort_8_banks_0(x258_lb_0_io_rPort_8_banks_0),
    .io_rPort_8_ofs_0(x258_lb_0_io_rPort_8_ofs_0),
    .io_rPort_8_en_0(x258_lb_0_io_rPort_8_en_0),
    .io_rPort_8_backpressure(x258_lb_0_io_rPort_8_backpressure),
    .io_rPort_8_output_0(x258_lb_0_io_rPort_8_output_0),
    .io_rPort_7_banks_1(x258_lb_0_io_rPort_7_banks_1),
    .io_rPort_7_banks_0(x258_lb_0_io_rPort_7_banks_0),
    .io_rPort_7_ofs_0(x258_lb_0_io_rPort_7_ofs_0),
    .io_rPort_7_en_0(x258_lb_0_io_rPort_7_en_0),
    .io_rPort_7_backpressure(x258_lb_0_io_rPort_7_backpressure),
    .io_rPort_7_output_0(x258_lb_0_io_rPort_7_output_0),
    .io_rPort_6_banks_1(x258_lb_0_io_rPort_6_banks_1),
    .io_rPort_6_banks_0(x258_lb_0_io_rPort_6_banks_0),
    .io_rPort_6_ofs_0(x258_lb_0_io_rPort_6_ofs_0),
    .io_rPort_6_en_0(x258_lb_0_io_rPort_6_en_0),
    .io_rPort_6_backpressure(x258_lb_0_io_rPort_6_backpressure),
    .io_rPort_6_output_0(x258_lb_0_io_rPort_6_output_0),
    .io_rPort_5_banks_1(x258_lb_0_io_rPort_5_banks_1),
    .io_rPort_5_banks_0(x258_lb_0_io_rPort_5_banks_0),
    .io_rPort_5_ofs_0(x258_lb_0_io_rPort_5_ofs_0),
    .io_rPort_5_en_0(x258_lb_0_io_rPort_5_en_0),
    .io_rPort_5_backpressure(x258_lb_0_io_rPort_5_backpressure),
    .io_rPort_5_output_0(x258_lb_0_io_rPort_5_output_0),
    .io_rPort_4_banks_1(x258_lb_0_io_rPort_4_banks_1),
    .io_rPort_4_banks_0(x258_lb_0_io_rPort_4_banks_0),
    .io_rPort_4_ofs_0(x258_lb_0_io_rPort_4_ofs_0),
    .io_rPort_4_en_0(x258_lb_0_io_rPort_4_en_0),
    .io_rPort_4_backpressure(x258_lb_0_io_rPort_4_backpressure),
    .io_rPort_4_output_0(x258_lb_0_io_rPort_4_output_0),
    .io_rPort_3_banks_1(x258_lb_0_io_rPort_3_banks_1),
    .io_rPort_3_banks_0(x258_lb_0_io_rPort_3_banks_0),
    .io_rPort_3_ofs_0(x258_lb_0_io_rPort_3_ofs_0),
    .io_rPort_3_en_0(x258_lb_0_io_rPort_3_en_0),
    .io_rPort_3_backpressure(x258_lb_0_io_rPort_3_backpressure),
    .io_rPort_3_output_0(x258_lb_0_io_rPort_3_output_0),
    .io_rPort_2_banks_1(x258_lb_0_io_rPort_2_banks_1),
    .io_rPort_2_banks_0(x258_lb_0_io_rPort_2_banks_0),
    .io_rPort_2_ofs_0(x258_lb_0_io_rPort_2_ofs_0),
    .io_rPort_2_en_0(x258_lb_0_io_rPort_2_en_0),
    .io_rPort_2_backpressure(x258_lb_0_io_rPort_2_backpressure),
    .io_rPort_2_output_0(x258_lb_0_io_rPort_2_output_0),
    .io_rPort_1_banks_1(x258_lb_0_io_rPort_1_banks_1),
    .io_rPort_1_banks_0(x258_lb_0_io_rPort_1_banks_0),
    .io_rPort_1_ofs_0(x258_lb_0_io_rPort_1_ofs_0),
    .io_rPort_1_en_0(x258_lb_0_io_rPort_1_en_0),
    .io_rPort_1_backpressure(x258_lb_0_io_rPort_1_backpressure),
    .io_rPort_1_output_0(x258_lb_0_io_rPort_1_output_0),
    .io_rPort_0_banks_1(x258_lb_0_io_rPort_0_banks_1),
    .io_rPort_0_banks_0(x258_lb_0_io_rPort_0_banks_0),
    .io_rPort_0_ofs_0(x258_lb_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x258_lb_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x258_lb_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x258_lb_0_io_rPort_0_output_0),
    .io_wPort_1_banks_1(x258_lb_0_io_wPort_1_banks_1),
    .io_wPort_1_banks_0(x258_lb_0_io_wPort_1_banks_0),
    .io_wPort_1_ofs_0(x258_lb_0_io_wPort_1_ofs_0),
    .io_wPort_1_data_0(x258_lb_0_io_wPort_1_data_0),
    .io_wPort_1_en_0(x258_lb_0_io_wPort_1_en_0),
    .io_wPort_0_banks_1(x258_lb_0_io_wPort_0_banks_1),
    .io_wPort_0_banks_0(x258_lb_0_io_wPort_0_banks_0),
    .io_wPort_0_ofs_0(x258_lb_0_io_wPort_0_ofs_0),
    .io_wPort_0_data_0(x258_lb_0_io_wPort_0_data_0),
    .io_wPort_0_en_0(x258_lb_0_io_wPort_0_en_0)
  );
  x452_sub x464_sub_1 ( // @[Math.scala 191:24:@25607.4]
    .clock(x464_sub_1_clock),
    .reset(x464_sub_1_reset),
    .io_a(x464_sub_1_io_a),
    .io_b(x464_sub_1_io_b),
    .io_flow(x464_sub_1_io_flow),
    .io_result(x464_sub_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_1 ( // @[package.scala 93:22:@25634.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x235_sum x267_sum_1 ( // @[Math.scala 150:24:@25643.4]
    .clock(x267_sum_1_clock),
    .reset(x267_sum_1_reset),
    .io_a(x267_sum_1_io_a),
    .io_b(x267_sum_1_io_b),
    .io_flow(x267_sum_1_io_flow),
    .io_result(x267_sum_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_2 ( // @[package.scala 93:22:@25653.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_3 ( // @[package.scala 93:22:@25662.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper_168 RetimeWrapper_4 ( // @[package.scala 93:22:@25671.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_5 ( // @[package.scala 93:22:@25680.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper_172 RetimeWrapper_6 ( // @[package.scala 93:22:@25689.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper_172 RetimeWrapper_7 ( // @[package.scala 93:22:@25698.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper_172 RetimeWrapper_8 ( // @[package.scala 93:22:@25709.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  x235_sum x269_rdcol_1 ( // @[Math.scala 150:24:@25732.4]
    .clock(x269_rdcol_1_clock),
    .reset(x269_rdcol_1_reset),
    .io_a(x269_rdcol_1_io_a),
    .io_b(x269_rdcol_1_io_b),
    .io_flow(x269_rdcol_1_io_flow),
    .io_result(x269_rdcol_1_io_result)
  );
  x235_sum x273_sum_1 ( // @[Math.scala 150:24:@25772.4]
    .clock(x273_sum_1_clock),
    .reset(x273_sum_1_reset),
    .io_a(x273_sum_1_io_a),
    .io_b(x273_sum_1_io_b),
    .io_flow(x273_sum_1_io_flow),
    .io_result(x273_sum_1_io_result)
  );
  RetimeWrapper_169 RetimeWrapper_9 ( // @[package.scala 93:22:@25782.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_10 ( // @[package.scala 93:22:@25791.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_11 ( // @[package.scala 93:22:@25800.4]
    .clock(RetimeWrapper_11_clock),
    .reset(RetimeWrapper_11_reset),
    .io_flow(RetimeWrapper_11_io_flow),
    .io_in(RetimeWrapper_11_io_in),
    .io_out(RetimeWrapper_11_io_out)
  );
  RetimeWrapper_172 RetimeWrapper_12 ( // @[package.scala 93:22:@25811.4]
    .clock(RetimeWrapper_12_clock),
    .reset(RetimeWrapper_12_reset),
    .io_flow(RetimeWrapper_12_io_flow),
    .io_in(RetimeWrapper_12_io_in),
    .io_out(RetimeWrapper_12_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_13 ( // @[package.scala 93:22:@25832.4]
    .clock(RetimeWrapper_13_clock),
    .reset(RetimeWrapper_13_reset),
    .io_flow(RetimeWrapper_13_io_flow),
    .io_in(RetimeWrapper_13_io_in),
    .io_out(RetimeWrapper_13_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_14 ( // @[package.scala 93:22:@25848.4]
    .clock(RetimeWrapper_14_clock),
    .reset(RetimeWrapper_14_reset),
    .io_flow(RetimeWrapper_14_io_flow),
    .io_in(RetimeWrapper_14_io_in),
    .io_out(RetimeWrapper_14_io_out)
  );
  RetimeWrapper RetimeWrapper_15 ( // @[package.scala 93:22:@25864.4]
    .clock(RetimeWrapper_15_clock),
    .reset(RetimeWrapper_15_reset),
    .io_flow(RetimeWrapper_15_io_flow),
    .io_in(RetimeWrapper_15_io_in),
    .io_out(RetimeWrapper_15_io_out)
  );
  RetimeWrapper_184 RetimeWrapper_16 ( // @[package.scala 93:22:@25879.4]
    .clock(RetimeWrapper_16_clock),
    .reset(RetimeWrapper_16_reset),
    .io_flow(RetimeWrapper_16_io_flow),
    .io_in(RetimeWrapper_16_io_in),
    .io_out(RetimeWrapper_16_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_17 ( // @[package.scala 93:22:@25888.4]
    .clock(RetimeWrapper_17_clock),
    .reset(RetimeWrapper_17_reset),
    .io_flow(RetimeWrapper_17_io_flow),
    .io_in(RetimeWrapper_17_io_in),
    .io_out(RetimeWrapper_17_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_18 ( // @[package.scala 93:22:@25897.4]
    .clock(RetimeWrapper_18_clock),
    .reset(RetimeWrapper_18_reset),
    .io_flow(RetimeWrapper_18_io_flow),
    .io_in(RetimeWrapper_18_io_in),
    .io_out(RetimeWrapper_18_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_19 ( // @[package.scala 93:22:@25906.4]
    .clock(RetimeWrapper_19_clock),
    .reset(RetimeWrapper_19_reset),
    .io_flow(RetimeWrapper_19_io_flow),
    .io_in(RetimeWrapper_19_io_in),
    .io_out(RetimeWrapper_19_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_20 ( // @[package.scala 93:22:@25915.4]
    .clock(RetimeWrapper_20_clock),
    .reset(RetimeWrapper_20_reset),
    .io_flow(RetimeWrapper_20_io_flow),
    .io_in(RetimeWrapper_20_io_in),
    .io_out(RetimeWrapper_20_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_21 ( // @[package.scala 93:22:@25924.4]
    .clock(RetimeWrapper_21_clock),
    .reset(RetimeWrapper_21_reset),
    .io_flow(RetimeWrapper_21_io_flow),
    .io_in(RetimeWrapper_21_io_in),
    .io_out(RetimeWrapper_21_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_22 ( // @[package.scala 93:22:@25936.4]
    .clock(RetimeWrapper_22_clock),
    .reset(RetimeWrapper_22_reset),
    .io_flow(RetimeWrapper_22_io_flow),
    .io_in(RetimeWrapper_22_io_in),
    .io_out(RetimeWrapper_22_io_out)
  );
  RetimeWrapper_181 RetimeWrapper_23 ( // @[package.scala 93:22:@25957.4]
    .clock(RetimeWrapper_23_clock),
    .reset(RetimeWrapper_23_reset),
    .io_flow(RetimeWrapper_23_io_flow),
    .io_in(RetimeWrapper_23_io_in),
    .io_out(RetimeWrapper_23_io_out)
  );
  RetimeWrapper_172 RetimeWrapper_24 ( // @[package.scala 93:22:@25981.4]
    .clock(RetimeWrapper_24_clock),
    .reset(RetimeWrapper_24_reset),
    .io_flow(RetimeWrapper_24_io_flow),
    .io_in(RetimeWrapper_24_io_in),
    .io_out(RetimeWrapper_24_io_out)
  );
  RetimeWrapper_184 RetimeWrapper_25 ( // @[package.scala 93:22:@25990.4]
    .clock(RetimeWrapper_25_clock),
    .reset(RetimeWrapper_25_reset),
    .io_flow(RetimeWrapper_25_io_flow),
    .io_in(RetimeWrapper_25_io_in),
    .io_out(RetimeWrapper_25_io_out)
  );
  RetimeWrapper_188 RetimeWrapper_26 ( // @[package.scala 93:22:@25999.4]
    .clock(RetimeWrapper_26_clock),
    .reset(RetimeWrapper_26_reset),
    .io_flow(RetimeWrapper_26_io_flow),
    .io_in(RetimeWrapper_26_io_in),
    .io_out(RetimeWrapper_26_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_27 ( // @[package.scala 93:22:@26011.4]
    .clock(RetimeWrapper_27_clock),
    .reset(RetimeWrapper_27_reset),
    .io_flow(RetimeWrapper_27_io_flow),
    .io_in(RetimeWrapper_27_io_in),
    .io_out(RetimeWrapper_27_io_out)
  );
  x235_sum x287_rdcol_1 ( // @[Math.scala 150:24:@26034.4]
    .clock(x287_rdcol_1_clock),
    .reset(x287_rdcol_1_reset),
    .io_a(x287_rdcol_1_io_a),
    .io_b(x287_rdcol_1_io_b),
    .io_flow(x287_rdcol_1_io_flow),
    .io_result(x287_rdcol_1_io_result)
  );
  RetimeWrapper_181 RetimeWrapper_28 ( // @[package.scala 93:22:@26085.4]
    .clock(RetimeWrapper_28_clock),
    .reset(RetimeWrapper_28_reset),
    .io_flow(RetimeWrapper_28_io_flow),
    .io_in(RetimeWrapper_28_io_in),
    .io_out(RetimeWrapper_28_io_out)
  );
  x235_sum x293_sum_1 ( // @[Math.scala 150:24:@26094.4]
    .clock(x293_sum_1_clock),
    .reset(x293_sum_1_reset),
    .io_a(x293_sum_1_io_a),
    .io_b(x293_sum_1_io_b),
    .io_flow(x293_sum_1_io_flow),
    .io_result(x293_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_29 ( // @[package.scala 93:22:@26104.4]
    .clock(RetimeWrapper_29_clock),
    .reset(RetimeWrapper_29_reset),
    .io_flow(RetimeWrapper_29_io_flow),
    .io_in(RetimeWrapper_29_io_in),
    .io_out(RetimeWrapper_29_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_30 ( // @[package.scala 93:22:@26113.4]
    .clock(RetimeWrapper_30_clock),
    .reset(RetimeWrapper_30_reset),
    .io_flow(RetimeWrapper_30_io_flow),
    .io_in(RetimeWrapper_30_io_in),
    .io_out(RetimeWrapper_30_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_31 ( // @[package.scala 93:22:@26122.4]
    .clock(RetimeWrapper_31_clock),
    .reset(RetimeWrapper_31_reset),
    .io_flow(RetimeWrapper_31_io_flow),
    .io_in(RetimeWrapper_31_io_in),
    .io_out(RetimeWrapper_31_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_32 ( // @[package.scala 93:22:@26134.4]
    .clock(RetimeWrapper_32_clock),
    .reset(RetimeWrapper_32_reset),
    .io_flow(RetimeWrapper_32_io_flow),
    .io_in(RetimeWrapper_32_io_in),
    .io_out(RetimeWrapper_32_io_out)
  );
  x235_sum x296_rdcol_1 ( // @[Math.scala 150:24:@26157.4]
    .clock(x296_rdcol_1_clock),
    .reset(x296_rdcol_1_reset),
    .io_a(x296_rdcol_1_io_a),
    .io_b(x296_rdcol_1_io_b),
    .io_flow(x296_rdcol_1_io_flow),
    .io_result(x296_rdcol_1_io_result)
  );
  x235_sum x302_sum_1 ( // @[Math.scala 150:24:@26208.4]
    .clock(x302_sum_1_clock),
    .reset(x302_sum_1_reset),
    .io_a(x302_sum_1_io_a),
    .io_b(x302_sum_1_io_b),
    .io_flow(x302_sum_1_io_flow),
    .io_result(x302_sum_1_io_result)
  );
  RetimeWrapper_29 RetimeWrapper_33 ( // @[package.scala 93:22:@26218.4]
    .clock(RetimeWrapper_33_clock),
    .reset(RetimeWrapper_33_reset),
    .io_flow(RetimeWrapper_33_io_flow),
    .io_in(RetimeWrapper_33_io_in),
    .io_out(RetimeWrapper_33_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_34 ( // @[package.scala 93:22:@26227.4]
    .clock(RetimeWrapper_34_clock),
    .reset(RetimeWrapper_34_reset),
    .io_flow(RetimeWrapper_34_io_flow),
    .io_in(RetimeWrapper_34_io_in),
    .io_out(RetimeWrapper_34_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_35 ( // @[package.scala 93:22:@26236.4]
    .clock(RetimeWrapper_35_clock),
    .reset(RetimeWrapper_35_reset),
    .io_flow(RetimeWrapper_35_io_flow),
    .io_in(RetimeWrapper_35_io_in),
    .io_out(RetimeWrapper_35_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_36 ( // @[package.scala 93:22:@26248.4]
    .clock(RetimeWrapper_36_clock),
    .reset(RetimeWrapper_36_reset),
    .io_flow(RetimeWrapper_36_io_flow),
    .io_in(RetimeWrapper_36_io_in),
    .io_out(RetimeWrapper_36_io_out)
  );
  x452_sub x305_rdrow_1 ( // @[Math.scala 191:24:@26271.4]
    .clock(x305_rdrow_1_clock),
    .reset(x305_rdrow_1_reset),
    .io_a(x305_rdrow_1_io_a),
    .io_b(x305_rdrow_1_io_b),
    .io_flow(x305_rdrow_1_io_flow),
    .io_result(x305_rdrow_1_io_result)
  );
  x452_sub x472_sub_1 ( // @[Math.scala 191:24:@26343.4]
    .clock(x472_sub_1_clock),
    .reset(x472_sub_1_reset),
    .io_a(x472_sub_1_io_a),
    .io_b(x472_sub_1_io_b),
    .io_flow(x472_sub_1_io_flow),
    .io_result(x472_sub_1_io_result)
  );
  RetimeWrapper_188 RetimeWrapper_37 ( // @[package.scala 93:22:@26353.4]
    .clock(RetimeWrapper_37_clock),
    .reset(RetimeWrapper_37_reset),
    .io_flow(RetimeWrapper_37_io_flow),
    .io_in(RetimeWrapper_37_io_in),
    .io_out(RetimeWrapper_37_io_out)
  );
  x235_sum x313_sum_1 ( // @[Math.scala 150:24:@26362.4]
    .clock(x313_sum_1_clock),
    .reset(x313_sum_1_reset),
    .io_a(x313_sum_1_io_a),
    .io_b(x313_sum_1_io_b),
    .io_flow(x313_sum_1_io_flow),
    .io_result(x313_sum_1_io_result)
  );
  RetimeWrapper_169 RetimeWrapper_38 ( // @[package.scala 93:22:@26372.4]
    .clock(RetimeWrapper_38_clock),
    .reset(RetimeWrapper_38_reset),
    .io_flow(RetimeWrapper_38_io_flow),
    .io_in(RetimeWrapper_38_io_in),
    .io_out(RetimeWrapper_38_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_39 ( // @[package.scala 93:22:@26381.4]
    .clock(RetimeWrapper_39_clock),
    .reset(RetimeWrapper_39_reset),
    .io_flow(RetimeWrapper_39_io_flow),
    .io_in(RetimeWrapper_39_io_in),
    .io_out(RetimeWrapper_39_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_40 ( // @[package.scala 93:22:@26393.4]
    .clock(RetimeWrapper_40_clock),
    .reset(RetimeWrapper_40_reset),
    .io_flow(RetimeWrapper_40_io_flow),
    .io_in(RetimeWrapper_40_io_in),
    .io_out(RetimeWrapper_40_io_out)
  );
  RetimeWrapper RetimeWrapper_41 ( // @[package.scala 93:22:@26414.4]
    .clock(RetimeWrapper_41_clock),
    .reset(RetimeWrapper_41_reset),
    .io_flow(RetimeWrapper_41_io_flow),
    .io_in(RetimeWrapper_41_io_in),
    .io_out(RetimeWrapper_41_io_out)
  );
  RetimeWrapper_187 RetimeWrapper_42 ( // @[package.scala 93:22:@26429.4]
    .clock(RetimeWrapper_42_clock),
    .reset(RetimeWrapper_42_reset),
    .io_flow(RetimeWrapper_42_io_flow),
    .io_in(RetimeWrapper_42_io_in),
    .io_out(RetimeWrapper_42_io_out)
  );
  x235_sum x318_sum_1 ( // @[Math.scala 150:24:@26440.4]
    .clock(x318_sum_1_clock),
    .reset(x318_sum_1_reset),
    .io_a(x318_sum_1_io_a),
    .io_b(x318_sum_1_io_b),
    .io_flow(x318_sum_1_io_flow),
    .io_result(x318_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_43 ( // @[package.scala 93:22:@26450.4]
    .clock(RetimeWrapper_43_clock),
    .reset(RetimeWrapper_43_reset),
    .io_flow(RetimeWrapper_43_io_flow),
    .io_in(RetimeWrapper_43_io_in),
    .io_out(RetimeWrapper_43_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_44 ( // @[package.scala 93:22:@26462.4]
    .clock(RetimeWrapper_44_clock),
    .reset(RetimeWrapper_44_reset),
    .io_flow(RetimeWrapper_44_io_flow),
    .io_in(RetimeWrapper_44_io_in),
    .io_out(RetimeWrapper_44_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_45 ( // @[package.scala 93:22:@26489.4]
    .clock(RetimeWrapper_45_clock),
    .reset(RetimeWrapper_45_reset),
    .io_flow(RetimeWrapper_45_io_flow),
    .io_in(RetimeWrapper_45_io_in),
    .io_out(RetimeWrapper_45_io_out)
  );
  x235_sum x323_sum_1 ( // @[Math.scala 150:24:@26498.4]
    .clock(x323_sum_1_clock),
    .reset(x323_sum_1_reset),
    .io_a(x323_sum_1_io_a),
    .io_b(x323_sum_1_io_b),
    .io_flow(x323_sum_1_io_flow),
    .io_result(x323_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_46 ( // @[package.scala 93:22:@26508.4]
    .clock(RetimeWrapper_46_clock),
    .reset(RetimeWrapper_46_reset),
    .io_flow(RetimeWrapper_46_io_flow),
    .io_in(RetimeWrapper_46_io_in),
    .io_out(RetimeWrapper_46_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_47 ( // @[package.scala 93:22:@26520.4]
    .clock(RetimeWrapper_47_clock),
    .reset(RetimeWrapper_47_reset),
    .io_flow(RetimeWrapper_47_io_flow),
    .io_in(RetimeWrapper_47_io_in),
    .io_out(RetimeWrapper_47_io_out)
  );
  RetimeWrapper_29 RetimeWrapper_48 ( // @[package.scala 93:22:@26547.4]
    .clock(RetimeWrapper_48_clock),
    .reset(RetimeWrapper_48_reset),
    .io_flow(RetimeWrapper_48_io_flow),
    .io_in(RetimeWrapper_48_io_in),
    .io_out(RetimeWrapper_48_io_out)
  );
  x235_sum x328_sum_1 ( // @[Math.scala 150:24:@26556.4]
    .clock(x328_sum_1_clock),
    .reset(x328_sum_1_reset),
    .io_a(x328_sum_1_io_a),
    .io_b(x328_sum_1_io_b),
    .io_flow(x328_sum_1_io_flow),
    .io_result(x328_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_49 ( // @[package.scala 93:22:@26566.4]
    .clock(RetimeWrapper_49_clock),
    .reset(RetimeWrapper_49_reset),
    .io_flow(RetimeWrapper_49_io_flow),
    .io_in(RetimeWrapper_49_io_in),
    .io_out(RetimeWrapper_49_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_50 ( // @[package.scala 93:22:@26578.4]
    .clock(RetimeWrapper_50_clock),
    .reset(RetimeWrapper_50_reset),
    .io_flow(RetimeWrapper_50_io_flow),
    .io_in(RetimeWrapper_50_io_in),
    .io_out(RetimeWrapper_50_io_out)
  );
  x452_sub x331_rdrow_1 ( // @[Math.scala 191:24:@26601.4]
    .clock(x331_rdrow_1_clock),
    .reset(x331_rdrow_1_reset),
    .io_a(x331_rdrow_1_io_a),
    .io_b(x331_rdrow_1_io_b),
    .io_flow(x331_rdrow_1_io_flow),
    .io_result(x331_rdrow_1_io_result)
  );
  x452_sub x477_sub_1 ( // @[Math.scala 191:24:@26673.4]
    .clock(x477_sub_1_clock),
    .reset(x477_sub_1_reset),
    .io_a(x477_sub_1_io_a),
    .io_b(x477_sub_1_io_b),
    .io_flow(x477_sub_1_io_flow),
    .io_result(x477_sub_1_io_result)
  );
  x235_sum x339_sum_1 ( // @[Math.scala 150:24:@26683.4]
    .clock(x339_sum_1_clock),
    .reset(x339_sum_1_reset),
    .io_a(x339_sum_1_io_a),
    .io_b(x339_sum_1_io_b),
    .io_flow(x339_sum_1_io_flow),
    .io_result(x339_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_51 ( // @[package.scala 93:22:@26693.4]
    .clock(RetimeWrapper_51_clock),
    .reset(RetimeWrapper_51_reset),
    .io_flow(RetimeWrapper_51_io_flow),
    .io_in(RetimeWrapper_51_io_in),
    .io_out(RetimeWrapper_51_io_out)
  );
  RetimeWrapper_169 RetimeWrapper_52 ( // @[package.scala 93:22:@26702.4]
    .clock(RetimeWrapper_52_clock),
    .reset(RetimeWrapper_52_reset),
    .io_flow(RetimeWrapper_52_io_flow),
    .io_in(RetimeWrapper_52_io_in),
    .io_out(RetimeWrapper_52_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_53 ( // @[package.scala 93:22:@26714.4]
    .clock(RetimeWrapper_53_clock),
    .reset(RetimeWrapper_53_reset),
    .io_flow(RetimeWrapper_53_io_flow),
    .io_in(RetimeWrapper_53_io_in),
    .io_out(RetimeWrapper_53_io_out)
  );
  x235_sum x344_sum_1 ( // @[Math.scala 150:24:@26741.4]
    .clock(x344_sum_1_clock),
    .reset(x344_sum_1_reset),
    .io_a(x344_sum_1_io_a),
    .io_b(x344_sum_1_io_b),
    .io_flow(x344_sum_1_io_flow),
    .io_result(x344_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_54 ( // @[package.scala 93:22:@26751.4]
    .clock(RetimeWrapper_54_clock),
    .reset(RetimeWrapper_54_reset),
    .io_flow(RetimeWrapper_54_io_flow),
    .io_in(RetimeWrapper_54_io_in),
    .io_out(RetimeWrapper_54_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_55 ( // @[package.scala 93:22:@26763.4]
    .clock(RetimeWrapper_55_clock),
    .reset(RetimeWrapper_55_reset),
    .io_flow(RetimeWrapper_55_io_flow),
    .io_in(RetimeWrapper_55_io_in),
    .io_out(RetimeWrapper_55_io_out)
  );
  x235_sum x349_sum_1 ( // @[Math.scala 150:24:@26790.4]
    .clock(x349_sum_1_clock),
    .reset(x349_sum_1_reset),
    .io_a(x349_sum_1_io_a),
    .io_b(x349_sum_1_io_b),
    .io_flow(x349_sum_1_io_flow),
    .io_result(x349_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_56 ( // @[package.scala 93:22:@26800.4]
    .clock(RetimeWrapper_56_clock),
    .reset(RetimeWrapper_56_reset),
    .io_flow(RetimeWrapper_56_io_flow),
    .io_in(RetimeWrapper_56_io_in),
    .io_out(RetimeWrapper_56_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_57 ( // @[package.scala 93:22:@26812.4]
    .clock(RetimeWrapper_57_clock),
    .reset(RetimeWrapper_57_reset),
    .io_flow(RetimeWrapper_57_io_flow),
    .io_in(RetimeWrapper_57_io_in),
    .io_out(RetimeWrapper_57_io_out)
  );
  x235_sum x354_sum_1 ( // @[Math.scala 150:24:@26841.4]
    .clock(x354_sum_1_clock),
    .reset(x354_sum_1_reset),
    .io_a(x354_sum_1_io_a),
    .io_b(x354_sum_1_io_b),
    .io_flow(x354_sum_1_io_flow),
    .io_result(x354_sum_1_io_result)
  );
  RetimeWrapper_6 RetimeWrapper_58 ( // @[package.scala 93:22:@26851.4]
    .clock(RetimeWrapper_58_clock),
    .reset(RetimeWrapper_58_reset),
    .io_flow(RetimeWrapper_58_io_flow),
    .io_in(RetimeWrapper_58_io_in),
    .io_out(RetimeWrapper_58_io_out)
  );
  RetimeWrapper_186 RetimeWrapper_59 ( // @[package.scala 93:22:@26863.4]
    .clock(RetimeWrapper_59_clock),
    .reset(RetimeWrapper_59_reset),
    .io_flow(RetimeWrapper_59_io_flow),
    .io_in(RetimeWrapper_59_io_in),
    .io_out(RetimeWrapper_59_io_out)
  );
  x357 x357_1 ( // @[Math.scala 262:24:@26886.4]
    .clock(x357_1_clock),
    .io_a(x357_1_io_a),
    .io_b(x357_1_io_b),
    .io_flow(x357_1_io_flow),
    .io_result(x357_1_io_result)
  );
  x357 x358_1 ( // @[Math.scala 262:24:@26898.4]
    .clock(x358_1_clock),
    .io_a(x358_1_io_a),
    .io_b(x358_1_io_b),
    .io_flow(x358_1_io_flow),
    .io_result(x358_1_io_result)
  );
  x357 x359_1 ( // @[Math.scala 262:24:@26910.4]
    .clock(x359_1_clock),
    .io_a(x359_1_io_a),
    .io_b(x359_1_io_b),
    .io_flow(x359_1_io_flow),
    .io_result(x359_1_io_result)
  );
  x357 x360_1 ( // @[Math.scala 262:24:@26922.4]
    .clock(x360_1_clock),
    .io_a(x360_1_io_a),
    .io_b(x360_1_io_b),
    .io_flow(x360_1_io_flow),
    .io_result(x360_1_io_result)
  );
  x357 x361_1 ( // @[Math.scala 262:24:@26934.4]
    .clock(x361_1_clock),
    .io_a(x361_1_io_a),
    .io_b(x361_1_io_b),
    .io_flow(x361_1_io_flow),
    .io_result(x361_1_io_result)
  );
  x357 x362_1 ( // @[Math.scala 262:24:@26946.4]
    .clock(x362_1_clock),
    .io_a(x362_1_io_a),
    .io_b(x362_1_io_b),
    .io_flow(x362_1_io_flow),
    .io_result(x362_1_io_result)
  );
  x357 x363_1 ( // @[Math.scala 262:24:@26958.4]
    .clock(x363_1_clock),
    .io_a(x363_1_io_a),
    .io_b(x363_1_io_b),
    .io_flow(x363_1_io_flow),
    .io_result(x363_1_io_result)
  );
  x357 x364_1 ( // @[Math.scala 262:24:@26970.4]
    .clock(x364_1_clock),
    .io_a(x364_1_io_a),
    .io_b(x364_1_io_b),
    .io_flow(x364_1_io_flow),
    .io_result(x364_1_io_result)
  );
  x357 x365_1 ( // @[Math.scala 262:24:@26982.4]
    .clock(x365_1_clock),
    .io_a(x365_1_io_a),
    .io_b(x365_1_io_b),
    .io_flow(x365_1_io_flow),
    .io_result(x365_1_io_result)
  );
  x366_x3 x366_x3_1 ( // @[Math.scala 150:24:@26992.4]
    .clock(x366_x3_1_clock),
    .reset(x366_x3_1_reset),
    .io_a(x366_x3_1_io_a),
    .io_b(x366_x3_1_io_b),
    .io_flow(x366_x3_1_io_flow),
    .io_result(x366_x3_1_io_result)
  );
  x366_x3 x367_x4_1 ( // @[Math.scala 150:24:@27002.4]
    .clock(x367_x4_1_clock),
    .reset(x367_x4_1_reset),
    .io_a(x367_x4_1_io_a),
    .io_b(x367_x4_1_io_b),
    .io_flow(x367_x4_1_io_flow),
    .io_result(x367_x4_1_io_result)
  );
  x366_x3 x368_x3_1 ( // @[Math.scala 150:24:@27012.4]
    .clock(x368_x3_1_clock),
    .reset(x368_x3_1_reset),
    .io_a(x368_x3_1_io_a),
    .io_b(x368_x3_1_io_b),
    .io_flow(x368_x3_1_io_flow),
    .io_result(x368_x3_1_io_result)
  );
  x366_x3 x369_x4_1 ( // @[Math.scala 150:24:@27022.4]
    .clock(x369_x4_1_clock),
    .reset(x369_x4_1_reset),
    .io_a(x369_x4_1_io_a),
    .io_b(x369_x4_1_io_b),
    .io_flow(x369_x4_1_io_flow),
    .io_result(x369_x4_1_io_result)
  );
  x366_x3 x370_x3_1 ( // @[Math.scala 150:24:@27032.4]
    .clock(x370_x3_1_clock),
    .reset(x370_x3_1_reset),
    .io_a(x370_x3_1_io_a),
    .io_b(x370_x3_1_io_b),
    .io_flow(x370_x3_1_io_flow),
    .io_result(x370_x3_1_io_result)
  );
  x366_x3 x371_x4_1 ( // @[Math.scala 150:24:@27042.4]
    .clock(x371_x4_1_clock),
    .reset(x371_x4_1_reset),
    .io_a(x371_x4_1_io_a),
    .io_b(x371_x4_1_io_b),
    .io_flow(x371_x4_1_io_flow),
    .io_result(x371_x4_1_io_result)
  );
  x366_x3 x372_x3_1 ( // @[Math.scala 150:24:@27052.4]
    .clock(x372_x3_1_clock),
    .reset(x372_x3_1_reset),
    .io_a(x372_x3_1_io_a),
    .io_b(x372_x3_1_io_b),
    .io_flow(x372_x3_1_io_flow),
    .io_result(x372_x3_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_60 ( // @[package.scala 93:22:@27062.4]
    .clock(RetimeWrapper_60_clock),
    .reset(RetimeWrapper_60_reset),
    .io_flow(RetimeWrapper_60_io_flow),
    .io_in(RetimeWrapper_60_io_in),
    .io_out(RetimeWrapper_60_io_out)
  );
  x366_x3 x373_sum_1 ( // @[Math.scala 150:24:@27071.4]
    .clock(x373_sum_1_clock),
    .reset(x373_sum_1_reset),
    .io_a(x373_sum_1_io_a),
    .io_b(x373_sum_1_io_b),
    .io_flow(x373_sum_1_io_flow),
    .io_result(x373_sum_1_io_result)
  );
  x374 x374_1 ( // @[Math.scala 720:24:@27081.4]
    .io_b(x374_1_io_b),
    .io_result(x374_1_io_result)
  );
  x375_mul x375_mul_1 ( // @[Math.scala 262:24:@27092.4]
    .clock(x375_mul_1_clock),
    .io_a(x375_mul_1_io_a),
    .io_flow(x375_mul_1_io_flow),
    .io_result(x375_mul_1_io_result)
  );
  x376 x376_1 ( // @[Math.scala 720:24:@27102.4]
    .io_b(x376_1_io_b),
    .io_result(x376_1_io_result)
  );
  x357 x377_1 ( // @[Math.scala 262:24:@27113.4]
    .clock(x377_1_clock),
    .io_a(x377_1_io_a),
    .io_b(x377_1_io_b),
    .io_flow(x377_1_io_flow),
    .io_result(x377_1_io_result)
  );
  x357 x378_1 ( // @[Math.scala 262:24:@27125.4]
    .clock(x378_1_clock),
    .io_a(x378_1_io_a),
    .io_b(x378_1_io_b),
    .io_flow(x378_1_io_flow),
    .io_result(x378_1_io_result)
  );
  x357 x379_1 ( // @[Math.scala 262:24:@27137.4]
    .clock(x379_1_clock),
    .io_a(x379_1_io_a),
    .io_b(x379_1_io_b),
    .io_flow(x379_1_io_flow),
    .io_result(x379_1_io_result)
  );
  x357 x380_1 ( // @[Math.scala 262:24:@27149.4]
    .clock(x380_1_clock),
    .io_a(x380_1_io_a),
    .io_b(x380_1_io_b),
    .io_flow(x380_1_io_flow),
    .io_result(x380_1_io_result)
  );
  x357 x381_1 ( // @[Math.scala 262:24:@27161.4]
    .clock(x381_1_clock),
    .io_a(x381_1_io_a),
    .io_b(x381_1_io_b),
    .io_flow(x381_1_io_flow),
    .io_result(x381_1_io_result)
  );
  x357 x382_1 ( // @[Math.scala 262:24:@27173.4]
    .clock(x382_1_clock),
    .io_a(x382_1_io_a),
    .io_b(x382_1_io_b),
    .io_flow(x382_1_io_flow),
    .io_result(x382_1_io_result)
  );
  x357 x383_1 ( // @[Math.scala 262:24:@27185.4]
    .clock(x383_1_clock),
    .io_a(x383_1_io_a),
    .io_b(x383_1_io_b),
    .io_flow(x383_1_io_flow),
    .io_result(x383_1_io_result)
  );
  x357 x384_1 ( // @[Math.scala 262:24:@27197.4]
    .clock(x384_1_clock),
    .io_a(x384_1_io_a),
    .io_b(x384_1_io_b),
    .io_flow(x384_1_io_flow),
    .io_result(x384_1_io_result)
  );
  x357 x385_1 ( // @[Math.scala 262:24:@27209.4]
    .clock(x385_1_clock),
    .io_a(x385_1_io_a),
    .io_b(x385_1_io_b),
    .io_flow(x385_1_io_flow),
    .io_result(x385_1_io_result)
  );
  x366_x3 x386_x3_1 ( // @[Math.scala 150:24:@27219.4]
    .clock(x386_x3_1_clock),
    .reset(x386_x3_1_reset),
    .io_a(x386_x3_1_io_a),
    .io_b(x386_x3_1_io_b),
    .io_flow(x386_x3_1_io_flow),
    .io_result(x386_x3_1_io_result)
  );
  x366_x3 x387_x4_1 ( // @[Math.scala 150:24:@27229.4]
    .clock(x387_x4_1_clock),
    .reset(x387_x4_1_reset),
    .io_a(x387_x4_1_io_a),
    .io_b(x387_x4_1_io_b),
    .io_flow(x387_x4_1_io_flow),
    .io_result(x387_x4_1_io_result)
  );
  x366_x3 x388_x3_1 ( // @[Math.scala 150:24:@27239.4]
    .clock(x388_x3_1_clock),
    .reset(x388_x3_1_reset),
    .io_a(x388_x3_1_io_a),
    .io_b(x388_x3_1_io_b),
    .io_flow(x388_x3_1_io_flow),
    .io_result(x388_x3_1_io_result)
  );
  x366_x3 x389_x4_1 ( // @[Math.scala 150:24:@27249.4]
    .clock(x389_x4_1_clock),
    .reset(x389_x4_1_reset),
    .io_a(x389_x4_1_io_a),
    .io_b(x389_x4_1_io_b),
    .io_flow(x389_x4_1_io_flow),
    .io_result(x389_x4_1_io_result)
  );
  x366_x3 x390_x3_1 ( // @[Math.scala 150:24:@27259.4]
    .clock(x390_x3_1_clock),
    .reset(x390_x3_1_reset),
    .io_a(x390_x3_1_io_a),
    .io_b(x390_x3_1_io_b),
    .io_flow(x390_x3_1_io_flow),
    .io_result(x390_x3_1_io_result)
  );
  x366_x3 x391_x4_1 ( // @[Math.scala 150:24:@27269.4]
    .clock(x391_x4_1_clock),
    .reset(x391_x4_1_reset),
    .io_a(x391_x4_1_io_a),
    .io_b(x391_x4_1_io_b),
    .io_flow(x391_x4_1_io_flow),
    .io_result(x391_x4_1_io_result)
  );
  x366_x3 x392_x3_1 ( // @[Math.scala 150:24:@27279.4]
    .clock(x392_x3_1_clock),
    .reset(x392_x3_1_reset),
    .io_a(x392_x3_1_io_a),
    .io_b(x392_x3_1_io_b),
    .io_flow(x392_x3_1_io_flow),
    .io_result(x392_x3_1_io_result)
  );
  RetimeWrapper_168 RetimeWrapper_61 ( // @[package.scala 93:22:@27289.4]
    .clock(RetimeWrapper_61_clock),
    .reset(RetimeWrapper_61_reset),
    .io_flow(RetimeWrapper_61_io_flow),
    .io_in(RetimeWrapper_61_io_in),
    .io_out(RetimeWrapper_61_io_out)
  );
  x366_x3 x393_sum_1 ( // @[Math.scala 150:24:@27298.4]
    .clock(x393_sum_1_clock),
    .reset(x393_sum_1_reset),
    .io_a(x393_sum_1_io_a),
    .io_b(x393_sum_1_io_b),
    .io_flow(x393_sum_1_io_flow),
    .io_result(x393_sum_1_io_result)
  );
  x374 x394_1 ( // @[Math.scala 720:24:@27308.4]
    .io_b(x394_1_io_b),
    .io_result(x394_1_io_result)
  );
  x375_mul x395_mul_1 ( // @[Math.scala 262:24:@27319.4]
    .clock(x395_mul_1_clock),
    .io_a(x395_mul_1_io_a),
    .io_flow(x395_mul_1_io_flow),
    .io_result(x395_mul_1_io_result)
  );
  x376 x396_1 ( // @[Math.scala 720:24:@27329.4]
    .io_b(x396_1_io_b),
    .io_result(x396_1_io_result)
  );
  RetimeWrapper_262 RetimeWrapper_62 ( // @[package.scala 93:22:@27344.4]
    .clock(RetimeWrapper_62_clock),
    .reset(RetimeWrapper_62_reset),
    .io_flow(RetimeWrapper_62_io_flow),
    .io_in(RetimeWrapper_62_io_in),
    .io_out(RetimeWrapper_62_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_63 ( // @[package.scala 93:22:@27353.4]
    .clock(RetimeWrapper_63_clock),
    .reset(RetimeWrapper_63_reset),
    .io_flow(RetimeWrapper_63_io_flow),
    .io_in(RetimeWrapper_63_io_in),
    .io_out(RetimeWrapper_63_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_64 ( // @[package.scala 93:22:@27362.4]
    .clock(RetimeWrapper_64_clock),
    .reset(RetimeWrapper_64_reset),
    .io_flow(RetimeWrapper_64_io_flow),
    .io_in(RetimeWrapper_64_io_in),
    .io_out(RetimeWrapper_64_io_out)
  );
  RetimeWrapper_48 RetimeWrapper_65 ( // @[package.scala 93:22:@27371.4]
    .clock(RetimeWrapper_65_clock),
    .reset(RetimeWrapper_65_reset),
    .io_flow(RetimeWrapper_65_io_flow),
    .io_in(RetimeWrapper_65_io_in),
    .io_out(RetimeWrapper_65_io_out)
  );
  assign b254 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 62:18:@25419.4]
  assign b255 = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 63:18:@25420.4]
  assign _T_205 = b254 & b255; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 67:30:@25422.4]
  assign _T_206 = _T_205 & io_sigsIn_datapathEn; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 67:37:@25423.4]
  assign _T_210 = io_in_x221_TID == 8'h0; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 69:76:@25428.4]
  assign _T_211 = _T_206 & _T_210; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 69:62:@25429.4]
  assign _T_213 = io_in_x221_TDEST == 8'h0; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 69:101:@25430.4]
  assign x483_x256_D1_0_number = RetimeWrapper_io_out; // @[package.scala 96:25:@25439.4 package.scala 96:25:@25440.4]
  assign b252_number = __io_result; // @[Math.scala 723:22:@25404.4 Math.scala 724:14:@25405.4]
  assign _T_243 = $signed(b252_number); // @[Math.scala 406:49:@25548.4]
  assign _T_245 = $signed(_T_243) & $signed(32'sh3); // @[Math.scala 406:56:@25550.4]
  assign _T_246 = $signed(_T_245); // @[Math.scala 406:56:@25551.4]
  assign x459_number = $unsigned(_T_246); // @[implicits.scala 133:21:@25552.4]
  assign _T_256 = $signed(x459_number); // @[Math.scala 406:49:@25561.4]
  assign _T_258 = $signed(_T_256) & $signed(32'sh3); // @[Math.scala 406:56:@25563.4]
  assign _T_259 = $signed(_T_258); // @[Math.scala 406:56:@25564.4]
  assign b253_number = __1_io_result; // @[Math.scala 723:22:@25416.4 Math.scala 724:14:@25417.4]
  assign _T_268 = $signed(b253_number); // @[Math.scala 406:49:@25572.4]
  assign _T_270 = $signed(_T_268) & $signed(32'sh3); // @[Math.scala 406:56:@25574.4]
  assign _T_271 = $signed(_T_270); // @[Math.scala 406:56:@25575.4]
  assign _T_275 = x459_number[31]; // @[FixedPoint.scala 50:25:@25581.4]
  assign _T_279 = _T_275 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25583.4]
  assign _T_280 = x459_number[31:2]; // @[FixedPoint.scala 18:52:@25584.4]
  assign _T_286 = _T_280 == 30'h3fffffff; // @[Math.scala 451:55:@25586.4]
  assign _T_287 = x459_number[1:0]; // @[FixedPoint.scala 18:52:@25587.4]
  assign _T_293 = _T_287 != 2'h0; // @[Math.scala 451:110:@25589.4]
  assign _T_294 = _T_286 & _T_293; // @[Math.scala 451:94:@25590.4]
  assign _T_296 = {_T_279,_T_280}; // @[Cat.scala 30:58:@25592.4]
  assign x264_1_number = _T_294 ? 32'h0 : _T_296; // @[Math.scala 454:20:@25593.4]
  assign _GEN_0 = {{9'd0}, x264_1_number}; // @[Math.scala 461:32:@25598.4]
  assign _T_301 = _GEN_0 << 9; // @[Math.scala 461:32:@25598.4]
  assign _GEN_1 = {{5'd0}, x264_1_number}; // @[Math.scala 461:32:@25603.4]
  assign _T_304 = _GEN_1 << 5; // @[Math.scala 461:32:@25603.4]
  assign _T_310 = b253_number[31]; // @[FixedPoint.scala 50:25:@25618.4]
  assign _T_314 = _T_310 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25620.4]
  assign _T_315 = b253_number[31:2]; // @[FixedPoint.scala 18:52:@25621.4]
  assign _T_321 = _T_315 == 30'h3fffffff; // @[Math.scala 451:55:@25623.4]
  assign _T_322 = b253_number[1:0]; // @[FixedPoint.scala 18:52:@25624.4]
  assign _T_328 = _T_322 != 2'h0; // @[Math.scala 451:110:@25626.4]
  assign _T_329 = _T_321 & _T_328; // @[Math.scala 451:94:@25627.4]
  assign _T_331 = {_T_314,_T_315}; // @[Cat.scala 30:58:@25629.4]
  assign _T_359 = ~ io_sigsIn_break; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:101:@25706.4]
  assign _T_363 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@25714.4 package.scala 96:25:@25715.4]
  assign _T_365 = io_rr ? _T_363 : 1'h0; // @[implicits.scala 55:10:@25716.4]
  assign _T_366 = _T_359 & _T_365; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:118:@25717.4]
  assign _T_368 = _T_366 & _T_359; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:206:@25719.4]
  assign _T_369 = _T_368 & io_sigsIn_backpressure; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:225:@25720.4]
  assign x490_b254_D3 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@25703.4 package.scala 96:25:@25704.4]
  assign _T_370 = _T_369 & x490_b254_D3; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 117:251:@25721.4]
  assign x489_b255_D3 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@25694.4 package.scala 96:25:@25695.4]
  assign x269_rdcol_number = x269_rdcol_1_io_result; // @[Math.scala 154:22:@25738.4 Math.scala 155:14:@25739.4]
  assign _T_387 = $signed(x269_rdcol_number); // @[Math.scala 406:49:@25747.4]
  assign _T_389 = $signed(_T_387) & $signed(32'sh3); // @[Math.scala 406:56:@25749.4]
  assign _T_390 = $signed(_T_389); // @[Math.scala 406:56:@25750.4]
  assign _T_394 = x269_rdcol_number[31]; // @[FixedPoint.scala 50:25:@25756.4]
  assign _T_398 = _T_394 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@25758.4]
  assign _T_399 = x269_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@25759.4]
  assign _T_405 = _T_399 == 30'h3fffffff; // @[Math.scala 451:55:@25761.4]
  assign _T_406 = x269_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@25762.4]
  assign _T_412 = _T_406 != 2'h0; // @[Math.scala 451:110:@25764.4]
  assign _T_413 = _T_405 & _T_412; // @[Math.scala 451:94:@25765.4]
  assign _T_415 = {_T_398,_T_399}; // @[Cat.scala 30:58:@25767.4]
  assign _T_435 = RetimeWrapper_12_io_out; // @[package.scala 96:25:@25816.4 package.scala 96:25:@25817.4]
  assign _T_437 = io_rr ? _T_435 : 1'h0; // @[implicits.scala 55:10:@25818.4]
  assign _T_438 = _T_359 & _T_437; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 138:118:@25819.4]
  assign _T_440 = _T_438 & _T_359; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 138:206:@25821.4]
  assign _T_441 = _T_440 & io_sigsIn_backpressure; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 138:225:@25822.4]
  assign _T_442 = _T_441 & x490_b254_D3; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 138:251:@25823.4]
  assign x494_b252_D6_number = RetimeWrapper_13_io_out; // @[package.scala 96:25:@25837.4 package.scala 96:25:@25838.4]
  assign _T_452 = $signed(x494_b252_D6_number); // @[Math.scala 476:37:@25843.4]
  assign x276 = $signed(_T_452) < $signed(32'sh0); // @[Math.scala 476:44:@25845.4]
  assign x495_x269_rdcol_D6_number = RetimeWrapper_14_io_out; // @[package.scala 96:25:@25853.4 package.scala 96:25:@25854.4]
  assign _T_463 = $signed(x495_x269_rdcol_D6_number); // @[Math.scala 476:37:@25859.4]
  assign x277 = $signed(_T_463) < $signed(32'sh0); // @[Math.scala 476:44:@25861.4]
  assign x496_x276_D1 = RetimeWrapper_15_io_out; // @[package.scala 96:25:@25869.4 package.scala 96:25:@25870.4]
  assign x278 = x496_x276_D1 | x277; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 151:24:@25873.4]
  assign _T_502 = RetimeWrapper_22_io_out; // @[package.scala 96:25:@25941.4 package.scala 96:25:@25942.4]
  assign _T_504 = io_rr ? _T_502 : 1'h0; // @[implicits.scala 55:10:@25943.4]
  assign _T_505 = _T_359 & _T_504; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 170:146:@25944.4]
  assign x498_x279_D2 = RetimeWrapper_17_io_out; // @[package.scala 96:25:@25893.4 package.scala 96:25:@25894.4]
  assign _T_506 = _T_505 & x498_x279_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 170:234:@25945.4]
  assign x502_b254_D9 = RetimeWrapper_21_io_out; // @[package.scala 96:25:@25929.4 package.scala 96:25:@25930.4]
  assign _T_507 = _T_506 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 170:242:@25946.4]
  assign x499_b255_D9 = RetimeWrapper_18_io_out; // @[package.scala 96:25:@25902.4 package.scala 96:25:@25903.4]
  assign x503_b253_D6_number = RetimeWrapper_23_io_out; // @[package.scala 96:25:@25962.4 package.scala 96:25:@25963.4]
  assign _T_520 = $signed(x503_b253_D6_number); // @[Math.scala 476:37:@25970.4]
  assign x282 = $signed(_T_520) < $signed(32'sh0); // @[Math.scala 476:44:@25972.4]
  assign x283 = x276 | x282; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 186:59:@25975.4]
  assign _T_547 = RetimeWrapper_27_io_out; // @[package.scala 96:25:@26016.4 package.scala 96:25:@26017.4]
  assign _T_549 = io_rr ? _T_547 : 1'h0; // @[implicits.scala 55:10:@26018.4]
  assign _T_550 = _T_359 & _T_549; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 199:194:@26019.4]
  assign x504_x284_D3 = RetimeWrapper_24_io_out; // @[package.scala 96:25:@25986.4 package.scala 96:25:@25987.4]
  assign _T_551 = _T_550 & x504_x284_D3; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 199:282:@26020.4]
  assign _T_552 = _T_551 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 199:290:@26021.4]
  assign x287_rdcol_number = x287_rdcol_1_io_result; // @[Math.scala 154:22:@26040.4 Math.scala 155:14:@26041.4]
  assign _T_567 = $signed(x287_rdcol_number); // @[Math.scala 476:37:@26046.4]
  assign x288 = $signed(_T_567) < $signed(32'sh0); // @[Math.scala 476:44:@26048.4]
  assign x289 = x496_x276_D1 | x288; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 207:59:@26051.4]
  assign _T_583 = $signed(_T_567) & $signed(32'sh3); // @[Math.scala 406:56:@26062.4]
  assign _T_584 = $signed(_T_583); // @[Math.scala 406:56:@26063.4]
  assign _T_588 = x287_rdcol_number[31]; // @[FixedPoint.scala 50:25:@26069.4]
  assign _T_592 = _T_588 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26071.4]
  assign _T_593 = x287_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@26072.4]
  assign _T_599 = _T_593 == 30'h3fffffff; // @[Math.scala 451:55:@26074.4]
  assign _T_600 = x287_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@26075.4]
  assign _T_606 = _T_600 != 2'h0; // @[Math.scala 451:110:@26077.4]
  assign _T_607 = _T_599 & _T_606; // @[Math.scala 451:94:@26078.4]
  assign _T_609 = {_T_592,_T_593}; // @[Cat.scala 30:58:@26080.4]
  assign _T_638 = RetimeWrapper_32_io_out; // @[package.scala 96:25:@26139.4 package.scala 96:25:@26140.4]
  assign _T_640 = io_rr ? _T_638 : 1'h0; // @[implicits.scala 55:10:@26141.4]
  assign _T_641 = _T_359 & _T_640; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 228:194:@26142.4]
  assign x510_x290_D2 = RetimeWrapper_31_io_out; // @[package.scala 96:25:@26127.4 package.scala 96:25:@26128.4]
  assign _T_642 = _T_641 & x510_x290_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 228:282:@26143.4]
  assign _T_643 = _T_642 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 228:290:@26144.4]
  assign x296_rdcol_number = x296_rdcol_1_io_result; // @[Math.scala 154:22:@26163.4 Math.scala 155:14:@26164.4]
  assign _T_658 = $signed(x296_rdcol_number); // @[Math.scala 476:37:@26169.4]
  assign x297 = $signed(_T_658) < $signed(32'sh0); // @[Math.scala 476:44:@26171.4]
  assign x298 = x496_x276_D1 | x297; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 236:59:@26174.4]
  assign _T_674 = $signed(_T_658) & $signed(32'sh3); // @[Math.scala 406:56:@26185.4]
  assign _T_675 = $signed(_T_674); // @[Math.scala 406:56:@26186.4]
  assign _T_679 = x296_rdcol_number[31]; // @[FixedPoint.scala 50:25:@26192.4]
  assign _T_683 = _T_679 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26194.4]
  assign _T_684 = x296_rdcol_number[31:2]; // @[FixedPoint.scala 18:52:@26195.4]
  assign _T_690 = _T_684 == 30'h3fffffff; // @[Math.scala 451:55:@26197.4]
  assign _T_691 = x296_rdcol_number[1:0]; // @[FixedPoint.scala 18:52:@26198.4]
  assign _T_697 = _T_691 != 2'h0; // @[Math.scala 451:110:@26200.4]
  assign _T_698 = _T_690 & _T_697; // @[Math.scala 451:94:@26201.4]
  assign _T_700 = {_T_683,_T_684}; // @[Cat.scala 30:58:@26203.4]
  assign _T_726 = RetimeWrapper_36_io_out; // @[package.scala 96:25:@26253.4 package.scala 96:25:@26254.4]
  assign _T_728 = io_rr ? _T_726 : 1'h0; // @[implicits.scala 55:10:@26255.4]
  assign _T_729 = _T_359 & _T_728; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 255:194:@26256.4]
  assign x513_x299_D2 = RetimeWrapper_35_io_out; // @[package.scala 96:25:@26241.4 package.scala 96:25:@26242.4]
  assign _T_730 = _T_729 & x513_x299_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 255:282:@26257.4]
  assign _T_731 = _T_730 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 255:290:@26258.4]
  assign x305_rdrow_number = x305_rdrow_1_io_result; // @[Math.scala 195:22:@26277.4 Math.scala 196:14:@26278.4]
  assign _T_748 = $signed(x305_rdrow_number); // @[Math.scala 406:49:@26284.4]
  assign _T_750 = $signed(_T_748) & $signed(32'sh3); // @[Math.scala 406:56:@26286.4]
  assign _T_751 = $signed(_T_750); // @[Math.scala 406:56:@26287.4]
  assign x468_number = $unsigned(_T_751); // @[implicits.scala 133:21:@26288.4]
  assign x307 = $signed(_T_748) < $signed(32'sh0); // @[Math.scala 476:44:@26296.4]
  assign x308 = x307 | x277; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 265:24:@26299.4]
  assign _T_772 = $signed(x468_number); // @[Math.scala 406:49:@26308.4]
  assign _T_774 = $signed(_T_772) & $signed(32'sh3); // @[Math.scala 406:56:@26310.4]
  assign _T_775 = $signed(_T_774); // @[Math.scala 406:56:@26311.4]
  assign _T_779 = x468_number[31]; // @[FixedPoint.scala 50:25:@26317.4]
  assign _T_783 = _T_779 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26319.4]
  assign _T_784 = x468_number[31:2]; // @[FixedPoint.scala 18:52:@26320.4]
  assign _T_790 = _T_784 == 30'h3fffffff; // @[Math.scala 451:55:@26322.4]
  assign _T_791 = x468_number[1:0]; // @[FixedPoint.scala 18:52:@26323.4]
  assign _T_797 = _T_791 != 2'h0; // @[Math.scala 451:110:@26325.4]
  assign _T_798 = _T_790 & _T_797; // @[Math.scala 451:94:@26326.4]
  assign _T_800 = {_T_783,_T_784}; // @[Cat.scala 30:58:@26328.4]
  assign x311_1_number = _T_798 ? 32'h0 : _T_800; // @[Math.scala 454:20:@26329.4]
  assign _GEN_2 = {{9'd0}, x311_1_number}; // @[Math.scala 461:32:@26334.4]
  assign _T_805 = _GEN_2 << 9; // @[Math.scala 461:32:@26334.4]
  assign _GEN_3 = {{5'd0}, x311_1_number}; // @[Math.scala 461:32:@26339.4]
  assign _T_808 = _GEN_3 << 5; // @[Math.scala 461:32:@26339.4]
  assign _T_835 = RetimeWrapper_40_io_out; // @[package.scala 96:25:@26398.4 package.scala 96:25:@26399.4]
  assign _T_837 = io_rr ? _T_835 : 1'h0; // @[implicits.scala 55:10:@26400.4]
  assign _T_838 = _T_359 & _T_837; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 290:194:@26401.4]
  assign x516_x309_D2 = RetimeWrapper_39_io_out; // @[package.scala 96:25:@26386.4 package.scala 96:25:@26387.4]
  assign _T_839 = _T_838 & x516_x309_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 290:282:@26402.4]
  assign _T_840 = _T_839 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 290:290:@26403.4]
  assign x517_x282_D1 = RetimeWrapper_41_io_out; // @[package.scala 96:25:@26419.4 package.scala 96:25:@26420.4]
  assign x316 = x307 | x517_x282_D1; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 302:59:@26423.4]
  assign _T_872 = RetimeWrapper_44_io_out; // @[package.scala 96:25:@26467.4 package.scala 96:25:@26468.4]
  assign _T_874 = io_rr ? _T_872 : 1'h0; // @[implicits.scala 55:10:@26469.4]
  assign _T_875 = _T_359 & _T_874; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 317:194:@26470.4]
  assign x519_x317_D2 = RetimeWrapper_43_io_out; // @[package.scala 96:25:@26455.4 package.scala 96:25:@26456.4]
  assign _T_876 = _T_875 & x519_x317_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 317:282:@26471.4]
  assign _T_877 = _T_876 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 317:290:@26472.4]
  assign x321 = x307 | x288; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 321:59:@26483.4]
  assign _T_904 = RetimeWrapper_47_io_out; // @[package.scala 96:25:@26525.4 package.scala 96:25:@26526.4]
  assign _T_906 = io_rr ? _T_904 : 1'h0; // @[implicits.scala 55:10:@26527.4]
  assign _T_907 = _T_359 & _T_906; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 334:194:@26528.4]
  assign x521_x322_D2 = RetimeWrapper_46_io_out; // @[package.scala 96:25:@26513.4 package.scala 96:25:@26514.4]
  assign _T_908 = _T_907 & x521_x322_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 334:282:@26529.4]
  assign _T_909 = _T_908 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 334:290:@26530.4]
  assign x326 = x307 | x297; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 338:59:@26541.4]
  assign _T_936 = RetimeWrapper_50_io_out; // @[package.scala 96:25:@26583.4 package.scala 96:25:@26584.4]
  assign _T_938 = io_rr ? _T_936 : 1'h0; // @[implicits.scala 55:10:@26585.4]
  assign _T_939 = _T_359 & _T_938; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 351:194:@26586.4]
  assign x523_x327_D2 = RetimeWrapper_49_io_out; // @[package.scala 96:25:@26571.4 package.scala 96:25:@26572.4]
  assign _T_940 = _T_939 & x523_x327_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 351:282:@26587.4]
  assign _T_941 = _T_940 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 351:290:@26588.4]
  assign x331_rdrow_number = x331_rdrow_1_io_result; // @[Math.scala 195:22:@26607.4 Math.scala 196:14:@26608.4]
  assign _T_958 = $signed(x331_rdrow_number); // @[Math.scala 406:49:@26614.4]
  assign _T_960 = $signed(_T_958) & $signed(32'sh3); // @[Math.scala 406:56:@26616.4]
  assign _T_961 = $signed(_T_960); // @[Math.scala 406:56:@26617.4]
  assign x473_number = $unsigned(_T_961); // @[implicits.scala 133:21:@26618.4]
  assign x333 = $signed(_T_958) < $signed(32'sh0); // @[Math.scala 476:44:@26626.4]
  assign x334 = x333 | x277; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 361:24:@26629.4]
  assign _T_982 = $signed(x473_number); // @[Math.scala 406:49:@26638.4]
  assign _T_984 = $signed(_T_982) & $signed(32'sh3); // @[Math.scala 406:56:@26640.4]
  assign _T_985 = $signed(_T_984); // @[Math.scala 406:56:@26641.4]
  assign _T_989 = x473_number[31]; // @[FixedPoint.scala 50:25:@26647.4]
  assign _T_993 = _T_989 ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12:@26649.4]
  assign _T_994 = x473_number[31:2]; // @[FixedPoint.scala 18:52:@26650.4]
  assign _T_1000 = _T_994 == 30'h3fffffff; // @[Math.scala 451:55:@26652.4]
  assign _T_1001 = x473_number[1:0]; // @[FixedPoint.scala 18:52:@26653.4]
  assign _T_1007 = _T_1001 != 2'h0; // @[Math.scala 451:110:@26655.4]
  assign _T_1008 = _T_1000 & _T_1007; // @[Math.scala 451:94:@26656.4]
  assign _T_1010 = {_T_993,_T_994}; // @[Cat.scala 30:58:@26658.4]
  assign x337_1_number = _T_1008 ? 32'h0 : _T_1010; // @[Math.scala 454:20:@26659.4]
  assign _GEN_4 = {{9'd0}, x337_1_number}; // @[Math.scala 461:32:@26664.4]
  assign _T_1015 = _GEN_4 << 9; // @[Math.scala 461:32:@26664.4]
  assign _GEN_5 = {{5'd0}, x337_1_number}; // @[Math.scala 461:32:@26669.4]
  assign _T_1018 = _GEN_5 << 5; // @[Math.scala 461:32:@26669.4]
  assign _T_1042 = RetimeWrapper_53_io_out; // @[package.scala 96:25:@26719.4 package.scala 96:25:@26720.4]
  assign _T_1044 = io_rr ? _T_1042 : 1'h0; // @[implicits.scala 55:10:@26721.4]
  assign _T_1045 = _T_359 & _T_1044; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 384:194:@26722.4]
  assign x524_x335_D2 = RetimeWrapper_51_io_out; // @[package.scala 96:25:@26698.4 package.scala 96:25:@26699.4]
  assign _T_1046 = _T_1045 & x524_x335_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 384:282:@26723.4]
  assign _T_1047 = _T_1046 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 384:290:@26724.4]
  assign x342 = x333 | x517_x282_D1; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 388:24:@26735.4]
  assign _T_1071 = RetimeWrapper_55_io_out; // @[package.scala 96:25:@26768.4 package.scala 96:25:@26769.4]
  assign _T_1073 = io_rr ? _T_1071 : 1'h0; // @[implicits.scala 55:10:@26770.4]
  assign _T_1074 = _T_359 & _T_1073; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 399:194:@26771.4]
  assign x526_x343_D2 = RetimeWrapper_54_io_out; // @[package.scala 96:25:@26756.4 package.scala 96:25:@26757.4]
  assign _T_1075 = _T_1074 & x526_x343_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 399:282:@26772.4]
  assign _T_1076 = _T_1075 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 399:290:@26773.4]
  assign x347 = x333 | x288; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 403:24:@26784.4]
  assign _T_1100 = RetimeWrapper_57_io_out; // @[package.scala 96:25:@26817.4 package.scala 96:25:@26818.4]
  assign _T_1102 = io_rr ? _T_1100 : 1'h0; // @[implicits.scala 55:10:@26819.4]
  assign _T_1103 = _T_359 & _T_1102; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 414:194:@26820.4]
  assign x527_x348_D2 = RetimeWrapper_56_io_out; // @[package.scala 96:25:@26805.4 package.scala 96:25:@26806.4]
  assign _T_1104 = _T_1103 & x527_x348_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 414:282:@26821.4]
  assign _T_1105 = _T_1104 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 414:290:@26822.4]
  assign x352 = x333 | x297; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 424:59:@26833.4]
  assign _T_1131 = RetimeWrapper_59_io_out; // @[package.scala 96:25:@26868.4 package.scala 96:25:@26869.4]
  assign _T_1133 = io_rr ? _T_1131 : 1'h0; // @[implicits.scala 55:10:@26870.4]
  assign _T_1134 = _T_359 & _T_1133; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 437:194:@26871.4]
  assign x528_x353_D2 = RetimeWrapper_58_io_out; // @[package.scala 96:25:@26856.4 package.scala 96:25:@26857.4]
  assign _T_1135 = _T_1134 & x528_x353_D2; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 437:282:@26872.4]
  assign _T_1136 = _T_1135 & x502_b254_D9; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 437:290:@26873.4]
  assign x376_number = x376_1_io_result; // @[Math.scala 723:22:@27107.4 Math.scala 724:14:@27108.4]
  assign x396_number = x396_1_io_result; // @[Math.scala 723:22:@27334.4 Math.scala 724:14:@27335.4]
  assign _T_1366 = RetimeWrapper_65_io_out; // @[package.scala 96:25:@27376.4 package.scala 96:25:@27377.4]
  assign _T_1368 = io_rr ? _T_1366 : 1'h0; // @[implicits.scala 55:10:@27378.4]
  assign x531_b254_D30 = RetimeWrapper_63_io_out; // @[package.scala 96:25:@27358.4 package.scala 96:25:@27359.4]
  assign _T_1369 = _T_1368 & x531_b254_D30; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 539:117:@27379.4]
  assign x532_b255_D30 = RetimeWrapper_64_io_out; // @[package.scala 96:25:@27367.4 package.scala 96:25:@27368.4]
  assign _T_1370 = _T_1369 & x532_b255_D30; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 539:123:@27380.4]
  assign x485_x460_D3_number = RetimeWrapper_2_io_out; // @[package.scala 96:25:@25658.4 package.scala 96:25:@25659.4]
  assign x487_x461_D3_number = RetimeWrapper_4_io_out; // @[package.scala 96:25:@25676.4 package.scala 96:25:@25677.4]
  assign x488_x267_sum_D1_number = RetimeWrapper_5_io_out; // @[package.scala 96:25:@25685.4 package.scala 96:25:@25686.4]
  assign x492_x465_D2_number = RetimeWrapper_10_io_out; // @[package.scala 96:25:@25796.4 package.scala 96:25:@25797.4]
  assign x493_x273_sum_D1_number = RetimeWrapper_11_io_out; // @[package.scala 96:25:@25805.4 package.scala 96:25:@25806.4]
  assign x497_x460_D9_number = RetimeWrapper_16_io_out; // @[package.scala 96:25:@25884.4 package.scala 96:25:@25885.4]
  assign x500_x465_D8_number = RetimeWrapper_19_io_out; // @[package.scala 96:25:@25911.4 package.scala 96:25:@25912.4]
  assign x501_x273_sum_D7_number = RetimeWrapper_20_io_out; // @[package.scala 96:25:@25920.4 package.scala 96:25:@25921.4]
  assign x505_x461_D9_number = RetimeWrapper_25_io_out; // @[package.scala 96:25:@25995.4 package.scala 96:25:@25996.4]
  assign x506_x267_sum_D7_number = RetimeWrapper_26_io_out; // @[package.scala 96:25:@26004.4 package.scala 96:25:@26005.4]
  assign x508_x293_sum_D1_number = RetimeWrapper_29_io_out; // @[package.scala 96:25:@26109.4 package.scala 96:25:@26110.4]
  assign x509_x466_D2_number = RetimeWrapper_30_io_out; // @[package.scala 96:25:@26118.4 package.scala 96:25:@26119.4]
  assign x511_x302_sum_D1_number = RetimeWrapper_33_io_out; // @[package.scala 96:25:@26223.4 package.scala 96:25:@26224.4]
  assign x512_x467_D2_number = RetimeWrapper_34_io_out; // @[package.scala 96:25:@26232.4 package.scala 96:25:@26233.4]
  assign x313_sum_number = x313_sum_1_io_result; // @[Math.scala 154:22:@26368.4 Math.scala 155:14:@26369.4]
  assign x515_x469_D2_number = RetimeWrapper_38_io_out; // @[package.scala 96:25:@26377.4 package.scala 96:25:@26378.4]
  assign x318_sum_number = x318_sum_1_io_result; // @[Math.scala 154:22:@26446.4 Math.scala 155:14:@26447.4]
  assign x323_sum_number = x323_sum_1_io_result; // @[Math.scala 154:22:@26504.4 Math.scala 155:14:@26505.4]
  assign x328_sum_number = x328_sum_1_io_result; // @[Math.scala 154:22:@26562.4 Math.scala 155:14:@26563.4]
  assign x339_sum_number = x339_sum_1_io_result; // @[Math.scala 154:22:@26689.4 Math.scala 155:14:@26690.4]
  assign x525_x474_D2_number = RetimeWrapper_52_io_out; // @[package.scala 96:25:@26707.4 package.scala 96:25:@26708.4]
  assign x344_sum_number = x344_sum_1_io_result; // @[Math.scala 154:22:@26747.4 Math.scala 155:14:@26748.4]
  assign x349_sum_number = x349_sum_1_io_result; // @[Math.scala 154:22:@26796.4 Math.scala 155:14:@26797.4]
  assign x354_sum_number = x354_sum_1_io_result; // @[Math.scala 154:22:@26847.4 Math.scala 155:14:@26848.4]
  assign io_in_x221_TREADY = _T_211 & _T_213; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 67:22:@25424.4 sm_x401_inr_Foreach_SAMPLER_BOX.scala 69:22:@25432.4]
  assign io_in_x222_TVALID = _T_1370 & io_sigsIn_backpressure; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 539:22:@27382.4]
  assign io_in_x222_TDATA = {{192'd0}, RetimeWrapper_62_io_out}; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 540:24:@27383.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@25402.4]
  assign __1_io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_1); // @[Math.scala 721:17:@25414.4]
  assign RetimeWrapper_clock = clock; // @[:@25435.4]
  assign RetimeWrapper_reset = reset; // @[:@25436.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25438.4]
  assign RetimeWrapper_io_in = io_in_x221_TDATA[63:0]; // @[package.scala 94:16:@25437.4]
  assign x258_lb_0_clock = clock; // @[:@25445.4]
  assign x258_lb_0_reset = reset; // @[:@25446.4]
  assign x258_lb_0_io_rPort_11_banks_1 = x509_x466_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26147.4]
  assign x258_lb_0_io_rPort_11_banks_0 = x497_x460_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26146.4]
  assign x258_lb_0_io_rPort_11_ofs_0 = x508_x293_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@26148.4]
  assign x258_lb_0_io_rPort_11_en_0 = _T_643 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26150.4]
  assign x258_lb_0_io_rPort_11_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26149.4]
  assign x258_lb_0_io_rPort_10_banks_1 = x505_x461_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26475.4]
  assign x258_lb_0_io_rPort_10_banks_0 = x515_x469_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26474.4]
  assign x258_lb_0_io_rPort_10_ofs_0 = x318_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@26476.4]
  assign x258_lb_0_io_rPort_10_en_0 = _T_877 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26478.4]
  assign x258_lb_0_io_rPort_10_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26477.4]
  assign x258_lb_0_io_rPort_9_banks_1 = x500_x465_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@26406.4]
  assign x258_lb_0_io_rPort_9_banks_0 = x515_x469_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26405.4]
  assign x258_lb_0_io_rPort_9_ofs_0 = x313_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@26407.4]
  assign x258_lb_0_io_rPort_9_en_0 = _T_840 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26409.4]
  assign x258_lb_0_io_rPort_9_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26408.4]
  assign x258_lb_0_io_rPort_8_banks_1 = x512_x467_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26876.4]
  assign x258_lb_0_io_rPort_8_banks_0 = x525_x474_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26875.4]
  assign x258_lb_0_io_rPort_8_ofs_0 = x354_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@26877.4]
  assign x258_lb_0_io_rPort_8_en_0 = _T_1136 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26879.4]
  assign x258_lb_0_io_rPort_8_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26878.4]
  assign x258_lb_0_io_rPort_7_banks_1 = x505_x461_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26776.4]
  assign x258_lb_0_io_rPort_7_banks_0 = x525_x474_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26775.4]
  assign x258_lb_0_io_rPort_7_ofs_0 = x344_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@26777.4]
  assign x258_lb_0_io_rPort_7_en_0 = _T_1076 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26779.4]
  assign x258_lb_0_io_rPort_7_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26778.4]
  assign x258_lb_0_io_rPort_6_banks_1 = x512_x467_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26261.4]
  assign x258_lb_0_io_rPort_6_banks_0 = x497_x460_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26260.4]
  assign x258_lb_0_io_rPort_6_ofs_0 = x511_x302_sum_D1_number[8:0]; // @[MemInterfaceType.scala 107:54:@26262.4]
  assign x258_lb_0_io_rPort_6_en_0 = _T_731 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26264.4]
  assign x258_lb_0_io_rPort_6_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26263.4]
  assign x258_lb_0_io_rPort_5_banks_1 = x509_x466_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26825.4]
  assign x258_lb_0_io_rPort_5_banks_0 = x525_x474_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26824.4]
  assign x258_lb_0_io_rPort_5_ofs_0 = x349_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@26826.4]
  assign x258_lb_0_io_rPort_5_en_0 = _T_1105 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26828.4]
  assign x258_lb_0_io_rPort_5_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26827.4]
  assign x258_lb_0_io_rPort_4_banks_1 = x505_x461_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26024.4]
  assign x258_lb_0_io_rPort_4_banks_0 = x497_x460_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@26023.4]
  assign x258_lb_0_io_rPort_4_ofs_0 = x506_x267_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@26025.4]
  assign x258_lb_0_io_rPort_4_en_0 = _T_552 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26027.4]
  assign x258_lb_0_io_rPort_4_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26026.4]
  assign x258_lb_0_io_rPort_3_banks_1 = x509_x466_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26533.4]
  assign x258_lb_0_io_rPort_3_banks_0 = x515_x469_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26532.4]
  assign x258_lb_0_io_rPort_3_ofs_0 = x323_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@26534.4]
  assign x258_lb_0_io_rPort_3_en_0 = _T_909 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26536.4]
  assign x258_lb_0_io_rPort_3_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26535.4]
  assign x258_lb_0_io_rPort_2_banks_1 = x512_x467_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26591.4]
  assign x258_lb_0_io_rPort_2_banks_0 = x515_x469_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26590.4]
  assign x258_lb_0_io_rPort_2_ofs_0 = x328_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@26592.4]
  assign x258_lb_0_io_rPort_2_en_0 = _T_941 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26594.4]
  assign x258_lb_0_io_rPort_2_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26593.4]
  assign x258_lb_0_io_rPort_1_banks_1 = x500_x465_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@25949.4]
  assign x258_lb_0_io_rPort_1_banks_0 = x497_x460_D9_number[2:0]; // @[MemInterfaceType.scala 106:58:@25948.4]
  assign x258_lb_0_io_rPort_1_ofs_0 = x501_x273_sum_D7_number[8:0]; // @[MemInterfaceType.scala 107:54:@25950.4]
  assign x258_lb_0_io_rPort_1_en_0 = _T_507 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@25952.4]
  assign x258_lb_0_io_rPort_1_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@25951.4]
  assign x258_lb_0_io_rPort_0_banks_1 = x500_x465_D8_number[2:0]; // @[MemInterfaceType.scala 106:58:@26727.4]
  assign x258_lb_0_io_rPort_0_banks_0 = x525_x474_D2_number[2:0]; // @[MemInterfaceType.scala 106:58:@26726.4]
  assign x258_lb_0_io_rPort_0_ofs_0 = x339_sum_number[8:0]; // @[MemInterfaceType.scala 107:54:@26728.4]
  assign x258_lb_0_io_rPort_0_en_0 = _T_1047 & x499_b255_D9; // @[MemInterfaceType.scala 110:79:@26730.4]
  assign x258_lb_0_io_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@26729.4]
  assign x258_lb_0_io_wPort_1_banks_1 = x492_x465_D2_number[2:0]; // @[MemInterfaceType.scala 88:58:@25826.4]
  assign x258_lb_0_io_wPort_1_banks_0 = x485_x460_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@25825.4]
  assign x258_lb_0_io_wPort_1_ofs_0 = x493_x273_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@25827.4]
  assign x258_lb_0_io_wPort_1_data_0 = RetimeWrapper_9_io_out; // @[MemInterfaceType.scala 90:56:@25828.4]
  assign x258_lb_0_io_wPort_1_en_0 = _T_442 & x489_b255_D3; // @[MemInterfaceType.scala 93:57:@25830.4]
  assign x258_lb_0_io_wPort_0_banks_1 = x487_x461_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@25724.4]
  assign x258_lb_0_io_wPort_0_banks_0 = x485_x460_D3_number[2:0]; // @[MemInterfaceType.scala 88:58:@25723.4]
  assign x258_lb_0_io_wPort_0_ofs_0 = x488_x267_sum_D1_number[8:0]; // @[MemInterfaceType.scala 89:54:@25725.4]
  assign x258_lb_0_io_wPort_0_data_0 = RetimeWrapper_3_io_out; // @[MemInterfaceType.scala 90:56:@25726.4]
  assign x258_lb_0_io_wPort_0_en_0 = _T_370 & x489_b255_D3; // @[MemInterfaceType.scala 93:57:@25728.4]
  assign x464_sub_1_clock = clock; // @[:@25608.4]
  assign x464_sub_1_reset = reset; // @[:@25609.4]
  assign x464_sub_1_io_a = _T_301[31:0]; // @[Math.scala 192:17:@25610.4]
  assign x464_sub_1_io_b = _T_304[31:0]; // @[Math.scala 193:17:@25611.4]
  assign x464_sub_1_io_flow = io_in_x222_TREADY; // @[Math.scala 194:20:@25612.4]
  assign RetimeWrapper_1_clock = clock; // @[:@25635.4]
  assign RetimeWrapper_1_reset = reset; // @[:@25636.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25638.4]
  assign RetimeWrapper_1_io_in = _T_329 ? 32'h0 : _T_331; // @[package.scala 94:16:@25637.4]
  assign x267_sum_1_clock = clock; // @[:@25644.4]
  assign x267_sum_1_reset = reset; // @[:@25645.4]
  assign x267_sum_1_io_a = x464_sub_1_io_result; // @[Math.scala 151:17:@25646.4]
  assign x267_sum_1_io_b = RetimeWrapper_1_io_out; // @[Math.scala 152:17:@25647.4]
  assign x267_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@25648.4]
  assign RetimeWrapper_2_clock = clock; // @[:@25654.4]
  assign RetimeWrapper_2_reset = reset; // @[:@25655.4]
  assign RetimeWrapper_2_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25657.4]
  assign RetimeWrapper_2_io_in = $unsigned(_T_259); // @[package.scala 94:16:@25656.4]
  assign RetimeWrapper_3_clock = clock; // @[:@25663.4]
  assign RetimeWrapper_3_reset = reset; // @[:@25664.4]
  assign RetimeWrapper_3_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25666.4]
  assign RetimeWrapper_3_io_in = x483_x256_D1_0_number[31:0]; // @[package.scala 94:16:@25665.4]
  assign RetimeWrapper_4_clock = clock; // @[:@25672.4]
  assign RetimeWrapper_4_reset = reset; // @[:@25673.4]
  assign RetimeWrapper_4_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25675.4]
  assign RetimeWrapper_4_io_in = $unsigned(_T_271); // @[package.scala 94:16:@25674.4]
  assign RetimeWrapper_5_clock = clock; // @[:@25681.4]
  assign RetimeWrapper_5_reset = reset; // @[:@25682.4]
  assign RetimeWrapper_5_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25684.4]
  assign RetimeWrapper_5_io_in = x267_sum_1_io_result; // @[package.scala 94:16:@25683.4]
  assign RetimeWrapper_6_clock = clock; // @[:@25690.4]
  assign RetimeWrapper_6_reset = reset; // @[:@25691.4]
  assign RetimeWrapper_6_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25693.4]
  assign RetimeWrapper_6_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@25692.4]
  assign RetimeWrapper_7_clock = clock; // @[:@25699.4]
  assign RetimeWrapper_7_reset = reset; // @[:@25700.4]
  assign RetimeWrapper_7_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25702.4]
  assign RetimeWrapper_7_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@25701.4]
  assign RetimeWrapper_8_clock = clock; // @[:@25710.4]
  assign RetimeWrapper_8_reset = reset; // @[:@25711.4]
  assign RetimeWrapper_8_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25713.4]
  assign RetimeWrapper_8_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25712.4]
  assign x269_rdcol_1_clock = clock; // @[:@25733.4]
  assign x269_rdcol_1_reset = reset; // @[:@25734.4]
  assign x269_rdcol_1_io_a = __1_io_result; // @[Math.scala 151:17:@25735.4]
  assign x269_rdcol_1_io_b = 32'h1; // @[Math.scala 152:17:@25736.4]
  assign x269_rdcol_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@25737.4]
  assign x273_sum_1_clock = clock; // @[:@25773.4]
  assign x273_sum_1_reset = reset; // @[:@25774.4]
  assign x273_sum_1_io_a = x464_sub_1_io_result; // @[Math.scala 151:17:@25775.4]
  assign x273_sum_1_io_b = _T_413 ? 32'h0 : _T_415; // @[Math.scala 152:17:@25776.4]
  assign x273_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@25777.4]
  assign RetimeWrapper_9_clock = clock; // @[:@25783.4]
  assign RetimeWrapper_9_reset = reset; // @[:@25784.4]
  assign RetimeWrapper_9_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25786.4]
  assign RetimeWrapper_9_io_in = x483_x256_D1_0_number[63:32]; // @[package.scala 94:16:@25785.4]
  assign RetimeWrapper_10_clock = clock; // @[:@25792.4]
  assign RetimeWrapper_10_reset = reset; // @[:@25793.4]
  assign RetimeWrapper_10_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25795.4]
  assign RetimeWrapper_10_io_in = $unsigned(_T_390); // @[package.scala 94:16:@25794.4]
  assign RetimeWrapper_11_clock = clock; // @[:@25801.4]
  assign RetimeWrapper_11_reset = reset; // @[:@25802.4]
  assign RetimeWrapper_11_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25804.4]
  assign RetimeWrapper_11_io_in = x273_sum_1_io_result; // @[package.scala 94:16:@25803.4]
  assign RetimeWrapper_12_clock = clock; // @[:@25812.4]
  assign RetimeWrapper_12_reset = reset; // @[:@25813.4]
  assign RetimeWrapper_12_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25815.4]
  assign RetimeWrapper_12_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25814.4]
  assign RetimeWrapper_13_clock = clock; // @[:@25833.4]
  assign RetimeWrapper_13_reset = reset; // @[:@25834.4]
  assign RetimeWrapper_13_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25836.4]
  assign RetimeWrapper_13_io_in = __io_result; // @[package.scala 94:16:@25835.4]
  assign RetimeWrapper_14_clock = clock; // @[:@25849.4]
  assign RetimeWrapper_14_reset = reset; // @[:@25850.4]
  assign RetimeWrapper_14_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25852.4]
  assign RetimeWrapper_14_io_in = x269_rdcol_1_io_result; // @[package.scala 94:16:@25851.4]
  assign RetimeWrapper_15_clock = clock; // @[:@25865.4]
  assign RetimeWrapper_15_reset = reset; // @[:@25866.4]
  assign RetimeWrapper_15_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25868.4]
  assign RetimeWrapper_15_io_in = $signed(_T_452) < $signed(32'sh0); // @[package.scala 94:16:@25867.4]
  assign RetimeWrapper_16_clock = clock; // @[:@25880.4]
  assign RetimeWrapper_16_reset = reset; // @[:@25881.4]
  assign RetimeWrapper_16_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25883.4]
  assign RetimeWrapper_16_io_in = $unsigned(_T_259); // @[package.scala 94:16:@25882.4]
  assign RetimeWrapper_17_clock = clock; // @[:@25889.4]
  assign RetimeWrapper_17_reset = reset; // @[:@25890.4]
  assign RetimeWrapper_17_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25892.4]
  assign RetimeWrapper_17_io_in = ~ x278; // @[package.scala 94:16:@25891.4]
  assign RetimeWrapper_18_clock = clock; // @[:@25898.4]
  assign RetimeWrapper_18_reset = reset; // @[:@25899.4]
  assign RetimeWrapper_18_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25901.4]
  assign RetimeWrapper_18_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@25900.4]
  assign RetimeWrapper_19_clock = clock; // @[:@25907.4]
  assign RetimeWrapper_19_reset = reset; // @[:@25908.4]
  assign RetimeWrapper_19_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25910.4]
  assign RetimeWrapper_19_io_in = $unsigned(_T_390); // @[package.scala 94:16:@25909.4]
  assign RetimeWrapper_20_clock = clock; // @[:@25916.4]
  assign RetimeWrapper_20_reset = reset; // @[:@25917.4]
  assign RetimeWrapper_20_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25919.4]
  assign RetimeWrapper_20_io_in = x273_sum_1_io_result; // @[package.scala 94:16:@25918.4]
  assign RetimeWrapper_21_clock = clock; // @[:@25925.4]
  assign RetimeWrapper_21_reset = reset; // @[:@25926.4]
  assign RetimeWrapper_21_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25928.4]
  assign RetimeWrapper_21_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@25927.4]
  assign RetimeWrapper_22_clock = clock; // @[:@25937.4]
  assign RetimeWrapper_22_reset = reset; // @[:@25938.4]
  assign RetimeWrapper_22_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25940.4]
  assign RetimeWrapper_22_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@25939.4]
  assign RetimeWrapper_23_clock = clock; // @[:@25958.4]
  assign RetimeWrapper_23_reset = reset; // @[:@25959.4]
  assign RetimeWrapper_23_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25961.4]
  assign RetimeWrapper_23_io_in = __1_io_result; // @[package.scala 94:16:@25960.4]
  assign RetimeWrapper_24_clock = clock; // @[:@25982.4]
  assign RetimeWrapper_24_reset = reset; // @[:@25983.4]
  assign RetimeWrapper_24_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25985.4]
  assign RetimeWrapper_24_io_in = ~ x283; // @[package.scala 94:16:@25984.4]
  assign RetimeWrapper_25_clock = clock; // @[:@25991.4]
  assign RetimeWrapper_25_reset = reset; // @[:@25992.4]
  assign RetimeWrapper_25_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@25994.4]
  assign RetimeWrapper_25_io_in = $unsigned(_T_271); // @[package.scala 94:16:@25993.4]
  assign RetimeWrapper_26_clock = clock; // @[:@26000.4]
  assign RetimeWrapper_26_reset = reset; // @[:@26001.4]
  assign RetimeWrapper_26_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26003.4]
  assign RetimeWrapper_26_io_in = x267_sum_1_io_result; // @[package.scala 94:16:@26002.4]
  assign RetimeWrapper_27_clock = clock; // @[:@26012.4]
  assign RetimeWrapper_27_reset = reset; // @[:@26013.4]
  assign RetimeWrapper_27_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26015.4]
  assign RetimeWrapper_27_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26014.4]
  assign x287_rdcol_1_clock = clock; // @[:@26035.4]
  assign x287_rdcol_1_reset = reset; // @[:@26036.4]
  assign x287_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@26037.4]
  assign x287_rdcol_1_io_b = 32'hffffffff; // @[Math.scala 152:17:@26038.4]
  assign x287_rdcol_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26039.4]
  assign RetimeWrapper_28_clock = clock; // @[:@26086.4]
  assign RetimeWrapper_28_reset = reset; // @[:@26087.4]
  assign RetimeWrapper_28_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26089.4]
  assign RetimeWrapper_28_io_in = x464_sub_1_io_result; // @[package.scala 94:16:@26088.4]
  assign x293_sum_1_clock = clock; // @[:@26095.4]
  assign x293_sum_1_reset = reset; // @[:@26096.4]
  assign x293_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@26097.4]
  assign x293_sum_1_io_b = _T_607 ? 32'h0 : _T_609; // @[Math.scala 152:17:@26098.4]
  assign x293_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26099.4]
  assign RetimeWrapper_29_clock = clock; // @[:@26105.4]
  assign RetimeWrapper_29_reset = reset; // @[:@26106.4]
  assign RetimeWrapper_29_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26108.4]
  assign RetimeWrapper_29_io_in = x293_sum_1_io_result; // @[package.scala 94:16:@26107.4]
  assign RetimeWrapper_30_clock = clock; // @[:@26114.4]
  assign RetimeWrapper_30_reset = reset; // @[:@26115.4]
  assign RetimeWrapper_30_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26117.4]
  assign RetimeWrapper_30_io_in = $unsigned(_T_584); // @[package.scala 94:16:@26116.4]
  assign RetimeWrapper_31_clock = clock; // @[:@26123.4]
  assign RetimeWrapper_31_reset = reset; // @[:@26124.4]
  assign RetimeWrapper_31_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26126.4]
  assign RetimeWrapper_31_io_in = ~ x289; // @[package.scala 94:16:@26125.4]
  assign RetimeWrapper_32_clock = clock; // @[:@26135.4]
  assign RetimeWrapper_32_reset = reset; // @[:@26136.4]
  assign RetimeWrapper_32_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26138.4]
  assign RetimeWrapper_32_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26137.4]
  assign x296_rdcol_1_clock = clock; // @[:@26158.4]
  assign x296_rdcol_1_reset = reset; // @[:@26159.4]
  assign x296_rdcol_1_io_a = RetimeWrapper_23_io_out; // @[Math.scala 151:17:@26160.4]
  assign x296_rdcol_1_io_b = 32'hfffffffe; // @[Math.scala 152:17:@26161.4]
  assign x296_rdcol_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26162.4]
  assign x302_sum_1_clock = clock; // @[:@26209.4]
  assign x302_sum_1_reset = reset; // @[:@26210.4]
  assign x302_sum_1_io_a = RetimeWrapper_28_io_out; // @[Math.scala 151:17:@26211.4]
  assign x302_sum_1_io_b = _T_698 ? 32'h0 : _T_700; // @[Math.scala 152:17:@26212.4]
  assign x302_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26213.4]
  assign RetimeWrapper_33_clock = clock; // @[:@26219.4]
  assign RetimeWrapper_33_reset = reset; // @[:@26220.4]
  assign RetimeWrapper_33_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26222.4]
  assign RetimeWrapper_33_io_in = x302_sum_1_io_result; // @[package.scala 94:16:@26221.4]
  assign RetimeWrapper_34_clock = clock; // @[:@26228.4]
  assign RetimeWrapper_34_reset = reset; // @[:@26229.4]
  assign RetimeWrapper_34_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26231.4]
  assign RetimeWrapper_34_io_in = $unsigned(_T_675); // @[package.scala 94:16:@26230.4]
  assign RetimeWrapper_35_clock = clock; // @[:@26237.4]
  assign RetimeWrapper_35_reset = reset; // @[:@26238.4]
  assign RetimeWrapper_35_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26240.4]
  assign RetimeWrapper_35_io_in = ~ x298; // @[package.scala 94:16:@26239.4]
  assign RetimeWrapper_36_clock = clock; // @[:@26249.4]
  assign RetimeWrapper_36_reset = reset; // @[:@26250.4]
  assign RetimeWrapper_36_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26252.4]
  assign RetimeWrapper_36_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26251.4]
  assign x305_rdrow_1_clock = clock; // @[:@26272.4]
  assign x305_rdrow_1_reset = reset; // @[:@26273.4]
  assign x305_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@26274.4]
  assign x305_rdrow_1_io_b = 32'h1; // @[Math.scala 193:17:@26275.4]
  assign x305_rdrow_1_io_flow = io_in_x222_TREADY; // @[Math.scala 194:20:@26276.4]
  assign x472_sub_1_clock = clock; // @[:@26344.4]
  assign x472_sub_1_reset = reset; // @[:@26345.4]
  assign x472_sub_1_io_a = _T_805[31:0]; // @[Math.scala 192:17:@26346.4]
  assign x472_sub_1_io_b = _T_808[31:0]; // @[Math.scala 193:17:@26347.4]
  assign x472_sub_1_io_flow = io_in_x222_TREADY; // @[Math.scala 194:20:@26348.4]
  assign RetimeWrapper_37_clock = clock; // @[:@26354.4]
  assign RetimeWrapper_37_reset = reset; // @[:@26355.4]
  assign RetimeWrapper_37_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26357.4]
  assign RetimeWrapper_37_io_in = _T_413 ? 32'h0 : _T_415; // @[package.scala 94:16:@26356.4]
  assign x313_sum_1_clock = clock; // @[:@26363.4]
  assign x313_sum_1_reset = reset; // @[:@26364.4]
  assign x313_sum_1_io_a = x472_sub_1_io_result; // @[Math.scala 151:17:@26365.4]
  assign x313_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@26366.4]
  assign x313_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26367.4]
  assign RetimeWrapper_38_clock = clock; // @[:@26373.4]
  assign RetimeWrapper_38_reset = reset; // @[:@26374.4]
  assign RetimeWrapper_38_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26376.4]
  assign RetimeWrapper_38_io_in = $unsigned(_T_775); // @[package.scala 94:16:@26375.4]
  assign RetimeWrapper_39_clock = clock; // @[:@26382.4]
  assign RetimeWrapper_39_reset = reset; // @[:@26383.4]
  assign RetimeWrapper_39_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26385.4]
  assign RetimeWrapper_39_io_in = ~ x308; // @[package.scala 94:16:@26384.4]
  assign RetimeWrapper_40_clock = clock; // @[:@26394.4]
  assign RetimeWrapper_40_reset = reset; // @[:@26395.4]
  assign RetimeWrapper_40_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26397.4]
  assign RetimeWrapper_40_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26396.4]
  assign RetimeWrapper_41_clock = clock; // @[:@26415.4]
  assign RetimeWrapper_41_reset = reset; // @[:@26416.4]
  assign RetimeWrapper_41_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26418.4]
  assign RetimeWrapper_41_io_in = $signed(_T_520) < $signed(32'sh0); // @[package.scala 94:16:@26417.4]
  assign RetimeWrapper_42_clock = clock; // @[:@26430.4]
  assign RetimeWrapper_42_reset = reset; // @[:@26431.4]
  assign RetimeWrapper_42_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26433.4]
  assign RetimeWrapper_42_io_in = _T_329 ? 32'h0 : _T_331; // @[package.scala 94:16:@26432.4]
  assign x318_sum_1_clock = clock; // @[:@26441.4]
  assign x318_sum_1_reset = reset; // @[:@26442.4]
  assign x318_sum_1_io_a = x472_sub_1_io_result; // @[Math.scala 151:17:@26443.4]
  assign x318_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@26444.4]
  assign x318_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26445.4]
  assign RetimeWrapper_43_clock = clock; // @[:@26451.4]
  assign RetimeWrapper_43_reset = reset; // @[:@26452.4]
  assign RetimeWrapper_43_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26454.4]
  assign RetimeWrapper_43_io_in = ~ x316; // @[package.scala 94:16:@26453.4]
  assign RetimeWrapper_44_clock = clock; // @[:@26463.4]
  assign RetimeWrapper_44_reset = reset; // @[:@26464.4]
  assign RetimeWrapper_44_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26466.4]
  assign RetimeWrapper_44_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26465.4]
  assign RetimeWrapper_45_clock = clock; // @[:@26490.4]
  assign RetimeWrapper_45_reset = reset; // @[:@26491.4]
  assign RetimeWrapper_45_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26493.4]
  assign RetimeWrapper_45_io_in = _T_607 ? 32'h0 : _T_609; // @[package.scala 94:16:@26492.4]
  assign x323_sum_1_clock = clock; // @[:@26499.4]
  assign x323_sum_1_reset = reset; // @[:@26500.4]
  assign x323_sum_1_io_a = x472_sub_1_io_result; // @[Math.scala 151:17:@26501.4]
  assign x323_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@26502.4]
  assign x323_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26503.4]
  assign RetimeWrapper_46_clock = clock; // @[:@26509.4]
  assign RetimeWrapper_46_reset = reset; // @[:@26510.4]
  assign RetimeWrapper_46_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26512.4]
  assign RetimeWrapper_46_io_in = ~ x321; // @[package.scala 94:16:@26511.4]
  assign RetimeWrapper_47_clock = clock; // @[:@26521.4]
  assign RetimeWrapper_47_reset = reset; // @[:@26522.4]
  assign RetimeWrapper_47_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26524.4]
  assign RetimeWrapper_47_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26523.4]
  assign RetimeWrapper_48_clock = clock; // @[:@26548.4]
  assign RetimeWrapper_48_reset = reset; // @[:@26549.4]
  assign RetimeWrapper_48_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26551.4]
  assign RetimeWrapper_48_io_in = _T_698 ? 32'h0 : _T_700; // @[package.scala 94:16:@26550.4]
  assign x328_sum_1_clock = clock; // @[:@26557.4]
  assign x328_sum_1_reset = reset; // @[:@26558.4]
  assign x328_sum_1_io_a = x472_sub_1_io_result; // @[Math.scala 151:17:@26559.4]
  assign x328_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@26560.4]
  assign x328_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26561.4]
  assign RetimeWrapper_49_clock = clock; // @[:@26567.4]
  assign RetimeWrapper_49_reset = reset; // @[:@26568.4]
  assign RetimeWrapper_49_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26570.4]
  assign RetimeWrapper_49_io_in = ~ x326; // @[package.scala 94:16:@26569.4]
  assign RetimeWrapper_50_clock = clock; // @[:@26579.4]
  assign RetimeWrapper_50_reset = reset; // @[:@26580.4]
  assign RetimeWrapper_50_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26582.4]
  assign RetimeWrapper_50_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26581.4]
  assign x331_rdrow_1_clock = clock; // @[:@26602.4]
  assign x331_rdrow_1_reset = reset; // @[:@26603.4]
  assign x331_rdrow_1_io_a = RetimeWrapper_13_io_out; // @[Math.scala 192:17:@26604.4]
  assign x331_rdrow_1_io_b = 32'h2; // @[Math.scala 193:17:@26605.4]
  assign x331_rdrow_1_io_flow = io_in_x222_TREADY; // @[Math.scala 194:20:@26606.4]
  assign x477_sub_1_clock = clock; // @[:@26674.4]
  assign x477_sub_1_reset = reset; // @[:@26675.4]
  assign x477_sub_1_io_a = _T_1015[31:0]; // @[Math.scala 192:17:@26676.4]
  assign x477_sub_1_io_b = _T_1018[31:0]; // @[Math.scala 193:17:@26677.4]
  assign x477_sub_1_io_flow = io_in_x222_TREADY; // @[Math.scala 194:20:@26678.4]
  assign x339_sum_1_clock = clock; // @[:@26684.4]
  assign x339_sum_1_reset = reset; // @[:@26685.4]
  assign x339_sum_1_io_a = x477_sub_1_io_result; // @[Math.scala 151:17:@26686.4]
  assign x339_sum_1_io_b = RetimeWrapper_37_io_out; // @[Math.scala 152:17:@26687.4]
  assign x339_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26688.4]
  assign RetimeWrapper_51_clock = clock; // @[:@26694.4]
  assign RetimeWrapper_51_reset = reset; // @[:@26695.4]
  assign RetimeWrapper_51_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26697.4]
  assign RetimeWrapper_51_io_in = ~ x334; // @[package.scala 94:16:@26696.4]
  assign RetimeWrapper_52_clock = clock; // @[:@26703.4]
  assign RetimeWrapper_52_reset = reset; // @[:@26704.4]
  assign RetimeWrapper_52_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26706.4]
  assign RetimeWrapper_52_io_in = $unsigned(_T_985); // @[package.scala 94:16:@26705.4]
  assign RetimeWrapper_53_clock = clock; // @[:@26715.4]
  assign RetimeWrapper_53_reset = reset; // @[:@26716.4]
  assign RetimeWrapper_53_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26718.4]
  assign RetimeWrapper_53_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26717.4]
  assign x344_sum_1_clock = clock; // @[:@26742.4]
  assign x344_sum_1_reset = reset; // @[:@26743.4]
  assign x344_sum_1_io_a = x477_sub_1_io_result; // @[Math.scala 151:17:@26744.4]
  assign x344_sum_1_io_b = RetimeWrapper_42_io_out; // @[Math.scala 152:17:@26745.4]
  assign x344_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26746.4]
  assign RetimeWrapper_54_clock = clock; // @[:@26752.4]
  assign RetimeWrapper_54_reset = reset; // @[:@26753.4]
  assign RetimeWrapper_54_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26755.4]
  assign RetimeWrapper_54_io_in = ~ x342; // @[package.scala 94:16:@26754.4]
  assign RetimeWrapper_55_clock = clock; // @[:@26764.4]
  assign RetimeWrapper_55_reset = reset; // @[:@26765.4]
  assign RetimeWrapper_55_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26767.4]
  assign RetimeWrapper_55_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26766.4]
  assign x349_sum_1_clock = clock; // @[:@26791.4]
  assign x349_sum_1_reset = reset; // @[:@26792.4]
  assign x349_sum_1_io_a = x477_sub_1_io_result; // @[Math.scala 151:17:@26793.4]
  assign x349_sum_1_io_b = RetimeWrapper_45_io_out; // @[Math.scala 152:17:@26794.4]
  assign x349_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26795.4]
  assign RetimeWrapper_56_clock = clock; // @[:@26801.4]
  assign RetimeWrapper_56_reset = reset; // @[:@26802.4]
  assign RetimeWrapper_56_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26804.4]
  assign RetimeWrapper_56_io_in = ~ x347; // @[package.scala 94:16:@26803.4]
  assign RetimeWrapper_57_clock = clock; // @[:@26813.4]
  assign RetimeWrapper_57_reset = reset; // @[:@26814.4]
  assign RetimeWrapper_57_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26816.4]
  assign RetimeWrapper_57_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26815.4]
  assign x354_sum_1_clock = clock; // @[:@26842.4]
  assign x354_sum_1_reset = reset; // @[:@26843.4]
  assign x354_sum_1_io_a = x477_sub_1_io_result; // @[Math.scala 151:17:@26844.4]
  assign x354_sum_1_io_b = RetimeWrapper_48_io_out; // @[Math.scala 152:17:@26845.4]
  assign x354_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26846.4]
  assign RetimeWrapper_58_clock = clock; // @[:@26852.4]
  assign RetimeWrapper_58_reset = reset; // @[:@26853.4]
  assign RetimeWrapper_58_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26855.4]
  assign RetimeWrapper_58_io_in = ~ x352; // @[package.scala 94:16:@26854.4]
  assign RetimeWrapper_59_clock = clock; // @[:@26864.4]
  assign RetimeWrapper_59_reset = reset; // @[:@26865.4]
  assign RetimeWrapper_59_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@26867.4]
  assign RetimeWrapper_59_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@26866.4]
  assign x357_1_clock = clock; // @[:@26887.4]
  assign x357_1_io_a = x258_lb_0_io_rPort_1_output_0; // @[Math.scala 263:17:@26889.4]
  assign x357_1_io_b = 32'h1; // @[Math.scala 264:17:@26890.4]
  assign x357_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26891.4]
  assign x358_1_clock = clock; // @[:@26899.4]
  assign x358_1_io_a = x258_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@26901.4]
  assign x358_1_io_b = 32'h2; // @[Math.scala 264:17:@26902.4]
  assign x358_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26903.4]
  assign x359_1_clock = clock; // @[:@26911.4]
  assign x359_1_io_a = x258_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@26913.4]
  assign x359_1_io_b = 32'h1; // @[Math.scala 264:17:@26914.4]
  assign x359_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26915.4]
  assign x360_1_clock = clock; // @[:@26923.4]
  assign x360_1_io_a = x258_lb_0_io_rPort_9_output_0; // @[Math.scala 263:17:@26925.4]
  assign x360_1_io_b = 32'h2; // @[Math.scala 264:17:@26926.4]
  assign x360_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26927.4]
  assign x361_1_clock = clock; // @[:@26935.4]
  assign x361_1_io_a = x258_lb_0_io_rPort_10_output_0; // @[Math.scala 263:17:@26937.4]
  assign x361_1_io_b = 32'h4; // @[Math.scala 264:17:@26938.4]
  assign x361_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26939.4]
  assign x362_1_clock = clock; // @[:@26947.4]
  assign x362_1_io_a = x258_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@26949.4]
  assign x362_1_io_b = 32'h2; // @[Math.scala 264:17:@26950.4]
  assign x362_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26951.4]
  assign x363_1_clock = clock; // @[:@26959.4]
  assign x363_1_io_a = x258_lb_0_io_rPort_0_output_0; // @[Math.scala 263:17:@26961.4]
  assign x363_1_io_b = 32'h1; // @[Math.scala 264:17:@26962.4]
  assign x363_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26963.4]
  assign x364_1_clock = clock; // @[:@26971.4]
  assign x364_1_io_a = x258_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@26973.4]
  assign x364_1_io_b = 32'h2; // @[Math.scala 264:17:@26974.4]
  assign x364_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26975.4]
  assign x365_1_clock = clock; // @[:@26983.4]
  assign x365_1_io_a = x258_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@26985.4]
  assign x365_1_io_b = 32'h1; // @[Math.scala 264:17:@26986.4]
  assign x365_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@26987.4]
  assign x366_x3_1_clock = clock; // @[:@26993.4]
  assign x366_x3_1_reset = reset; // @[:@26994.4]
  assign x366_x3_1_io_a = x357_1_io_result; // @[Math.scala 151:17:@26995.4]
  assign x366_x3_1_io_b = x358_1_io_result; // @[Math.scala 152:17:@26996.4]
  assign x366_x3_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@26997.4]
  assign x367_x4_1_clock = clock; // @[:@27003.4]
  assign x367_x4_1_reset = reset; // @[:@27004.4]
  assign x367_x4_1_io_a = x359_1_io_result; // @[Math.scala 151:17:@27005.4]
  assign x367_x4_1_io_b = x360_1_io_result; // @[Math.scala 152:17:@27006.4]
  assign x367_x4_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27007.4]
  assign x368_x3_1_clock = clock; // @[:@27013.4]
  assign x368_x3_1_reset = reset; // @[:@27014.4]
  assign x368_x3_1_io_a = x361_1_io_result; // @[Math.scala 151:17:@27015.4]
  assign x368_x3_1_io_b = x362_1_io_result; // @[Math.scala 152:17:@27016.4]
  assign x368_x3_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27017.4]
  assign x369_x4_1_clock = clock; // @[:@27023.4]
  assign x369_x4_1_reset = reset; // @[:@27024.4]
  assign x369_x4_1_io_a = x363_1_io_result; // @[Math.scala 151:17:@27025.4]
  assign x369_x4_1_io_b = x364_1_io_result; // @[Math.scala 152:17:@27026.4]
  assign x369_x4_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27027.4]
  assign x370_x3_1_clock = clock; // @[:@27033.4]
  assign x370_x3_1_reset = reset; // @[:@27034.4]
  assign x370_x3_1_io_a = x366_x3_1_io_result; // @[Math.scala 151:17:@27035.4]
  assign x370_x3_1_io_b = x367_x4_1_io_result; // @[Math.scala 152:17:@27036.4]
  assign x370_x3_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27037.4]
  assign x371_x4_1_clock = clock; // @[:@27043.4]
  assign x371_x4_1_reset = reset; // @[:@27044.4]
  assign x371_x4_1_io_a = x368_x3_1_io_result; // @[Math.scala 151:17:@27045.4]
  assign x371_x4_1_io_b = x369_x4_1_io_result; // @[Math.scala 152:17:@27046.4]
  assign x371_x4_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27047.4]
  assign x372_x3_1_clock = clock; // @[:@27053.4]
  assign x372_x3_1_reset = reset; // @[:@27054.4]
  assign x372_x3_1_io_a = x370_x3_1_io_result; // @[Math.scala 151:17:@27055.4]
  assign x372_x3_1_io_b = x371_x4_1_io_result; // @[Math.scala 152:17:@27056.4]
  assign x372_x3_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27057.4]
  assign RetimeWrapper_60_clock = clock; // @[:@27063.4]
  assign RetimeWrapper_60_reset = reset; // @[:@27064.4]
  assign RetimeWrapper_60_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27066.4]
  assign RetimeWrapper_60_io_in = x365_1_io_result; // @[package.scala 94:16:@27065.4]
  assign x373_sum_1_clock = clock; // @[:@27072.4]
  assign x373_sum_1_reset = reset; // @[:@27073.4]
  assign x373_sum_1_io_a = x372_x3_1_io_result; // @[Math.scala 151:17:@27074.4]
  assign x373_sum_1_io_b = RetimeWrapper_60_io_out; // @[Math.scala 152:17:@27075.4]
  assign x373_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27076.4]
  assign x374_1_io_b = x373_sum_1_io_result; // @[Math.scala 721:17:@27084.4]
  assign x375_mul_1_clock = clock; // @[:@27093.4]
  assign x375_mul_1_io_a = x374_1_io_result; // @[Math.scala 263:17:@27095.4]
  assign x375_mul_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27097.4]
  assign x376_1_io_b = x375_mul_1_io_result; // @[Math.scala 721:17:@27105.4]
  assign x377_1_clock = clock; // @[:@27114.4]
  assign x377_1_io_a = x258_lb_0_io_rPort_4_output_0; // @[Math.scala 263:17:@27116.4]
  assign x377_1_io_b = 32'h1; // @[Math.scala 264:17:@27117.4]
  assign x377_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27118.4]
  assign x378_1_clock = clock; // @[:@27126.4]
  assign x378_1_io_a = x258_lb_0_io_rPort_11_output_0; // @[Math.scala 263:17:@27128.4]
  assign x378_1_io_b = 32'h2; // @[Math.scala 264:17:@27129.4]
  assign x378_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27130.4]
  assign x379_1_clock = clock; // @[:@27138.4]
  assign x379_1_io_a = x258_lb_0_io_rPort_6_output_0; // @[Math.scala 263:17:@27140.4]
  assign x379_1_io_b = 32'h1; // @[Math.scala 264:17:@27141.4]
  assign x379_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27142.4]
  assign x380_1_clock = clock; // @[:@27150.4]
  assign x380_1_io_a = x258_lb_0_io_rPort_10_output_0; // @[Math.scala 263:17:@27152.4]
  assign x380_1_io_b = 32'h2; // @[Math.scala 264:17:@27153.4]
  assign x380_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27154.4]
  assign x381_1_clock = clock; // @[:@27162.4]
  assign x381_1_io_a = x258_lb_0_io_rPort_3_output_0; // @[Math.scala 263:17:@27164.4]
  assign x381_1_io_b = 32'h4; // @[Math.scala 264:17:@27165.4]
  assign x381_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27166.4]
  assign x382_1_clock = clock; // @[:@27174.4]
  assign x382_1_io_a = x258_lb_0_io_rPort_2_output_0; // @[Math.scala 263:17:@27176.4]
  assign x382_1_io_b = 32'h2; // @[Math.scala 264:17:@27177.4]
  assign x382_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27178.4]
  assign x383_1_clock = clock; // @[:@27186.4]
  assign x383_1_io_a = x258_lb_0_io_rPort_7_output_0; // @[Math.scala 263:17:@27188.4]
  assign x383_1_io_b = 32'h1; // @[Math.scala 264:17:@27189.4]
  assign x383_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27190.4]
  assign x384_1_clock = clock; // @[:@27198.4]
  assign x384_1_io_a = x258_lb_0_io_rPort_5_output_0; // @[Math.scala 263:17:@27200.4]
  assign x384_1_io_b = 32'h2; // @[Math.scala 264:17:@27201.4]
  assign x384_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27202.4]
  assign x385_1_clock = clock; // @[:@27210.4]
  assign x385_1_io_a = x258_lb_0_io_rPort_8_output_0; // @[Math.scala 263:17:@27212.4]
  assign x385_1_io_b = 32'h1; // @[Math.scala 264:17:@27213.4]
  assign x385_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27214.4]
  assign x386_x3_1_clock = clock; // @[:@27220.4]
  assign x386_x3_1_reset = reset; // @[:@27221.4]
  assign x386_x3_1_io_a = x377_1_io_result; // @[Math.scala 151:17:@27222.4]
  assign x386_x3_1_io_b = x378_1_io_result; // @[Math.scala 152:17:@27223.4]
  assign x386_x3_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27224.4]
  assign x387_x4_1_clock = clock; // @[:@27230.4]
  assign x387_x4_1_reset = reset; // @[:@27231.4]
  assign x387_x4_1_io_a = x379_1_io_result; // @[Math.scala 151:17:@27232.4]
  assign x387_x4_1_io_b = x380_1_io_result; // @[Math.scala 152:17:@27233.4]
  assign x387_x4_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27234.4]
  assign x388_x3_1_clock = clock; // @[:@27240.4]
  assign x388_x3_1_reset = reset; // @[:@27241.4]
  assign x388_x3_1_io_a = x381_1_io_result; // @[Math.scala 151:17:@27242.4]
  assign x388_x3_1_io_b = x382_1_io_result; // @[Math.scala 152:17:@27243.4]
  assign x388_x3_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27244.4]
  assign x389_x4_1_clock = clock; // @[:@27250.4]
  assign x389_x4_1_reset = reset; // @[:@27251.4]
  assign x389_x4_1_io_a = x383_1_io_result; // @[Math.scala 151:17:@27252.4]
  assign x389_x4_1_io_b = x384_1_io_result; // @[Math.scala 152:17:@27253.4]
  assign x389_x4_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27254.4]
  assign x390_x3_1_clock = clock; // @[:@27260.4]
  assign x390_x3_1_reset = reset; // @[:@27261.4]
  assign x390_x3_1_io_a = x386_x3_1_io_result; // @[Math.scala 151:17:@27262.4]
  assign x390_x3_1_io_b = x387_x4_1_io_result; // @[Math.scala 152:17:@27263.4]
  assign x390_x3_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27264.4]
  assign x391_x4_1_clock = clock; // @[:@27270.4]
  assign x391_x4_1_reset = reset; // @[:@27271.4]
  assign x391_x4_1_io_a = x388_x3_1_io_result; // @[Math.scala 151:17:@27272.4]
  assign x391_x4_1_io_b = x389_x4_1_io_result; // @[Math.scala 152:17:@27273.4]
  assign x391_x4_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27274.4]
  assign x392_x3_1_clock = clock; // @[:@27280.4]
  assign x392_x3_1_reset = reset; // @[:@27281.4]
  assign x392_x3_1_io_a = x390_x3_1_io_result; // @[Math.scala 151:17:@27282.4]
  assign x392_x3_1_io_b = x391_x4_1_io_result; // @[Math.scala 152:17:@27283.4]
  assign x392_x3_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27284.4]
  assign RetimeWrapper_61_clock = clock; // @[:@27290.4]
  assign RetimeWrapper_61_reset = reset; // @[:@27291.4]
  assign RetimeWrapper_61_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27293.4]
  assign RetimeWrapper_61_io_in = x385_1_io_result; // @[package.scala 94:16:@27292.4]
  assign x393_sum_1_clock = clock; // @[:@27299.4]
  assign x393_sum_1_reset = reset; // @[:@27300.4]
  assign x393_sum_1_io_a = x392_x3_1_io_result; // @[Math.scala 151:17:@27301.4]
  assign x393_sum_1_io_b = RetimeWrapper_61_io_out; // @[Math.scala 152:17:@27302.4]
  assign x393_sum_1_io_flow = io_in_x222_TREADY; // @[Math.scala 153:20:@27303.4]
  assign x394_1_io_b = x393_sum_1_io_result; // @[Math.scala 721:17:@27311.4]
  assign x395_mul_1_clock = clock; // @[:@27320.4]
  assign x395_mul_1_io_a = x394_1_io_result; // @[Math.scala 263:17:@27322.4]
  assign x395_mul_1_io_flow = io_in_x222_TREADY; // @[Math.scala 265:20:@27324.4]
  assign x396_1_io_b = x395_mul_1_io_result; // @[Math.scala 721:17:@27332.4]
  assign RetimeWrapper_62_clock = clock; // @[:@27345.4]
  assign RetimeWrapper_62_reset = reset; // @[:@27346.4]
  assign RetimeWrapper_62_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27348.4]
  assign RetimeWrapper_62_io_in = {x376_number,x396_number}; // @[package.scala 94:16:@27347.4]
  assign RetimeWrapper_63_clock = clock; // @[:@27354.4]
  assign RetimeWrapper_63_reset = reset; // @[:@27355.4]
  assign RetimeWrapper_63_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27357.4]
  assign RetimeWrapper_63_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@27356.4]
  assign RetimeWrapper_64_clock = clock; // @[:@27363.4]
  assign RetimeWrapper_64_reset = reset; // @[:@27364.4]
  assign RetimeWrapper_64_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27366.4]
  assign RetimeWrapper_64_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_1; // @[package.scala 94:16:@27365.4]
  assign RetimeWrapper_65_clock = clock; // @[:@27372.4]
  assign RetimeWrapper_65_reset = reset; // @[:@27373.4]
  assign RetimeWrapper_65_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@27375.4]
  assign RetimeWrapper_65_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@27374.4]
endmodule
module x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1( // @[:@27393.2]
  input          clock, // @[:@27394.4]
  input          reset, // @[:@27395.4]
  input          io_in_x221_TVALID, // @[:@27396.4]
  output         io_in_x221_TREADY, // @[:@27396.4]
  input  [255:0] io_in_x221_TDATA, // @[:@27396.4]
  input  [7:0]   io_in_x221_TID, // @[:@27396.4]
  input  [7:0]   io_in_x221_TDEST, // @[:@27396.4]
  output         io_in_x222_TVALID, // @[:@27396.4]
  input          io_in_x222_TREADY, // @[:@27396.4]
  output [255:0] io_in_x222_TDATA, // @[:@27396.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@27396.4]
  input          io_sigsIn_smChildAcks_0, // @[:@27396.4]
  output         io_sigsOut_smDoneIn_0, // @[:@27396.4]
  input          io_rr // @[:@27396.4]
);
  wire  x251_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire  x251_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire  x251_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire  x251_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire [12:0] x251_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire [12:0] x251_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire  x251_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire  x251_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire  x251_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@27430.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_clock; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_reset; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_enable; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_parentAck; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_backpressure; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@27518.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@27518.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@27518.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@27518.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@27518.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@27560.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@27560.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@27560.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@27560.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@27560.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@27568.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@27568.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@27568.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@27568.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@27568.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_clock; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_reset; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TREADY; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire [255:0] x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TDATA; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire [7:0] x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TID; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire [7:0] x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TDEST; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TVALID; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TREADY; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire [255:0] x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TDATA; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire [31:0] x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire [31:0] x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_rr; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
  wire  _T_240; // @[package.scala 96:25:@27523.4 package.scala 96:25:@27524.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[sm_x402_outr_UnitPipe.scala 69:66:@27529.4]
  wire  _T_253; // @[package.scala 96:25:@27565.4 package.scala 96:25:@27566.4]
  wire  _T_259; // @[package.scala 96:25:@27573.4 package.scala 96:25:@27574.4]
  wire  _T_262; // @[SpatialBlocks.scala 138:93:@27576.4]
  wire  x401_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@27577.4]
  wire  _T_264; // @[SpatialBlocks.scala 157:36:@27585.4]
  wire  _T_265; // @[SpatialBlocks.scala 157:78:@27586.4]
  wire  _T_272; // @[SpatialBlocks.scala 159:58:@27598.4]
  x229_ctrchain x251_ctrchain ( // @[SpatialBlocks.scala 37:22:@27430.4]
    .clock(x251_ctrchain_clock),
    .reset(x251_ctrchain_reset),
    .io_input_reset(x251_ctrchain_io_input_reset),
    .io_input_enable(x251_ctrchain_io_input_enable),
    .io_output_counts_1(x251_ctrchain_io_output_counts_1),
    .io_output_counts_0(x251_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x251_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x251_ctrchain_io_output_oobs_1),
    .io_output_done(x251_ctrchain_io_output_done)
  );
  x401_inr_Foreach_SAMPLER_BOX_sm x401_inr_Foreach_SAMPLER_BOX_sm ( // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 32:18:@27490.4]
    .clock(x401_inr_Foreach_SAMPLER_BOX_sm_clock),
    .reset(x401_inr_Foreach_SAMPLER_BOX_sm_reset),
    .io_enable(x401_inr_Foreach_SAMPLER_BOX_sm_io_enable),
    .io_done(x401_inr_Foreach_SAMPLER_BOX_sm_io_done),
    .io_doneLatch(x401_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch),
    .io_ctrDone(x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone),
    .io_datapathEn(x401_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn),
    .io_ctrInc(x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc),
    .io_ctrRst(x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst),
    .io_parentAck(x401_inr_Foreach_SAMPLER_BOX_sm_io_parentAck),
    .io_backpressure(x401_inr_Foreach_SAMPLER_BOX_sm_io_backpressure),
    .io_break(x401_inr_Foreach_SAMPLER_BOX_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@27518.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@27560.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@27568.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1 x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1 ( // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 552:24:@27602.4]
    .clock(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_clock),
    .reset(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_reset),
    .io_in_x221_TREADY(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TREADY),
    .io_in_x221_TDATA(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TDATA),
    .io_in_x221_TID(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TID),
    .io_in_x221_TDEST(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TDEST),
    .io_in_x222_TVALID(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TVALID),
    .io_in_x222_TREADY(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TREADY),
    .io_in_x222_TDATA(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TDATA),
    .io_sigsIn_backpressure(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_rr)
  );
  assign _T_240 = RetimeWrapper_io_out; // @[package.scala 96:25:@27523.4 package.scala 96:25:@27524.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure = io_in_x221_TVALID | x401_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x402_outr_UnitPipe.scala 69:66:@27529.4]
  assign _T_253 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@27565.4 package.scala 96:25:@27566.4]
  assign _T_259 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@27573.4 package.scala 96:25:@27574.4]
  assign _T_262 = ~ _T_259; // @[SpatialBlocks.scala 138:93:@27576.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn = _T_253 & _T_262; // @[SpatialBlocks.scala 138:90:@27577.4]
  assign _T_264 = x401_inr_Foreach_SAMPLER_BOX_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@27585.4]
  assign _T_265 = ~ x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@27586.4]
  assign _T_272 = x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrInc; // @[SpatialBlocks.scala 159:58:@27598.4]
  assign io_in_x221_TREADY = x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TREADY; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 48:23:@27660.4]
  assign io_in_x222_TVALID = x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TVALID; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 49:23:@27670.4]
  assign io_in_x222_TDATA = x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TDATA; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 49:23:@27668.4]
  assign io_sigsOut_smDoneIn_0 = x401_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[SpatialBlocks.scala 156:53:@27583.4]
  assign x251_ctrchain_clock = clock; // @[:@27431.4]
  assign x251_ctrchain_reset = reset; // @[:@27432.4]
  assign x251_ctrchain_io_input_reset = x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@27601.4]
  assign x251_ctrchain_io_input_enable = _T_272 & x401_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 132:75:@27553.4 SpatialBlocks.scala 159:42:@27600.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sm_clock = clock; // @[:@27491.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sm_reset = reset; // @[:@27492.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sm_io_enable = x401_inr_Foreach_SAMPLER_BOX_sigsIn_baseEn & x401_inr_Foreach_SAMPLER_BOX_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@27580.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sm_io_ctrDone = io_rr ? _T_240 : 1'h0; // @[sm_x402_outr_UnitPipe.scala 67:50:@27526.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@27582.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sm_io_backpressure = io_in_x222_TREADY | x401_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@27554.4]
  assign x401_inr_Foreach_SAMPLER_BOX_sm_io_break = 1'h0; // @[sm_x402_outr_UnitPipe.scala 71:48:@27532.4]
  assign RetimeWrapper_clock = clock; // @[:@27519.4]
  assign RetimeWrapper_reset = reset; // @[:@27520.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@27522.4]
  assign RetimeWrapper_io_in = x251_ctrchain_io_output_done; // @[package.scala 94:16:@27521.4]
  assign RetimeWrapper_1_clock = clock; // @[:@27561.4]
  assign RetimeWrapper_1_reset = reset; // @[:@27562.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@27564.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@27563.4]
  assign RetimeWrapper_2_clock = clock; // @[:@27569.4]
  assign RetimeWrapper_2_reset = reset; // @[:@27570.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@27572.4]
  assign RetimeWrapper_2_io_in = x401_inr_Foreach_SAMPLER_BOX_sm_io_done; // @[package.scala 94:16:@27571.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_clock = clock; // @[:@27603.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_reset = reset; // @[:@27604.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TDATA = io_in_x221_TDATA; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 48:23:@27659.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TID = io_in_x221_TID; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 48:23:@27655.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x221_TDEST = io_in_x221_TDEST; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 48:23:@27654.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_in_x222_TREADY = io_in_x222_TREADY; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 49:23:@27669.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_backpressure = io_in_x222_TREADY | x401_inr_Foreach_SAMPLER_BOX_sm_io_doneLatch; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 557:22:@27687.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_datapathEn = _T_264 & _T_265; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 557:22:@27685.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_break = x401_inr_Foreach_SAMPLER_BOX_sm_io_break; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 557:22:@27683.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x251_ctrchain_io_output_counts_1[12]}},x251_ctrchain_io_output_counts_1}; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 557:22:@27678.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x251_ctrchain_io_output_counts_0[12]}},x251_ctrchain_io_output_counts_0}; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 557:22:@27677.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x251_ctrchain_io_output_oobs_0; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 557:22:@27675.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x251_ctrchain_io_output_oobs_1; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 557:22:@27676.4]
  assign x401_inr_Foreach_SAMPLER_BOX_kernelx401_inr_Foreach_SAMPLER_BOX_concrete1_io_rr = io_rr; // @[sm_x401_inr_Foreach_SAMPLER_BOX.scala 556:18:@27671.4]
endmodule
module x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1( // @[:@27701.2]
  input          clock, // @[:@27702.4]
  input          reset, // @[:@27703.4]
  input          io_in_x221_TVALID, // @[:@27704.4]
  output         io_in_x221_TREADY, // @[:@27704.4]
  input  [255:0] io_in_x221_TDATA, // @[:@27704.4]
  input  [7:0]   io_in_x221_TID, // @[:@27704.4]
  input  [7:0]   io_in_x221_TDEST, // @[:@27704.4]
  output         io_in_x222_TVALID, // @[:@27704.4]
  input          io_in_x222_TREADY, // @[:@27704.4]
  output [255:0] io_in_x222_TDATA, // @[:@27704.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@27704.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@27704.4]
  input          io_sigsIn_smChildAcks_0, // @[:@27704.4]
  input          io_sigsIn_smChildAcks_1, // @[:@27704.4]
  output         io_sigsOut_smDoneIn_0, // @[:@27704.4]
  output         io_sigsOut_smDoneIn_1, // @[:@27704.4]
  output         io_sigsOut_smCtrCopyDone_0, // @[:@27704.4]
  output         io_sigsOut_smCtrCopyDone_1, // @[:@27704.4]
  input          io_rr // @[:@27704.4]
);
  wire  x224_fifoinraw_0_clock; // @[m_x224_fifoinraw_0.scala 27:17:@27718.4]
  wire  x224_fifoinraw_0_reset; // @[m_x224_fifoinraw_0.scala 27:17:@27718.4]
  wire  x225_fifoinpacked_0_clock; // @[m_x225_fifoinpacked_0.scala 27:17:@27742.4]
  wire  x225_fifoinpacked_0_reset; // @[m_x225_fifoinpacked_0.scala 27:17:@27742.4]
  wire  x225_fifoinpacked_0_io_wPort_0_en_0; // @[m_x225_fifoinpacked_0.scala 27:17:@27742.4]
  wire  x225_fifoinpacked_0_io_full; // @[m_x225_fifoinpacked_0.scala 27:17:@27742.4]
  wire  x225_fifoinpacked_0_io_active_0_in; // @[m_x225_fifoinpacked_0.scala 27:17:@27742.4]
  wire  x225_fifoinpacked_0_io_active_0_out; // @[m_x225_fifoinpacked_0.scala 27:17:@27742.4]
  wire  x226_fifooutraw_0_clock; // @[m_x226_fifooutraw_0.scala 27:17:@27766.4]
  wire  x226_fifooutraw_0_reset; // @[m_x226_fifooutraw_0.scala 27:17:@27766.4]
  wire  x229_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire  x229_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire  x229_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire  x229_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire [12:0] x229_ctrchain_io_output_counts_1; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire [12:0] x229_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire  x229_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire  x229_ctrchain_io_output_oobs_1; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire  x229_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@27790.4]
  wire  x247_inr_Foreach_sm_clock; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_reset; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_enable; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_done; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_doneLatch; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_ctrDone; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_datapathEn; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_ctrInc; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_ctrRst; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_parentAck; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_backpressure; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  x247_inr_Foreach_sm_io_break; // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@27878.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@27878.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@27878.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@27878.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@27878.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@27924.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@27924.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@27924.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@27924.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@27924.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@27932.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@27932.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@27932.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@27932.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@27932.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_clock; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_reset; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_wPort_0_en_0; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_full; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_active_0_in; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_active_0_out; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire [31:0] x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire [31:0] x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_rr; // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
  wire  x402_outr_UnitPipe_sm_clock; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_reset; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_enable; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_done; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_rst; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_ctrDone; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_ctrInc; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_parentAck; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  x402_outr_UnitPipe_sm_io_childAck_0; // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@28156.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@28156.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@28156.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@28156.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@28156.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@28164.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@28164.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@28164.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@28164.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@28164.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_clock; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_reset; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TVALID; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TREADY; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire [255:0] x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TDATA; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire [7:0] x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TID; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire [7:0] x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TDEST; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TVALID; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TREADY; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire [255:0] x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TDATA; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_rr; // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
  wire  _T_254; // @[package.scala 96:25:@27883.4 package.scala 96:25:@27884.4]
  wire  _T_260; // @[implicits.scala 47:10:@27887.4]
  wire  _T_261; // @[sm_x403_outr_UnitPipe.scala 70:41:@27888.4]
  wire  _T_262; // @[sm_x403_outr_UnitPipe.scala 70:78:@27889.4]
  wire  _T_263; // @[sm_x403_outr_UnitPipe.scala 70:76:@27890.4]
  wire  _T_275; // @[package.scala 96:25:@27929.4 package.scala 96:25:@27930.4]
  wire  _T_281; // @[package.scala 96:25:@27937.4 package.scala 96:25:@27938.4]
  wire  _T_284; // @[SpatialBlocks.scala 138:93:@27940.4]
  wire  _T_286; // @[SpatialBlocks.scala 157:36:@27949.4]
  wire  _T_287; // @[SpatialBlocks.scala 157:78:@27950.4]
  wire  _T_354; // @[package.scala 100:49:@28127.4]
  reg  _T_357; // @[package.scala 48:56:@28128.4]
  reg [31:0] _RAND_0;
  wire  _T_371; // @[package.scala 96:25:@28161.4 package.scala 96:25:@28162.4]
  wire  _T_377; // @[package.scala 96:25:@28169.4 package.scala 96:25:@28170.4]
  wire  _T_380; // @[SpatialBlocks.scala 138:93:@28172.4]
  x224_fifoinraw_0 x224_fifoinraw_0 ( // @[m_x224_fifoinraw_0.scala 27:17:@27718.4]
    .clock(x224_fifoinraw_0_clock),
    .reset(x224_fifoinraw_0_reset)
  );
  x225_fifoinpacked_0 x225_fifoinpacked_0 ( // @[m_x225_fifoinpacked_0.scala 27:17:@27742.4]
    .clock(x225_fifoinpacked_0_clock),
    .reset(x225_fifoinpacked_0_reset),
    .io_wPort_0_en_0(x225_fifoinpacked_0_io_wPort_0_en_0),
    .io_full(x225_fifoinpacked_0_io_full),
    .io_active_0_in(x225_fifoinpacked_0_io_active_0_in),
    .io_active_0_out(x225_fifoinpacked_0_io_active_0_out)
  );
  x224_fifoinraw_0 x226_fifooutraw_0 ( // @[m_x226_fifooutraw_0.scala 27:17:@27766.4]
    .clock(x226_fifooutraw_0_clock),
    .reset(x226_fifooutraw_0_reset)
  );
  x229_ctrchain x229_ctrchain ( // @[SpatialBlocks.scala 37:22:@27790.4]
    .clock(x229_ctrchain_clock),
    .reset(x229_ctrchain_reset),
    .io_input_reset(x229_ctrchain_io_input_reset),
    .io_input_enable(x229_ctrchain_io_input_enable),
    .io_output_counts_1(x229_ctrchain_io_output_counts_1),
    .io_output_counts_0(x229_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x229_ctrchain_io_output_oobs_0),
    .io_output_oobs_1(x229_ctrchain_io_output_oobs_1),
    .io_output_done(x229_ctrchain_io_output_done)
  );
  x247_inr_Foreach_sm x247_inr_Foreach_sm ( // @[sm_x247_inr_Foreach.scala 32:18:@27850.4]
    .clock(x247_inr_Foreach_sm_clock),
    .reset(x247_inr_Foreach_sm_reset),
    .io_enable(x247_inr_Foreach_sm_io_enable),
    .io_done(x247_inr_Foreach_sm_io_done),
    .io_doneLatch(x247_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x247_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x247_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x247_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x247_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x247_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x247_inr_Foreach_sm_io_backpressure),
    .io_break(x247_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@27878.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@27924.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@27932.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  x247_inr_Foreach_kernelx247_inr_Foreach_concrete1 x247_inr_Foreach_kernelx247_inr_Foreach_concrete1 ( // @[sm_x247_inr_Foreach.scala 106:24:@27967.4]
    .clock(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_clock),
    .reset(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_reset),
    .io_in_x225_fifoinpacked_0_wPort_0_en_0(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_wPort_0_en_0),
    .io_in_x225_fifoinpacked_0_full(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_full),
    .io_in_x225_fifoinpacked_0_active_0_in(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_active_0_in),
    .io_in_x225_fifoinpacked_0_active_0_out(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_active_0_out),
    .io_sigsIn_backpressure(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_1(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1),
    .io_sigsIn_cchainOutputs_0_counts_0(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_sigsIn_cchainOutputs_0_oobs_1(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1),
    .io_rr(x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_rr)
  );
  RootController_sm x402_outr_UnitPipe_sm ( // @[sm_x402_outr_UnitPipe.scala 32:18:@28099.4]
    .clock(x402_outr_UnitPipe_sm_clock),
    .reset(x402_outr_UnitPipe_sm_reset),
    .io_enable(x402_outr_UnitPipe_sm_io_enable),
    .io_done(x402_outr_UnitPipe_sm_io_done),
    .io_rst(x402_outr_UnitPipe_sm_io_rst),
    .io_ctrDone(x402_outr_UnitPipe_sm_io_ctrDone),
    .io_ctrInc(x402_outr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x402_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x402_outr_UnitPipe_sm_io_doneIn_0),
    .io_enableOut_0(x402_outr_UnitPipe_sm_io_enableOut_0),
    .io_childAck_0(x402_outr_UnitPipe_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@28156.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@28164.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1 x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1 ( // @[sm_x402_outr_UnitPipe.scala 76:24:@28194.4]
    .clock(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_clock),
    .reset(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_reset),
    .io_in_x221_TVALID(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TVALID),
    .io_in_x221_TREADY(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TREADY),
    .io_in_x221_TDATA(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TDATA),
    .io_in_x221_TID(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TID),
    .io_in_x221_TDEST(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TDEST),
    .io_in_x222_TVALID(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TVALID),
    .io_in_x222_TREADY(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TREADY),
    .io_in_x222_TDATA(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TDATA),
    .io_sigsIn_smEnableOuts_0(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_254 = RetimeWrapper_io_out; // @[package.scala 96:25:@27883.4 package.scala 96:25:@27884.4]
  assign _T_260 = x225_fifoinpacked_0_io_full; // @[implicits.scala 47:10:@27887.4]
  assign _T_261 = ~ _T_260; // @[sm_x403_outr_UnitPipe.scala 70:41:@27888.4]
  assign _T_262 = ~ x225_fifoinpacked_0_io_active_0_out; // @[sm_x403_outr_UnitPipe.scala 70:78:@27889.4]
  assign _T_263 = _T_261 | _T_262; // @[sm_x403_outr_UnitPipe.scala 70:76:@27890.4]
  assign _T_275 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@27929.4 package.scala 96:25:@27930.4]
  assign _T_281 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@27937.4 package.scala 96:25:@27938.4]
  assign _T_284 = ~ _T_281; // @[SpatialBlocks.scala 138:93:@27940.4]
  assign _T_286 = x247_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@27949.4]
  assign _T_287 = ~ x247_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@27950.4]
  assign _T_354 = x402_outr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@28127.4]
  assign _T_371 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@28161.4 package.scala 96:25:@28162.4]
  assign _T_377 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@28169.4 package.scala 96:25:@28170.4]
  assign _T_380 = ~ _T_377; // @[SpatialBlocks.scala 138:93:@28172.4]
  assign io_in_x221_TREADY = x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TREADY; // @[sm_x402_outr_UnitPipe.scala 48:23:@28250.4]
  assign io_in_x222_TVALID = x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TVALID; // @[sm_x402_outr_UnitPipe.scala 49:23:@28260.4]
  assign io_in_x222_TDATA = x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TDATA; // @[sm_x402_outr_UnitPipe.scala 49:23:@28258.4]
  assign io_sigsOut_smDoneIn_0 = x247_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@27947.4]
  assign io_sigsOut_smDoneIn_1 = x402_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@28179.4]
  assign io_sigsOut_smCtrCopyDone_0 = x247_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@27966.4]
  assign io_sigsOut_smCtrCopyDone_1 = x402_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@28193.4]
  assign x224_fifoinraw_0_clock = clock; // @[:@27719.4]
  assign x224_fifoinraw_0_reset = reset; // @[:@27720.4]
  assign x225_fifoinpacked_0_clock = clock; // @[:@27743.4]
  assign x225_fifoinpacked_0_reset = reset; // @[:@27744.4]
  assign x225_fifoinpacked_0_io_wPort_0_en_0 = x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_wPort_0_en_0; // @[MemInterfaceType.scala 67:44:@28027.4]
  assign x225_fifoinpacked_0_io_active_0_in = x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_active_0_in; // @[MemInterfaceType.scala 167:86:@28026.4]
  assign x226_fifooutraw_0_clock = clock; // @[:@27767.4]
  assign x226_fifooutraw_0_reset = reset; // @[:@27768.4]
  assign x229_ctrchain_clock = clock; // @[:@27791.4]
  assign x229_ctrchain_reset = reset; // @[:@27792.4]
  assign x229_ctrchain_io_input_reset = x247_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@27965.4]
  assign x229_ctrchain_io_input_enable = x247_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@27917.4 SpatialBlocks.scala 159:42:@27964.4]
  assign x247_inr_Foreach_sm_clock = clock; // @[:@27851.4]
  assign x247_inr_Foreach_sm_reset = reset; // @[:@27852.4]
  assign x247_inr_Foreach_sm_io_enable = _T_275 & _T_284; // @[SpatialBlocks.scala 140:18:@27944.4]
  assign x247_inr_Foreach_sm_io_ctrDone = io_rr ? _T_254 : 1'h0; // @[sm_x403_outr_UnitPipe.scala 69:38:@27886.4]
  assign x247_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@27946.4]
  assign x247_inr_Foreach_sm_io_backpressure = _T_263 | x247_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@27918.4]
  assign x247_inr_Foreach_sm_io_break = 1'h0; // @[sm_x403_outr_UnitPipe.scala 73:36:@27896.4]
  assign RetimeWrapper_clock = clock; // @[:@27879.4]
  assign RetimeWrapper_reset = reset; // @[:@27880.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@27882.4]
  assign RetimeWrapper_io_in = x229_ctrchain_io_output_done; // @[package.scala 94:16:@27881.4]
  assign RetimeWrapper_1_clock = clock; // @[:@27925.4]
  assign RetimeWrapper_1_reset = reset; // @[:@27926.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@27928.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@27927.4]
  assign RetimeWrapper_2_clock = clock; // @[:@27933.4]
  assign RetimeWrapper_2_reset = reset; // @[:@27934.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@27936.4]
  assign RetimeWrapper_2_io_in = x247_inr_Foreach_sm_io_done; // @[package.scala 94:16:@27935.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_clock = clock; // @[:@27968.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_reset = reset; // @[:@27969.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_full = x225_fifoinpacked_0_io_full; // @[MemInterfaceType.scala 159:15:@28021.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_in_x225_fifoinpacked_0_active_0_out = x225_fifoinpacked_0_io_active_0_out; // @[MemInterfaceType.scala 158:75:@28020.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_backpressure = _T_263 | x247_inr_Foreach_sm_io_doneLatch; // @[sm_x247_inr_Foreach.scala 111:22:@28050.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_286 & _T_287; // @[sm_x247_inr_Foreach.scala 111:22:@28048.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_break = x247_inr_Foreach_sm_io_break; // @[sm_x247_inr_Foreach.scala 111:22:@28046.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_1 = {{19{x229_ctrchain_io_output_counts_1[12]}},x229_ctrchain_io_output_counts_1}; // @[sm_x247_inr_Foreach.scala 111:22:@28041.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{19{x229_ctrchain_io_output_counts_0[12]}},x229_ctrchain_io_output_counts_0}; // @[sm_x247_inr_Foreach.scala 111:22:@28040.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x229_ctrchain_io_output_oobs_0; // @[sm_x247_inr_Foreach.scala 111:22:@28038.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_1 = x229_ctrchain_io_output_oobs_1; // @[sm_x247_inr_Foreach.scala 111:22:@28039.4]
  assign x247_inr_Foreach_kernelx247_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x247_inr_Foreach.scala 110:18:@28034.4]
  assign x402_outr_UnitPipe_sm_clock = clock; // @[:@28100.4]
  assign x402_outr_UnitPipe_sm_reset = reset; // @[:@28101.4]
  assign x402_outr_UnitPipe_sm_io_enable = _T_371 & _T_380; // @[SpatialBlocks.scala 140:18:@28176.4]
  assign x402_outr_UnitPipe_sm_io_rst = 1'h0; // @[SpatialBlocks.scala 134:15:@28151.4]
  assign x402_outr_UnitPipe_sm_io_ctrDone = x402_outr_UnitPipe_sm_io_ctrInc & _T_357; // @[sm_x403_outr_UnitPipe.scala 78:40:@28131.4]
  assign x402_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@28178.4]
  assign x402_outr_UnitPipe_sm_io_doneIn_0 = x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@28148.4]
  assign RetimeWrapper_3_clock = clock; // @[:@28157.4]
  assign RetimeWrapper_3_reset = reset; // @[:@28158.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@28160.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@28159.4]
  assign RetimeWrapper_4_clock = clock; // @[:@28165.4]
  assign RetimeWrapper_4_reset = reset; // @[:@28166.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@28168.4]
  assign RetimeWrapper_4_io_in = x402_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@28167.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_clock = clock; // @[:@28195.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_reset = reset; // @[:@28196.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TVALID = io_in_x221_TVALID; // @[sm_x402_outr_UnitPipe.scala 48:23:@28251.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TDATA = io_in_x221_TDATA; // @[sm_x402_outr_UnitPipe.scala 48:23:@28249.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TID = io_in_x221_TID; // @[sm_x402_outr_UnitPipe.scala 48:23:@28245.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x221_TDEST = io_in_x221_TDEST; // @[sm_x402_outr_UnitPipe.scala 48:23:@28244.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_in_x222_TREADY = io_in_x222_TREADY; // @[sm_x402_outr_UnitPipe.scala 49:23:@28259.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x402_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x402_outr_UnitPipe.scala 81:22:@28269.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x402_outr_UnitPipe_sm_io_childAck_0; // @[sm_x402_outr_UnitPipe.scala 81:22:@28267.4]
  assign x402_outr_UnitPipe_kernelx402_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x402_outr_UnitPipe.scala 80:18:@28261.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_357 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_357 <= 1'h0;
    end else begin
      _T_357 <= _T_354;
    end
  end
endmodule
module x425_outr_UnitPipe_sm( // @[:@28758.2]
  input   clock, // @[:@28759.4]
  input   reset, // @[:@28760.4]
  input   io_enable, // @[:@28761.4]
  output  io_done, // @[:@28761.4]
  input   io_parentAck, // @[:@28761.4]
  input   io_doneIn_0, // @[:@28761.4]
  input   io_doneIn_1, // @[:@28761.4]
  input   io_doneIn_2, // @[:@28761.4]
  output  io_enableOut_0, // @[:@28761.4]
  output  io_enableOut_1, // @[:@28761.4]
  output  io_enableOut_2, // @[:@28761.4]
  output  io_childAck_0, // @[:@28761.4]
  output  io_childAck_1, // @[:@28761.4]
  output  io_childAck_2, // @[:@28761.4]
  input   io_ctrCopyDone_0, // @[:@28761.4]
  input   io_ctrCopyDone_1, // @[:@28761.4]
  input   io_ctrCopyDone_2 // @[:@28761.4]
);
  wire  active_0_clock; // @[Controllers.scala 76:50:@28764.4]
  wire  active_0_reset; // @[Controllers.scala 76:50:@28764.4]
  wire  active_0_io_input_set; // @[Controllers.scala 76:50:@28764.4]
  wire  active_0_io_input_reset; // @[Controllers.scala 76:50:@28764.4]
  wire  active_0_io_input_asyn_reset; // @[Controllers.scala 76:50:@28764.4]
  wire  active_0_io_output; // @[Controllers.scala 76:50:@28764.4]
  wire  active_1_clock; // @[Controllers.scala 76:50:@28767.4]
  wire  active_1_reset; // @[Controllers.scala 76:50:@28767.4]
  wire  active_1_io_input_set; // @[Controllers.scala 76:50:@28767.4]
  wire  active_1_io_input_reset; // @[Controllers.scala 76:50:@28767.4]
  wire  active_1_io_input_asyn_reset; // @[Controllers.scala 76:50:@28767.4]
  wire  active_1_io_output; // @[Controllers.scala 76:50:@28767.4]
  wire  active_2_clock; // @[Controllers.scala 76:50:@28770.4]
  wire  active_2_reset; // @[Controllers.scala 76:50:@28770.4]
  wire  active_2_io_input_set; // @[Controllers.scala 76:50:@28770.4]
  wire  active_2_io_input_reset; // @[Controllers.scala 76:50:@28770.4]
  wire  active_2_io_input_asyn_reset; // @[Controllers.scala 76:50:@28770.4]
  wire  active_2_io_output; // @[Controllers.scala 76:50:@28770.4]
  wire  done_0_clock; // @[Controllers.scala 77:48:@28773.4]
  wire  done_0_reset; // @[Controllers.scala 77:48:@28773.4]
  wire  done_0_io_input_set; // @[Controllers.scala 77:48:@28773.4]
  wire  done_0_io_input_reset; // @[Controllers.scala 77:48:@28773.4]
  wire  done_0_io_input_asyn_reset; // @[Controllers.scala 77:48:@28773.4]
  wire  done_0_io_output; // @[Controllers.scala 77:48:@28773.4]
  wire  done_1_clock; // @[Controllers.scala 77:48:@28776.4]
  wire  done_1_reset; // @[Controllers.scala 77:48:@28776.4]
  wire  done_1_io_input_set; // @[Controllers.scala 77:48:@28776.4]
  wire  done_1_io_input_reset; // @[Controllers.scala 77:48:@28776.4]
  wire  done_1_io_input_asyn_reset; // @[Controllers.scala 77:48:@28776.4]
  wire  done_1_io_output; // @[Controllers.scala 77:48:@28776.4]
  wire  done_2_clock; // @[Controllers.scala 77:48:@28779.4]
  wire  done_2_reset; // @[Controllers.scala 77:48:@28779.4]
  wire  done_2_io_input_set; // @[Controllers.scala 77:48:@28779.4]
  wire  done_2_io_input_reset; // @[Controllers.scala 77:48:@28779.4]
  wire  done_2_io_input_asyn_reset; // @[Controllers.scala 77:48:@28779.4]
  wire  done_2_io_output; // @[Controllers.scala 77:48:@28779.4]
  wire  iterDone_0_clock; // @[Controllers.scala 90:52:@28820.4]
  wire  iterDone_0_reset; // @[Controllers.scala 90:52:@28820.4]
  wire  iterDone_0_io_input_set; // @[Controllers.scala 90:52:@28820.4]
  wire  iterDone_0_io_input_reset; // @[Controllers.scala 90:52:@28820.4]
  wire  iterDone_0_io_input_asyn_reset; // @[Controllers.scala 90:52:@28820.4]
  wire  iterDone_0_io_output; // @[Controllers.scala 90:52:@28820.4]
  wire  iterDone_1_clock; // @[Controllers.scala 90:52:@28823.4]
  wire  iterDone_1_reset; // @[Controllers.scala 90:52:@28823.4]
  wire  iterDone_1_io_input_set; // @[Controllers.scala 90:52:@28823.4]
  wire  iterDone_1_io_input_reset; // @[Controllers.scala 90:52:@28823.4]
  wire  iterDone_1_io_input_asyn_reset; // @[Controllers.scala 90:52:@28823.4]
  wire  iterDone_1_io_output; // @[Controllers.scala 90:52:@28823.4]
  wire  iterDone_2_clock; // @[Controllers.scala 90:52:@28826.4]
  wire  iterDone_2_reset; // @[Controllers.scala 90:52:@28826.4]
  wire  iterDone_2_io_input_set; // @[Controllers.scala 90:52:@28826.4]
  wire  iterDone_2_io_input_reset; // @[Controllers.scala 90:52:@28826.4]
  wire  iterDone_2_io_input_asyn_reset; // @[Controllers.scala 90:52:@28826.4]
  wire  iterDone_2_io_output; // @[Controllers.scala 90:52:@28826.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@28877.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@28877.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@28877.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@28877.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@28877.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@28891.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@28891.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@28891.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@28891.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@28891.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@28909.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@28909.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@28909.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@28909.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@28909.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@28946.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@28946.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@28946.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@28946.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@28946.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@28960.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@28960.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@28960.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@28960.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@28960.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@28978.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@29015.4]
  wire  RetimeWrapper_7_clock; // @[package.scala 93:22:@29029.4]
  wire  RetimeWrapper_7_reset; // @[package.scala 93:22:@29029.4]
  wire  RetimeWrapper_7_io_flow; // @[package.scala 93:22:@29029.4]
  wire  RetimeWrapper_7_io_in; // @[package.scala 93:22:@29029.4]
  wire  RetimeWrapper_7_io_out; // @[package.scala 93:22:@29029.4]
  wire  RetimeWrapper_8_clock; // @[package.scala 93:22:@29047.4]
  wire  RetimeWrapper_8_reset; // @[package.scala 93:22:@29047.4]
  wire  RetimeWrapper_8_io_flow; // @[package.scala 93:22:@29047.4]
  wire  RetimeWrapper_8_io_in; // @[package.scala 93:22:@29047.4]
  wire  RetimeWrapper_8_io_out; // @[package.scala 93:22:@29047.4]
  wire  RetimeWrapper_9_clock; // @[package.scala 93:22:@29104.4]
  wire  RetimeWrapper_9_reset; // @[package.scala 93:22:@29104.4]
  wire  RetimeWrapper_9_io_flow; // @[package.scala 93:22:@29104.4]
  wire  RetimeWrapper_9_io_in; // @[package.scala 93:22:@29104.4]
  wire  RetimeWrapper_9_io_out; // @[package.scala 93:22:@29104.4]
  wire  RetimeWrapper_10_clock; // @[package.scala 93:22:@29121.4]
  wire  RetimeWrapper_10_reset; // @[package.scala 93:22:@29121.4]
  wire  RetimeWrapper_10_io_flow; // @[package.scala 93:22:@29121.4]
  wire  RetimeWrapper_10_io_in; // @[package.scala 93:22:@29121.4]
  wire  RetimeWrapper_10_io_out; // @[package.scala 93:22:@29121.4]
  wire  _T_77; // @[Controllers.scala 80:47:@28782.4]
  wire  allDone; // @[Controllers.scala 80:47:@28783.4]
  wire  _T_151; // @[Controllers.scala 165:35:@28861.4]
  wire  _T_153; // @[Controllers.scala 165:60:@28862.4]
  wire  _T_154; // @[Controllers.scala 165:58:@28863.4]
  wire  _T_156; // @[Controllers.scala 165:76:@28864.4]
  wire  _T_157; // @[Controllers.scala 165:74:@28865.4]
  wire  _T_161; // @[Controllers.scala 165:109:@28868.4]
  wire  _T_164; // @[Controllers.scala 165:141:@28870.4]
  wire  _T_172; // @[package.scala 96:25:@28882.4 package.scala 96:25:@28883.4]
  wire  _T_176; // @[Controllers.scala 167:54:@28885.4]
  wire  _T_177; // @[Controllers.scala 167:52:@28886.4]
  wire  _T_184; // @[package.scala 96:25:@28896.4 package.scala 96:25:@28897.4]
  wire  _T_202; // @[package.scala 96:25:@28914.4 package.scala 96:25:@28915.4]
  wire  _T_206; // @[Controllers.scala 169:67:@28917.4]
  wire  _T_207; // @[Controllers.scala 169:86:@28918.4]
  wire  _T_219; // @[Controllers.scala 165:35:@28930.4]
  wire  _T_221; // @[Controllers.scala 165:60:@28931.4]
  wire  _T_222; // @[Controllers.scala 165:58:@28932.4]
  wire  _T_224; // @[Controllers.scala 165:76:@28933.4]
  wire  _T_225; // @[Controllers.scala 165:74:@28934.4]
  wire  _T_229; // @[Controllers.scala 165:109:@28937.4]
  wire  _T_232; // @[Controllers.scala 165:141:@28939.4]
  wire  _T_240; // @[package.scala 96:25:@28951.4 package.scala 96:25:@28952.4]
  wire  _T_244; // @[Controllers.scala 167:54:@28954.4]
  wire  _T_245; // @[Controllers.scala 167:52:@28955.4]
  wire  _T_252; // @[package.scala 96:25:@28965.4 package.scala 96:25:@28966.4]
  wire  _T_270; // @[package.scala 96:25:@28983.4 package.scala 96:25:@28984.4]
  wire  _T_274; // @[Controllers.scala 169:67:@28986.4]
  wire  _T_275; // @[Controllers.scala 169:86:@28987.4]
  wire  _T_287; // @[Controllers.scala 165:35:@28999.4]
  wire  _T_289; // @[Controllers.scala 165:60:@29000.4]
  wire  _T_290; // @[Controllers.scala 165:58:@29001.4]
  wire  _T_292; // @[Controllers.scala 165:76:@29002.4]
  wire  _T_293; // @[Controllers.scala 165:74:@29003.4]
  wire  _T_297; // @[Controllers.scala 165:109:@29006.4]
  wire  _T_300; // @[Controllers.scala 165:141:@29008.4]
  wire  _T_308; // @[package.scala 96:25:@29020.4 package.scala 96:25:@29021.4]
  wire  _T_312; // @[Controllers.scala 167:54:@29023.4]
  wire  _T_313; // @[Controllers.scala 167:52:@29024.4]
  wire  _T_320; // @[package.scala 96:25:@29034.4 package.scala 96:25:@29035.4]
  wire  _T_338; // @[package.scala 96:25:@29052.4 package.scala 96:25:@29053.4]
  wire  _T_342; // @[Controllers.scala 169:67:@29055.4]
  wire  _T_343; // @[Controllers.scala 169:86:@29056.4]
  wire  _T_358; // @[Controllers.scala 213:68:@29074.4]
  wire  _T_360; // @[Controllers.scala 213:90:@29076.4]
  wire  _T_362; // @[Controllers.scala 213:132:@29078.4]
  wire  _T_366; // @[Controllers.scala 213:68:@29083.4]
  wire  _T_368; // @[Controllers.scala 213:90:@29085.4]
  wire  _T_374; // @[Controllers.scala 213:68:@29091.4]
  wire  _T_376; // @[Controllers.scala 213:90:@29093.4]
  wire  _T_383; // @[package.scala 100:49:@29099.4]
  reg  _T_386; // @[package.scala 48:56:@29100.4]
  reg [31:0] _RAND_0;
  wire  _T_387; // @[package.scala 100:41:@29102.4]
  reg  _T_400; // @[package.scala 48:56:@29118.4]
  reg [31:0] _RAND_1;
  SRFF active_0 ( // @[Controllers.scala 76:50:@28764.4]
    .clock(active_0_clock),
    .reset(active_0_reset),
    .io_input_set(active_0_io_input_set),
    .io_input_reset(active_0_io_input_reset),
    .io_input_asyn_reset(active_0_io_input_asyn_reset),
    .io_output(active_0_io_output)
  );
  SRFF active_1 ( // @[Controllers.scala 76:50:@28767.4]
    .clock(active_1_clock),
    .reset(active_1_reset),
    .io_input_set(active_1_io_input_set),
    .io_input_reset(active_1_io_input_reset),
    .io_input_asyn_reset(active_1_io_input_asyn_reset),
    .io_output(active_1_io_output)
  );
  SRFF active_2 ( // @[Controllers.scala 76:50:@28770.4]
    .clock(active_2_clock),
    .reset(active_2_reset),
    .io_input_set(active_2_io_input_set),
    .io_input_reset(active_2_io_input_reset),
    .io_input_asyn_reset(active_2_io_input_asyn_reset),
    .io_output(active_2_io_output)
  );
  SRFF done_0 ( // @[Controllers.scala 77:48:@28773.4]
    .clock(done_0_clock),
    .reset(done_0_reset),
    .io_input_set(done_0_io_input_set),
    .io_input_reset(done_0_io_input_reset),
    .io_input_asyn_reset(done_0_io_input_asyn_reset),
    .io_output(done_0_io_output)
  );
  SRFF done_1 ( // @[Controllers.scala 77:48:@28776.4]
    .clock(done_1_clock),
    .reset(done_1_reset),
    .io_input_set(done_1_io_input_set),
    .io_input_reset(done_1_io_input_reset),
    .io_input_asyn_reset(done_1_io_input_asyn_reset),
    .io_output(done_1_io_output)
  );
  SRFF done_2 ( // @[Controllers.scala 77:48:@28779.4]
    .clock(done_2_clock),
    .reset(done_2_reset),
    .io_input_set(done_2_io_input_set),
    .io_input_reset(done_2_io_input_reset),
    .io_input_asyn_reset(done_2_io_input_asyn_reset),
    .io_output(done_2_io_output)
  );
  SRFF iterDone_0 ( // @[Controllers.scala 90:52:@28820.4]
    .clock(iterDone_0_clock),
    .reset(iterDone_0_reset),
    .io_input_set(iterDone_0_io_input_set),
    .io_input_reset(iterDone_0_io_input_reset),
    .io_input_asyn_reset(iterDone_0_io_input_asyn_reset),
    .io_output(iterDone_0_io_output)
  );
  SRFF iterDone_1 ( // @[Controllers.scala 90:52:@28823.4]
    .clock(iterDone_1_clock),
    .reset(iterDone_1_reset),
    .io_input_set(iterDone_1_io_input_set),
    .io_input_reset(iterDone_1_io_input_reset),
    .io_input_asyn_reset(iterDone_1_io_input_asyn_reset),
    .io_output(iterDone_1_io_output)
  );
  SRFF iterDone_2 ( // @[Controllers.scala 90:52:@28826.4]
    .clock(iterDone_2_clock),
    .reset(iterDone_2_reset),
    .io_input_set(iterDone_2_io_input_set),
    .io_input_reset(iterDone_2_io_input_reset),
    .io_input_asyn_reset(iterDone_2_io_input_asyn_reset),
    .io_output(iterDone_2_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@28877.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@28891.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@28909.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@28946.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@28960.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@28978.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@29015.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  RetimeWrapper RetimeWrapper_7 ( // @[package.scala 93:22:@29029.4]
    .clock(RetimeWrapper_7_clock),
    .reset(RetimeWrapper_7_reset),
    .io_flow(RetimeWrapper_7_io_flow),
    .io_in(RetimeWrapper_7_io_in),
    .io_out(RetimeWrapper_7_io_out)
  );
  RetimeWrapper RetimeWrapper_8 ( // @[package.scala 93:22:@29047.4]
    .clock(RetimeWrapper_8_clock),
    .reset(RetimeWrapper_8_reset),
    .io_flow(RetimeWrapper_8_io_flow),
    .io_in(RetimeWrapper_8_io_in),
    .io_out(RetimeWrapper_8_io_out)
  );
  RetimeWrapper RetimeWrapper_9 ( // @[package.scala 93:22:@29104.4]
    .clock(RetimeWrapper_9_clock),
    .reset(RetimeWrapper_9_reset),
    .io_flow(RetimeWrapper_9_io_flow),
    .io_in(RetimeWrapper_9_io_in),
    .io_out(RetimeWrapper_9_io_out)
  );
  RetimeWrapper RetimeWrapper_10 ( // @[package.scala 93:22:@29121.4]
    .clock(RetimeWrapper_10_clock),
    .reset(RetimeWrapper_10_reset),
    .io_flow(RetimeWrapper_10_io_flow),
    .io_in(RetimeWrapper_10_io_in),
    .io_out(RetimeWrapper_10_io_out)
  );
  assign _T_77 = done_0_io_output & done_1_io_output; // @[Controllers.scala 80:47:@28782.4]
  assign allDone = _T_77 & done_2_io_output; // @[Controllers.scala 80:47:@28783.4]
  assign _T_151 = ~ iterDone_0_io_output; // @[Controllers.scala 165:35:@28861.4]
  assign _T_153 = io_doneIn_0 == 1'h0; // @[Controllers.scala 165:60:@28862.4]
  assign _T_154 = _T_151 & _T_153; // @[Controllers.scala 165:58:@28863.4]
  assign _T_156 = done_0_io_output == 1'h0; // @[Controllers.scala 165:76:@28864.4]
  assign _T_157 = _T_154 & _T_156; // @[Controllers.scala 165:74:@28865.4]
  assign _T_161 = _T_157 & io_enable; // @[Controllers.scala 165:109:@28868.4]
  assign _T_164 = io_ctrCopyDone_0 == 1'h0; // @[Controllers.scala 165:141:@28870.4]
  assign _T_172 = RetimeWrapper_io_out; // @[package.scala 96:25:@28882.4 package.scala 96:25:@28883.4]
  assign _T_176 = _T_172 == 1'h0; // @[Controllers.scala 167:54:@28885.4]
  assign _T_177 = io_doneIn_0 | _T_176; // @[Controllers.scala 167:52:@28886.4]
  assign _T_184 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@28896.4 package.scala 96:25:@28897.4]
  assign _T_202 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@28914.4 package.scala 96:25:@28915.4]
  assign _T_206 = _T_202 == 1'h0; // @[Controllers.scala 169:67:@28917.4]
  assign _T_207 = _T_206 & io_enable; // @[Controllers.scala 169:86:@28918.4]
  assign _T_219 = ~ iterDone_1_io_output; // @[Controllers.scala 165:35:@28930.4]
  assign _T_221 = io_doneIn_1 == 1'h0; // @[Controllers.scala 165:60:@28931.4]
  assign _T_222 = _T_219 & _T_221; // @[Controllers.scala 165:58:@28932.4]
  assign _T_224 = done_1_io_output == 1'h0; // @[Controllers.scala 165:76:@28933.4]
  assign _T_225 = _T_222 & _T_224; // @[Controllers.scala 165:74:@28934.4]
  assign _T_229 = _T_225 & io_enable; // @[Controllers.scala 165:109:@28937.4]
  assign _T_232 = io_ctrCopyDone_1 == 1'h0; // @[Controllers.scala 165:141:@28939.4]
  assign _T_240 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@28951.4 package.scala 96:25:@28952.4]
  assign _T_244 = _T_240 == 1'h0; // @[Controllers.scala 167:54:@28954.4]
  assign _T_245 = io_doneIn_1 | _T_244; // @[Controllers.scala 167:52:@28955.4]
  assign _T_252 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@28965.4 package.scala 96:25:@28966.4]
  assign _T_270 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@28983.4 package.scala 96:25:@28984.4]
  assign _T_274 = _T_270 == 1'h0; // @[Controllers.scala 169:67:@28986.4]
  assign _T_275 = _T_274 & io_enable; // @[Controllers.scala 169:86:@28987.4]
  assign _T_287 = ~ iterDone_2_io_output; // @[Controllers.scala 165:35:@28999.4]
  assign _T_289 = io_doneIn_2 == 1'h0; // @[Controllers.scala 165:60:@29000.4]
  assign _T_290 = _T_287 & _T_289; // @[Controllers.scala 165:58:@29001.4]
  assign _T_292 = done_2_io_output == 1'h0; // @[Controllers.scala 165:76:@29002.4]
  assign _T_293 = _T_290 & _T_292; // @[Controllers.scala 165:74:@29003.4]
  assign _T_297 = _T_293 & io_enable; // @[Controllers.scala 165:109:@29006.4]
  assign _T_300 = io_ctrCopyDone_2 == 1'h0; // @[Controllers.scala 165:141:@29008.4]
  assign _T_308 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@29020.4 package.scala 96:25:@29021.4]
  assign _T_312 = _T_308 == 1'h0; // @[Controllers.scala 167:54:@29023.4]
  assign _T_313 = io_doneIn_2 | _T_312; // @[Controllers.scala 167:52:@29024.4]
  assign _T_320 = RetimeWrapper_7_io_out; // @[package.scala 96:25:@29034.4 package.scala 96:25:@29035.4]
  assign _T_338 = RetimeWrapper_8_io_out; // @[package.scala 96:25:@29052.4 package.scala 96:25:@29053.4]
  assign _T_342 = _T_338 == 1'h0; // @[Controllers.scala 169:67:@29055.4]
  assign _T_343 = _T_342 & io_enable; // @[Controllers.scala 169:86:@29056.4]
  assign _T_358 = io_enable & active_0_io_output; // @[Controllers.scala 213:68:@29074.4]
  assign _T_360 = _T_358 & _T_151; // @[Controllers.scala 213:90:@29076.4]
  assign _T_362 = ~ allDone; // @[Controllers.scala 213:132:@29078.4]
  assign _T_366 = io_enable & active_1_io_output; // @[Controllers.scala 213:68:@29083.4]
  assign _T_368 = _T_366 & _T_219; // @[Controllers.scala 213:90:@29085.4]
  assign _T_374 = io_enable & active_2_io_output; // @[Controllers.scala 213:68:@29091.4]
  assign _T_376 = _T_374 & _T_287; // @[Controllers.scala 213:90:@29093.4]
  assign _T_383 = allDone == 1'h0; // @[package.scala 100:49:@29099.4]
  assign _T_387 = allDone & _T_386; // @[package.scala 100:41:@29102.4]
  assign io_done = RetimeWrapper_10_io_out; // @[Controllers.scala 245:13:@29128.4]
  assign io_enableOut_0 = _T_360 & _T_362; // @[Controllers.scala 213:55:@29082.4]
  assign io_enableOut_1 = _T_368 & _T_362; // @[Controllers.scala 213:55:@29090.4]
  assign io_enableOut_2 = _T_376 & _T_362; // @[Controllers.scala 213:55:@29098.4]
  assign io_childAck_0 = iterDone_0_io_output; // @[Controllers.scala 212:58:@29069.4]
  assign io_childAck_1 = iterDone_1_io_output; // @[Controllers.scala 212:58:@29071.4]
  assign io_childAck_2 = iterDone_2_io_output; // @[Controllers.scala 212:58:@29073.4]
  assign active_0_clock = clock; // @[:@28765.4]
  assign active_0_reset = reset; // @[:@28766.4]
  assign active_0_io_input_set = _T_161 & _T_164; // @[Controllers.scala 165:32:@28872.4]
  assign active_0_io_input_reset = io_ctrCopyDone_0 | io_parentAck; // @[Controllers.scala 166:34:@28876.4]
  assign active_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@28786.4]
  assign active_1_clock = clock; // @[:@28768.4]
  assign active_1_reset = reset; // @[:@28769.4]
  assign active_1_io_input_set = _T_229 & _T_232; // @[Controllers.scala 165:32:@28941.4]
  assign active_1_io_input_reset = io_ctrCopyDone_1 | io_parentAck; // @[Controllers.scala 166:34:@28945.4]
  assign active_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@28787.4]
  assign active_2_clock = clock; // @[:@28771.4]
  assign active_2_reset = reset; // @[:@28772.4]
  assign active_2_io_input_set = _T_297 & _T_300; // @[Controllers.scala 165:32:@29010.4]
  assign active_2_io_input_reset = io_ctrCopyDone_2 | io_parentAck; // @[Controllers.scala 166:34:@29014.4]
  assign active_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 84:40:@28788.4]
  assign done_0_clock = clock; // @[:@28774.4]
  assign done_0_reset = reset; // @[:@28775.4]
  assign done_0_io_input_set = io_ctrCopyDone_0 | _T_207; // @[Controllers.scala 169:30:@28922.4]
  assign done_0_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@28800.4 Controllers.scala 170:32:@28929.4]
  assign done_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@28789.4]
  assign done_1_clock = clock; // @[:@28777.4]
  assign done_1_reset = reset; // @[:@28778.4]
  assign done_1_io_input_set = io_ctrCopyDone_1 | _T_275; // @[Controllers.scala 169:30:@28991.4]
  assign done_1_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@28809.4 Controllers.scala 170:32:@28998.4]
  assign done_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@28790.4]
  assign done_2_clock = clock; // @[:@28780.4]
  assign done_2_reset = reset; // @[:@28781.4]
  assign done_2_io_input_set = io_ctrCopyDone_2 | _T_343; // @[Controllers.scala 169:30:@29060.4]
  assign done_2_io_input_reset = io_parentAck; // @[Controllers.scala 86:33:@28818.4 Controllers.scala 170:32:@29067.4]
  assign done_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 85:38:@28791.4]
  assign iterDone_0_clock = clock; // @[:@28821.4]
  assign iterDone_0_reset = reset; // @[:@28822.4]
  assign iterDone_0_io_input_set = _T_177 & io_enable; // @[Controllers.scala 167:34:@28890.4]
  assign iterDone_0_io_input_reset = _T_184 | io_parentAck; // @[Controllers.scala 92:37:@28840.4 Controllers.scala 168:36:@28906.4]
  assign iterDone_0_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@28829.4]
  assign iterDone_1_clock = clock; // @[:@28824.4]
  assign iterDone_1_reset = reset; // @[:@28825.4]
  assign iterDone_1_io_input_set = _T_245 & io_enable; // @[Controllers.scala 167:34:@28959.4]
  assign iterDone_1_io_input_reset = _T_252 | io_parentAck; // @[Controllers.scala 92:37:@28849.4 Controllers.scala 168:36:@28975.4]
  assign iterDone_1_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@28830.4]
  assign iterDone_2_clock = clock; // @[:@28827.4]
  assign iterDone_2_reset = reset; // @[:@28828.4]
  assign iterDone_2_io_input_set = _T_313 & io_enable; // @[Controllers.scala 167:34:@29028.4]
  assign iterDone_2_io_input_reset = _T_320 | io_parentAck; // @[Controllers.scala 92:37:@28858.4 Controllers.scala 168:36:@29044.4]
  assign iterDone_2_io_input_asyn_reset = 1'h0; // @[Controllers.scala 91:42:@28831.4]
  assign RetimeWrapper_clock = clock; // @[:@28878.4]
  assign RetimeWrapper_reset = reset; // @[:@28879.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@28881.4]
  assign RetimeWrapper_io_in = 1'h1; // @[package.scala 94:16:@28880.4]
  assign RetimeWrapper_1_clock = clock; // @[:@28892.4]
  assign RetimeWrapper_1_reset = reset; // @[:@28893.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@28895.4]
  assign RetimeWrapper_1_io_in = io_doneIn_0; // @[package.scala 94:16:@28894.4]
  assign RetimeWrapper_2_clock = clock; // @[:@28910.4]
  assign RetimeWrapper_2_reset = reset; // @[:@28911.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@28913.4]
  assign RetimeWrapper_2_io_in = 1'h1; // @[package.scala 94:16:@28912.4]
  assign RetimeWrapper_3_clock = clock; // @[:@28947.4]
  assign RetimeWrapper_3_reset = reset; // @[:@28948.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@28950.4]
  assign RetimeWrapper_3_io_in = 1'h1; // @[package.scala 94:16:@28949.4]
  assign RetimeWrapper_4_clock = clock; // @[:@28961.4]
  assign RetimeWrapper_4_reset = reset; // @[:@28962.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@28964.4]
  assign RetimeWrapper_4_io_in = io_doneIn_1; // @[package.scala 94:16:@28963.4]
  assign RetimeWrapper_5_clock = clock; // @[:@28979.4]
  assign RetimeWrapper_5_reset = reset; // @[:@28980.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@28982.4]
  assign RetimeWrapper_5_io_in = 1'h1; // @[package.scala 94:16:@28981.4]
  assign RetimeWrapper_6_clock = clock; // @[:@29016.4]
  assign RetimeWrapper_6_reset = reset; // @[:@29017.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@29019.4]
  assign RetimeWrapper_6_io_in = 1'h1; // @[package.scala 94:16:@29018.4]
  assign RetimeWrapper_7_clock = clock; // @[:@29030.4]
  assign RetimeWrapper_7_reset = reset; // @[:@29031.4]
  assign RetimeWrapper_7_io_flow = 1'h1; // @[package.scala 95:18:@29033.4]
  assign RetimeWrapper_7_io_in = io_doneIn_2; // @[package.scala 94:16:@29032.4]
  assign RetimeWrapper_8_clock = clock; // @[:@29048.4]
  assign RetimeWrapper_8_reset = reset; // @[:@29049.4]
  assign RetimeWrapper_8_io_flow = 1'h1; // @[package.scala 95:18:@29051.4]
  assign RetimeWrapper_8_io_in = 1'h1; // @[package.scala 94:16:@29050.4]
  assign RetimeWrapper_9_clock = clock; // @[:@29105.4]
  assign RetimeWrapper_9_reset = reset; // @[:@29106.4]
  assign RetimeWrapper_9_io_flow = 1'h1; // @[package.scala 95:18:@29108.4]
  assign RetimeWrapper_9_io_in = _T_387 | io_parentAck; // @[package.scala 94:16:@29107.4]
  assign RetimeWrapper_10_clock = clock; // @[:@29122.4]
  assign RetimeWrapper_10_reset = reset; // @[:@29123.4]
  assign RetimeWrapper_10_io_flow = io_enable; // @[package.scala 95:18:@29125.4]
  assign RetimeWrapper_10_io_in = allDone & _T_400; // @[package.scala 94:16:@29124.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_386 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_400 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_386 <= 1'h0;
    end else begin
      _T_386 <= _T_383;
    end
    if (reset) begin
      _T_400 <= 1'h0;
    end else begin
      _T_400 <= _T_383;
    end
  end
endmodule
module x411_inr_UnitPipe_sm( // @[:@29301.2]
  input   clock, // @[:@29302.4]
  input   reset, // @[:@29303.4]
  input   io_enable, // @[:@29304.4]
  output  io_done, // @[:@29304.4]
  output  io_doneLatch, // @[:@29304.4]
  input   io_ctrDone, // @[:@29304.4]
  output  io_datapathEn, // @[:@29304.4]
  output  io_ctrInc, // @[:@29304.4]
  input   io_parentAck, // @[:@29304.4]
  input   io_backpressure // @[:@29304.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@29306.4]
  wire  active_reset; // @[Controllers.scala 261:22:@29306.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@29306.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@29306.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@29306.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@29306.4]
  wire  done_clock; // @[Controllers.scala 262:20:@29309.4]
  wire  done_reset; // @[Controllers.scala 262:20:@29309.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@29309.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@29309.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@29309.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@29309.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29363.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29371.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29371.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29371.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29371.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29371.4]
  wire  _T_80; // @[Controllers.scala 264:48:@29314.4]
  wire  _T_81; // @[Controllers.scala 264:46:@29315.4]
  wire  _T_82; // @[Controllers.scala 264:62:@29316.4]
  wire  _T_83; // @[Controllers.scala 264:60:@29317.4]
  wire  _T_100; // @[package.scala 100:49:@29334.4]
  reg  _T_103; // @[package.scala 48:56:@29335.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 100:49:@29343.4]
  wire  _T_116; // @[Controllers.scala 283:41:@29351.4]
  wire  _T_117; // @[Controllers.scala 283:59:@29352.4]
  wire  _T_119; // @[Controllers.scala 284:37:@29355.4]
  reg  _T_125; // @[package.scala 48:56:@29359.4]
  reg [31:0] _RAND_1;
  reg  _T_142; // @[Controllers.scala 291:31:@29381.4]
  reg [31:0] _RAND_2;
  reg  _T_149; // @[package.scala 48:56:@29384.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:41:@29386.4]
  wire  _T_152; // @[Controllers.scala 292:61:@29387.4]
  wire  _T_153; // @[Controllers.scala 292:24:@29388.4]
  SRFF active ( // @[Controllers.scala 261:22:@29306.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@29309.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@29363.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@29371.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@29314.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@29315.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@29316.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@29317.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@29334.4]
  assign _T_108 = done_io_output == 1'h0; // @[package.scala 100:49:@29343.4]
  assign _T_116 = active_io_output & _T_82; // @[Controllers.scala 283:41:@29351.4]
  assign _T_117 = _T_116 & io_enable; // @[Controllers.scala 283:59:@29352.4]
  assign _T_119 = active_io_output & io_enable; // @[Controllers.scala 284:37:@29355.4]
  assign _T_150 = done_io_output & _T_149; // @[package.scala 100:41:@29386.4]
  assign _T_152 = _T_150 ? 1'h1 : _T_142; // @[Controllers.scala 292:61:@29387.4]
  assign _T_153 = io_parentAck ? 1'h0 : _T_152; // @[Controllers.scala 292:24:@29388.4]
  assign io_done = done_io_output & _T_125; // @[Controllers.scala 287:13:@29362.4]
  assign io_doneLatch = _T_142; // @[Controllers.scala 293:18:@29390.4]
  assign io_datapathEn = _T_117 & io_backpressure; // @[Controllers.scala 283:21:@29354.4]
  assign io_ctrInc = _T_119 & io_backpressure; // @[Controllers.scala 284:17:@29357.4]
  assign active_clock = clock; // @[:@29307.4]
  assign active_reset = reset; // @[:@29308.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@29319.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@29323.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@29324.4]
  assign done_clock = clock; // @[:@29310.4]
  assign done_reset = reset; // @[:@29311.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@29339.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@29332.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@29333.4]
  assign RetimeWrapper_clock = clock; // @[:@29364.4]
  assign RetimeWrapper_reset = reset; // @[:@29365.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@29367.4]
  assign RetimeWrapper_io_in = 1'h0; // @[package.scala 94:16:@29366.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29372.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29373.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@29375.4]
  assign RetimeWrapper_1_io_in = io_ctrDone; // @[package.scala 94:16:@29374.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_125 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_142 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_149 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_125 <= 1'h0;
    end else begin
      _T_125 <= _T_108;
    end
    if (reset) begin
      _T_142 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_142 <= 1'h0;
      end else begin
        if (_T_150) begin
          _T_142 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_149 <= 1'h0;
    end else begin
      _T_149 <= _T_108;
    end
  end
endmodule
module x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1( // @[:@29465.2]
  output        io_in_x404_valid, // @[:@29468.4]
  output [63:0] io_in_x404_bits_addr, // @[:@29468.4]
  output [31:0] io_in_x404_bits_size, // @[:@29468.4]
  input  [63:0] io_in_x219_outdram_number, // @[:@29468.4]
  input         io_sigsIn_backpressure, // @[:@29468.4]
  input         io_sigsIn_datapathEn, // @[:@29468.4]
  input         io_rr // @[:@29468.4]
);
  wire [96:0] x408_tuple; // @[Cat.scala 30:58:@29482.4]
  wire  _T_135; // @[implicits.scala 55:10:@29485.4]
  assign x408_tuple = {33'h7e9000,io_in_x219_outdram_number}; // @[Cat.scala 30:58:@29482.4]
  assign _T_135 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@29485.4]
  assign io_in_x404_valid = _T_135 & io_sigsIn_backpressure; // @[sm_x411_inr_UnitPipe.scala 65:18:@29488.4]
  assign io_in_x404_bits_addr = x408_tuple[63:0]; // @[sm_x411_inr_UnitPipe.scala 66:22:@29490.4]
  assign io_in_x404_bits_size = x408_tuple[95:64]; // @[sm_x411_inr_UnitPipe.scala 67:22:@29492.4]
endmodule
module FF_13( // @[:@29494.2]
  input         clock, // @[:@29495.4]
  input         reset, // @[:@29496.4]
  output [22:0] io_rPort_0_output_0, // @[:@29497.4]
  input  [22:0] io_wPort_0_data_0, // @[:@29497.4]
  input         io_wPort_0_reset, // @[:@29497.4]
  input         io_wPort_0_en_0 // @[:@29497.4]
);
  reg [22:0] ff; // @[MemPrimitives.scala 321:19:@29512.4]
  reg [31:0] _RAND_0;
  wire [22:0] _T_68; // @[MemPrimitives.scala 325:32:@29514.4]
  wire [22:0] _T_69; // @[MemPrimitives.scala 325:12:@29515.4]
  assign _T_68 = io_wPort_0_en_0 ? io_wPort_0_data_0 : ff; // @[MemPrimitives.scala 325:32:@29514.4]
  assign _T_69 = io_wPort_0_reset ? 23'h0 : _T_68; // @[MemPrimitives.scala 325:12:@29515.4]
  assign io_rPort_0_output_0 = ff; // @[MemPrimitives.scala 326:34:@29517.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff = _RAND_0[22:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      ff <= 23'h0;
    end else begin
      if (io_wPort_0_reset) begin
        ff <= 23'h0;
      end else begin
        if (io_wPort_0_en_0) begin
          ff <= io_wPort_0_data_0;
        end
      end
    end
  end
endmodule
module SingleCounter_5( // @[:@29532.2]
  input         clock, // @[:@29533.4]
  input         reset, // @[:@29534.4]
  input         io_input_reset, // @[:@29535.4]
  input         io_input_enable, // @[:@29535.4]
  output [22:0] io_output_count_0, // @[:@29535.4]
  output        io_output_oobs_0, // @[:@29535.4]
  output        io_output_done // @[:@29535.4]
);
  wire  bases_0_clock; // @[Counter.scala 261:53:@29548.4]
  wire  bases_0_reset; // @[Counter.scala 261:53:@29548.4]
  wire [22:0] bases_0_io_rPort_0_output_0; // @[Counter.scala 261:53:@29548.4]
  wire [22:0] bases_0_io_wPort_0_data_0; // @[Counter.scala 261:53:@29548.4]
  wire  bases_0_io_wPort_0_reset; // @[Counter.scala 261:53:@29548.4]
  wire  bases_0_io_wPort_0_en_0; // @[Counter.scala 261:53:@29548.4]
  wire  SRFF_clock; // @[Counter.scala 263:22:@29564.4]
  wire  SRFF_reset; // @[Counter.scala 263:22:@29564.4]
  wire  SRFF_io_input_set; // @[Counter.scala 263:22:@29564.4]
  wire  SRFF_io_input_reset; // @[Counter.scala 263:22:@29564.4]
  wire  SRFF_io_input_asyn_reset; // @[Counter.scala 263:22:@29564.4]
  wire  SRFF_io_output; // @[Counter.scala 263:22:@29564.4]
  wire  _T_36; // @[Counter.scala 264:45:@29567.4]
  wire [22:0] _T_48; // @[Counter.scala 287:52:@29592.4]
  wire [23:0] _T_50; // @[Counter.scala 291:33:@29593.4]
  wire [22:0] _T_51; // @[Counter.scala 291:33:@29594.4]
  wire [22:0] _T_52; // @[Counter.scala 291:33:@29595.4]
  wire  _T_57; // @[Counter.scala 293:18:@29597.4]
  wire [22:0] _T_68; // @[Counter.scala 299:115:@29605.4]
  wire [22:0] _T_71; // @[Counter.scala 299:152:@29608.4]
  wire [22:0] _T_72; // @[Counter.scala 299:74:@29609.4]
  wire  _T_75; // @[Counter.scala 322:102:@29613.4]
  wire  _T_77; // @[Counter.scala 322:130:@29614.4]
  FF_13 bases_0 ( // @[Counter.scala 261:53:@29548.4]
    .clock(bases_0_clock),
    .reset(bases_0_reset),
    .io_rPort_0_output_0(bases_0_io_rPort_0_output_0),
    .io_wPort_0_data_0(bases_0_io_wPort_0_data_0),
    .io_wPort_0_reset(bases_0_io_wPort_0_reset),
    .io_wPort_0_en_0(bases_0_io_wPort_0_en_0)
  );
  SRFF SRFF ( // @[Counter.scala 263:22:@29564.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  assign _T_36 = io_input_reset == 1'h0; // @[Counter.scala 264:45:@29567.4]
  assign _T_48 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 287:52:@29592.4]
  assign _T_50 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@29593.4]
  assign _T_51 = $signed(_T_48) + $signed(23'sh1); // @[Counter.scala 291:33:@29594.4]
  assign _T_52 = $signed(_T_51); // @[Counter.scala 291:33:@29595.4]
  assign _T_57 = $signed(_T_52) >= $signed(23'sh1fa400); // @[Counter.scala 293:18:@29597.4]
  assign _T_68 = $unsigned(_T_48); // @[Counter.scala 299:115:@29605.4]
  assign _T_71 = $unsigned(_T_52); // @[Counter.scala 299:152:@29608.4]
  assign _T_72 = _T_57 ? _T_68 : _T_71; // @[Counter.scala 299:74:@29609.4]
  assign _T_75 = $signed(_T_48) < $signed(23'sh0); // @[Counter.scala 322:102:@29613.4]
  assign _T_77 = $signed(_T_48) >= $signed(23'sh1fa400); // @[Counter.scala 322:130:@29614.4]
  assign io_output_count_0 = $signed(bases_0_io_rPort_0_output_0); // @[Counter.scala 304:28:@29612.4]
  assign io_output_oobs_0 = _T_75 | _T_77; // @[Counter.scala 322:60:@29616.4]
  assign io_output_done = io_input_enable & _T_57; // @[Counter.scala 333:20:@29618.4]
  assign bases_0_clock = clock; // @[:@29549.4]
  assign bases_0_reset = reset; // @[:@29550.4]
  assign bases_0_io_wPort_0_data_0 = io_input_reset ? 23'h0 : _T_72; // @[Counter.scala 299:31:@29611.4]
  assign bases_0_io_wPort_0_reset = io_input_reset; // @[Counter.scala 281:27:@29590.4]
  assign bases_0_io_wPort_0_en_0 = io_input_enable; // @[Counter.scala 284:29:@29591.4]
  assign SRFF_clock = clock; // @[:@29565.4]
  assign SRFF_reset = reset; // @[:@29566.4]
  assign SRFF_io_input_set = io_input_enable & _T_36; // @[Counter.scala 264:23:@29569.4]
  assign SRFF_io_input_reset = io_input_reset | io_output_done; // @[Counter.scala 265:25:@29571.4]
  assign SRFF_io_input_asyn_reset = 1'h0; // @[Counter.scala 266:30:@29572.4]
endmodule
module x413_ctrchain( // @[:@29623.2]
  input         clock, // @[:@29624.4]
  input         reset, // @[:@29625.4]
  input         io_input_reset, // @[:@29626.4]
  input         io_input_enable, // @[:@29626.4]
  output [22:0] io_output_counts_0, // @[:@29626.4]
  output        io_output_oobs_0, // @[:@29626.4]
  output        io_output_done // @[:@29626.4]
);
  wire  ctrs_0_clock; // @[Counter.scala 513:46:@29628.4]
  wire  ctrs_0_reset; // @[Counter.scala 513:46:@29628.4]
  wire  ctrs_0_io_input_reset; // @[Counter.scala 513:46:@29628.4]
  wire  ctrs_0_io_input_enable; // @[Counter.scala 513:46:@29628.4]
  wire [22:0] ctrs_0_io_output_count_0; // @[Counter.scala 513:46:@29628.4]
  wire  ctrs_0_io_output_oobs_0; // @[Counter.scala 513:46:@29628.4]
  wire  ctrs_0_io_output_done; // @[Counter.scala 513:46:@29628.4]
  reg  wasDone; // @[Counter.scala 542:24:@29637.4]
  reg [31:0] _RAND_0;
  wire  _T_45; // @[Counter.scala 546:69:@29643.4]
  wire  _T_47; // @[Counter.scala 546:80:@29644.4]
  reg  doneLatch; // @[Counter.scala 550:26:@29649.4]
  reg [31:0] _RAND_1;
  wire  _T_54; // @[Counter.scala 551:48:@29650.4]
  wire  _T_55; // @[Counter.scala 551:19:@29651.4]
  SingleCounter_5 ctrs_0 ( // @[Counter.scala 513:46:@29628.4]
    .clock(ctrs_0_clock),
    .reset(ctrs_0_reset),
    .io_input_reset(ctrs_0_io_input_reset),
    .io_input_enable(ctrs_0_io_input_enable),
    .io_output_count_0(ctrs_0_io_output_count_0),
    .io_output_oobs_0(ctrs_0_io_output_oobs_0),
    .io_output_done(ctrs_0_io_output_done)
  );
  assign _T_45 = io_input_enable & ctrs_0_io_output_done; // @[Counter.scala 546:69:@29643.4]
  assign _T_47 = wasDone == 1'h0; // @[Counter.scala 546:80:@29644.4]
  assign _T_54 = ctrs_0_io_output_done ? 1'h1 : doneLatch; // @[Counter.scala 551:48:@29650.4]
  assign _T_55 = io_input_reset ? 1'h0 : _T_54; // @[Counter.scala 551:19:@29651.4]
  assign io_output_counts_0 = ctrs_0_io_output_count_0; // @[Counter.scala 557:32:@29653.4]
  assign io_output_oobs_0 = ctrs_0_io_output_oobs_0 | doneLatch; // @[Counter.scala 558:30:@29655.4]
  assign io_output_done = _T_45 & _T_47; // @[Counter.scala 546:18:@29646.4]
  assign ctrs_0_clock = clock; // @[:@29629.4]
  assign ctrs_0_reset = reset; // @[:@29630.4]
  assign ctrs_0_io_input_reset = io_input_reset; // @[Counter.scala 520:24:@29634.4]
  assign ctrs_0_io_input_enable = io_input_enable; // @[Counter.scala 524:33:@29635.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  wasDone = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  doneLatch = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      wasDone <= 1'h0;
    end else begin
      wasDone <= ctrs_0_io_output_done;
    end
    if (reset) begin
      doneLatch <= 1'h0;
    end else begin
      if (io_input_reset) begin
        doneLatch <= 1'h0;
      end else begin
        if (ctrs_0_io_output_done) begin
          doneLatch <= 1'h1;
        end
      end
    end
  end
endmodule
module x420_inr_Foreach_sm( // @[:@29843.2]
  input   clock, // @[:@29844.4]
  input   reset, // @[:@29845.4]
  input   io_enable, // @[:@29846.4]
  output  io_done, // @[:@29846.4]
  output  io_doneLatch, // @[:@29846.4]
  input   io_ctrDone, // @[:@29846.4]
  output  io_datapathEn, // @[:@29846.4]
  output  io_ctrInc, // @[:@29846.4]
  output  io_ctrRst, // @[:@29846.4]
  input   io_parentAck, // @[:@29846.4]
  input   io_backpressure, // @[:@29846.4]
  input   io_break // @[:@29846.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@29848.4]
  wire  active_reset; // @[Controllers.scala 261:22:@29848.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@29848.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@29848.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@29848.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@29848.4]
  wire  done_clock; // @[Controllers.scala 262:20:@29851.4]
  wire  done_reset; // @[Controllers.scala 262:20:@29851.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@29851.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@29851.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@29851.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@29851.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@29885.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@29885.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@29885.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@29885.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@29885.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@29907.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@29907.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@29907.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@29907.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@29907.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@29919.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@29927.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@29927.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@29927.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@29927.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@29927.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@29943.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@29943.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@29943.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@29943.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@29943.4]
  wire  _T_80; // @[Controllers.scala 264:48:@29856.4]
  wire  _T_81; // @[Controllers.scala 264:46:@29857.4]
  wire  _T_82; // @[Controllers.scala 264:62:@29858.4]
  wire  _T_83; // @[Controllers.scala 264:60:@29859.4]
  wire  _T_100; // @[package.scala 100:49:@29876.4]
  reg  _T_103; // @[package.scala 48:56:@29877.4]
  reg [31:0] _RAND_0;
  wire  _T_108; // @[package.scala 96:25:@29890.4 package.scala 96:25:@29891.4]
  wire  _T_110; // @[package.scala 100:49:@29892.4]
  reg  _T_113; // @[package.scala 48:56:@29893.4]
  reg [31:0] _RAND_1;
  wire  _T_114; // @[package.scala 100:41:@29895.4]
  wire  _T_118; // @[Controllers.scala 283:41:@29900.4]
  wire  _T_119; // @[Controllers.scala 283:59:@29901.4]
  wire  _T_121; // @[Controllers.scala 284:37:@29904.4]
  wire  _T_124; // @[package.scala 96:25:@29912.4 package.scala 96:25:@29913.4]
  wire  _T_126; // @[package.scala 100:49:@29914.4]
  reg  _T_129; // @[package.scala 48:56:@29915.4]
  reg [31:0] _RAND_2;
  reg  _T_146; // @[Controllers.scala 291:31:@29937.4]
  reg [31:0] _RAND_3;
  wire  _T_150; // @[package.scala 100:49:@29939.4]
  reg  _T_153; // @[package.scala 48:56:@29940.4]
  reg [31:0] _RAND_4;
  wire  _T_156; // @[package.scala 96:25:@29948.4 package.scala 96:25:@29949.4]
  wire  _T_158; // @[Controllers.scala 292:61:@29950.4]
  wire  _T_159; // @[Controllers.scala 292:24:@29951.4]
  SRFF active ( // @[Controllers.scala 261:22:@29848.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@29851.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@29885.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@29907.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@29919.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@29927.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@29943.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@29856.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@29857.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@29858.4]
  assign _T_83 = _T_81 & _T_82; // @[Controllers.scala 264:60:@29859.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@29876.4]
  assign _T_108 = RetimeWrapper_io_out; // @[package.scala 96:25:@29890.4 package.scala 96:25:@29891.4]
  assign _T_110 = _T_108 == 1'h0; // @[package.scala 100:49:@29892.4]
  assign _T_114 = _T_108 & _T_113; // @[package.scala 100:41:@29895.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@29900.4]
  assign _T_119 = _T_118 & io_enable; // @[Controllers.scala 283:59:@29901.4]
  assign _T_121 = active_io_output & io_enable; // @[Controllers.scala 284:37:@29904.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@29912.4 package.scala 96:25:@29913.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@29914.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@29939.4]
  assign _T_156 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@29948.4 package.scala 96:25:@29949.4]
  assign _T_158 = _T_156 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@29950.4]
  assign _T_159 = io_parentAck ? 1'h0 : _T_158; // @[Controllers.scala 292:24:@29951.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@29918.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@29953.4]
  assign io_datapathEn = _T_119 & io_backpressure; // @[Controllers.scala 283:21:@29903.4]
  assign io_ctrInc = _T_121 & io_backpressure; // @[Controllers.scala 284:17:@29906.4]
  assign io_ctrRst = _T_114 | io_parentAck; // @[Controllers.scala 274:13:@29898.4]
  assign active_clock = clock; // @[:@29849.4]
  assign active_reset = reset; // @[:@29850.4]
  assign active_io_input_set = _T_83 & io_backpressure; // @[Controllers.scala 264:23:@29861.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@29865.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@29866.4]
  assign done_clock = clock; // @[:@29852.4]
  assign done_reset = reset; // @[:@29853.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@29881.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@29874.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@29875.4]
  assign RetimeWrapper_clock = clock; // @[:@29886.4]
  assign RetimeWrapper_reset = reset; // @[:@29887.4]
  assign RetimeWrapper_io_flow = io_backpressure; // @[package.scala 95:18:@29889.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@29888.4]
  assign RetimeWrapper_1_clock = clock; // @[:@29908.4]
  assign RetimeWrapper_1_reset = reset; // @[:@29909.4]
  assign RetimeWrapper_1_io_flow = io_backpressure; // @[package.scala 95:18:@29911.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@29910.4]
  assign RetimeWrapper_2_clock = clock; // @[:@29920.4]
  assign RetimeWrapper_2_reset = reset; // @[:@29921.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@29923.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@29922.4]
  assign RetimeWrapper_3_clock = clock; // @[:@29928.4]
  assign RetimeWrapper_3_reset = reset; // @[:@29929.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@29931.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@29930.4]
  assign RetimeWrapper_4_clock = clock; // @[:@29944.4]
  assign RetimeWrapper_4_reset = reset; // @[:@29945.4]
  assign RetimeWrapper_4_io_flow = io_backpressure; // @[package.scala 95:18:@29947.4]
  assign RetimeWrapper_4_io_in = done_io_output & _T_153; // @[package.scala 94:16:@29946.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_113 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_129 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_146 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_153 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_113 <= 1'h0;
    end else begin
      _T_113 <= _T_110;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_156) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x420_inr_Foreach_kernelx420_inr_Foreach_concrete1( // @[:@30160.2]
  input         clock, // @[:@30161.4]
  input         reset, // @[:@30162.4]
  output [20:0] io_in_x223_outbuf_0_rPort_0_ofs_0, // @[:@30163.4]
  output        io_in_x223_outbuf_0_rPort_0_en_0, // @[:@30163.4]
  output        io_in_x223_outbuf_0_rPort_0_backpressure, // @[:@30163.4]
  input  [31:0] io_in_x223_outbuf_0_rPort_0_output_0, // @[:@30163.4]
  output        io_in_x405_valid, // @[:@30163.4]
  output [31:0] io_in_x405_bits_wdata_0, // @[:@30163.4]
  output        io_in_x405_bits_wstrb, // @[:@30163.4]
  input         io_sigsIn_backpressure, // @[:@30163.4]
  input         io_sigsIn_datapathEn, // @[:@30163.4]
  input         io_sigsIn_break, // @[:@30163.4]
  input  [31:0] io_sigsIn_cchainOutputs_0_counts_0, // @[:@30163.4]
  input         io_sigsIn_cchainOutputs_0_oobs_0, // @[:@30163.4]
  input         io_rr // @[:@30163.4]
);
  wire [31:0] __io_b; // @[Math.scala 720:24:@30190.4]
  wire [31:0] __io_result; // @[Math.scala 720:24:@30190.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30219.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30219.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30219.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30219.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30219.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30228.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30228.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30228.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30228.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30228.4]
  wire  b415; // @[sm_x420_inr_Foreach.scala 62:18:@30198.4]
  wire  _T_274; // @[sm_x420_inr_Foreach.scala 67:129:@30202.4]
  wire  _T_278; // @[implicits.scala 55:10:@30205.4]
  wire  _T_279; // @[sm_x420_inr_Foreach.scala 67:146:@30206.4]
  wire [32:0] x418_tuple; // @[Cat.scala 30:58:@30216.4]
  wire  _T_290; // @[package.scala 96:25:@30233.4 package.scala 96:25:@30234.4]
  wire  _T_292; // @[implicits.scala 55:10:@30235.4]
  wire  x533_b415_D2; // @[package.scala 96:25:@30224.4 package.scala 96:25:@30225.4]
  wire  _T_293; // @[sm_x420_inr_Foreach.scala 74:112:@30236.4]
  wire [31:0] b414_number; // @[Math.scala 723:22:@30195.4 Math.scala 724:14:@30196.4]
  _ _ ( // @[Math.scala 720:24:@30190.4]
    .io_b(__io_b),
    .io_result(__io_result)
  );
  RetimeWrapper_6 RetimeWrapper ( // @[package.scala 93:22:@30219.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper_6 RetimeWrapper_1 ( // @[package.scala 93:22:@30228.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  assign b415 = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x420_inr_Foreach.scala 62:18:@30198.4]
  assign _T_274 = ~ io_sigsIn_break; // @[sm_x420_inr_Foreach.scala 67:129:@30202.4]
  assign _T_278 = io_rr ? io_sigsIn_datapathEn : 1'h0; // @[implicits.scala 55:10:@30205.4]
  assign _T_279 = _T_274 & _T_278; // @[sm_x420_inr_Foreach.scala 67:146:@30206.4]
  assign x418_tuple = {1'h1,io_in_x223_outbuf_0_rPort_0_output_0}; // @[Cat.scala 30:58:@30216.4]
  assign _T_290 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30233.4 package.scala 96:25:@30234.4]
  assign _T_292 = io_rr ? _T_290 : 1'h0; // @[implicits.scala 55:10:@30235.4]
  assign x533_b415_D2 = RetimeWrapper_io_out; // @[package.scala 96:25:@30224.4 package.scala 96:25:@30225.4]
  assign _T_293 = _T_292 & x533_b415_D2; // @[sm_x420_inr_Foreach.scala 74:112:@30236.4]
  assign b414_number = __io_result; // @[Math.scala 723:22:@30195.4 Math.scala 724:14:@30196.4]
  assign io_in_x223_outbuf_0_rPort_0_ofs_0 = b414_number[20:0]; // @[MemInterfaceType.scala 107:54:@30209.4]
  assign io_in_x223_outbuf_0_rPort_0_en_0 = _T_279 & b415; // @[MemInterfaceType.scala 110:79:@30211.4]
  assign io_in_x223_outbuf_0_rPort_0_backpressure = io_sigsIn_backpressure; // @[MemInterfaceType.scala 108:30:@30210.4]
  assign io_in_x405_valid = _T_293 & io_sigsIn_backpressure; // @[sm_x420_inr_Foreach.scala 74:18:@30238.4]
  assign io_in_x405_bits_wdata_0 = x418_tuple[31:0]; // @[sm_x420_inr_Foreach.scala 75:26:@30240.4]
  assign io_in_x405_bits_wstrb = x418_tuple[32]; // @[sm_x420_inr_Foreach.scala 76:23:@30242.4]
  assign __io_b = $unsigned(io_sigsIn_cchainOutputs_0_counts_0); // @[Math.scala 721:17:@30193.4]
  assign RetimeWrapper_clock = clock; // @[:@30220.4]
  assign RetimeWrapper_reset = reset; // @[:@30221.4]
  assign RetimeWrapper_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30223.4]
  assign RetimeWrapper_io_in = ~ io_sigsIn_cchainOutputs_0_oobs_0; // @[package.scala 94:16:@30222.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30229.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30230.4]
  assign RetimeWrapper_1_io_flow = io_sigsIn_backpressure; // @[package.scala 95:18:@30232.4]
  assign RetimeWrapper_1_io_in = io_sigsIn_datapathEn; // @[package.scala 94:16:@30231.4]
endmodule
module x424_inr_UnitPipe_sm( // @[:@30398.2]
  input   clock, // @[:@30399.4]
  input   reset, // @[:@30400.4]
  input   io_enable, // @[:@30401.4]
  output  io_done, // @[:@30401.4]
  output  io_doneLatch, // @[:@30401.4]
  input   io_ctrDone, // @[:@30401.4]
  output  io_datapathEn, // @[:@30401.4]
  output  io_ctrInc, // @[:@30401.4]
  input   io_parentAck // @[:@30401.4]
);
  wire  active_clock; // @[Controllers.scala 261:22:@30403.4]
  wire  active_reset; // @[Controllers.scala 261:22:@30403.4]
  wire  active_io_input_set; // @[Controllers.scala 261:22:@30403.4]
  wire  active_io_input_reset; // @[Controllers.scala 261:22:@30403.4]
  wire  active_io_input_asyn_reset; // @[Controllers.scala 261:22:@30403.4]
  wire  active_io_output; // @[Controllers.scala 261:22:@30403.4]
  wire  done_clock; // @[Controllers.scala 262:20:@30406.4]
  wire  done_reset; // @[Controllers.scala 262:20:@30406.4]
  wire  done_io_input_set; // @[Controllers.scala 262:20:@30406.4]
  wire  done_io_input_reset; // @[Controllers.scala 262:20:@30406.4]
  wire  done_io_input_asyn_reset; // @[Controllers.scala 262:20:@30406.4]
  wire  done_io_output; // @[Controllers.scala 262:20:@30406.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30440.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30440.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30440.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30440.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30440.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30462.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30462.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30462.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30462.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30462.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30474.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30474.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30474.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30474.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30474.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30482.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30482.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30482.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30482.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30482.4]
  wire  _T_80; // @[Controllers.scala 264:48:@30411.4]
  wire  _T_81; // @[Controllers.scala 264:46:@30412.4]
  wire  _T_82; // @[Controllers.scala 264:62:@30413.4]
  wire  _T_100; // @[package.scala 100:49:@30431.4]
  reg  _T_103; // @[package.scala 48:56:@30432.4]
  reg [31:0] _RAND_0;
  wire  _T_118; // @[Controllers.scala 283:41:@30455.4]
  wire  _T_124; // @[package.scala 96:25:@30467.4 package.scala 96:25:@30468.4]
  wire  _T_126; // @[package.scala 100:49:@30469.4]
  reg  _T_129; // @[package.scala 48:56:@30470.4]
  reg [31:0] _RAND_1;
  reg  _T_146; // @[Controllers.scala 291:31:@30492.4]
  reg [31:0] _RAND_2;
  wire  _T_150; // @[package.scala 100:49:@30494.4]
  reg  _T_153; // @[package.scala 48:56:@30495.4]
  reg [31:0] _RAND_3;
  wire  _T_154; // @[package.scala 100:41:@30497.4]
  wire  _T_156; // @[Controllers.scala 292:61:@30498.4]
  wire  _T_157; // @[Controllers.scala 292:24:@30499.4]
  SRFF active ( // @[Controllers.scala 261:22:@30403.4]
    .clock(active_clock),
    .reset(active_reset),
    .io_input_set(active_io_input_set),
    .io_input_reset(active_io_input_reset),
    .io_input_asyn_reset(active_io_input_asyn_reset),
    .io_output(active_io_output)
  );
  SRFF done ( // @[Controllers.scala 262:20:@30406.4]
    .clock(done_clock),
    .reset(done_reset),
    .io_input_set(done_io_input_set),
    .io_input_reset(done_io_input_reset),
    .io_input_asyn_reset(done_io_input_asyn_reset),
    .io_output(done_io_output)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30440.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30462.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30474.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30482.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  assign _T_80 = ~ io_ctrDone; // @[Controllers.scala 264:48:@30411.4]
  assign _T_81 = io_enable & _T_80; // @[Controllers.scala 264:46:@30412.4]
  assign _T_82 = ~ done_io_output; // @[Controllers.scala 264:62:@30413.4]
  assign _T_100 = io_ctrDone == 1'h0; // @[package.scala 100:49:@30431.4]
  assign _T_118 = active_io_output & _T_82; // @[Controllers.scala 283:41:@30455.4]
  assign _T_124 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30467.4 package.scala 96:25:@30468.4]
  assign _T_126 = _T_124 == 1'h0; // @[package.scala 100:49:@30469.4]
  assign _T_150 = done_io_output == 1'h0; // @[package.scala 100:49:@30494.4]
  assign _T_154 = done_io_output & _T_153; // @[package.scala 100:41:@30497.4]
  assign _T_156 = _T_154 ? 1'h1 : _T_146; // @[Controllers.scala 292:61:@30498.4]
  assign _T_157 = io_parentAck ? 1'h0 : _T_156; // @[Controllers.scala 292:24:@30499.4]
  assign io_done = _T_124 & _T_129; // @[Controllers.scala 287:13:@30473.4]
  assign io_doneLatch = _T_146; // @[Controllers.scala 293:18:@30501.4]
  assign io_datapathEn = _T_118 & io_enable; // @[Controllers.scala 283:21:@30458.4]
  assign io_ctrInc = active_io_output & io_enable; // @[Controllers.scala 284:17:@30461.4]
  assign active_clock = clock; // @[:@30404.4]
  assign active_reset = reset; // @[:@30405.4]
  assign active_io_input_set = _T_81 & _T_82; // @[Controllers.scala 264:23:@30416.4]
  assign active_io_input_reset = io_ctrDone | io_parentAck; // @[Controllers.scala 265:25:@30420.4]
  assign active_io_input_asyn_reset = 1'h0; // @[Controllers.scala 266:30:@30421.4]
  assign done_clock = clock; // @[:@30407.4]
  assign done_reset = reset; // @[:@30408.4]
  assign done_io_input_set = io_ctrDone & _T_103; // @[Controllers.scala 269:104:@30436.4]
  assign done_io_input_reset = io_parentAck; // @[Controllers.scala 267:23:@30429.4]
  assign done_io_input_asyn_reset = 1'h0; // @[Controllers.scala 268:28:@30430.4]
  assign RetimeWrapper_clock = clock; // @[:@30441.4]
  assign RetimeWrapper_reset = reset; // @[:@30442.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30444.4]
  assign RetimeWrapper_io_in = done_io_output; // @[package.scala 94:16:@30443.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30463.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30464.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30466.4]
  assign RetimeWrapper_1_io_in = done_io_output; // @[package.scala 94:16:@30465.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30475.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30476.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30478.4]
  assign RetimeWrapper_2_io_in = 1'h0; // @[package.scala 94:16:@30477.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30483.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30484.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30486.4]
  assign RetimeWrapper_3_io_in = io_ctrDone; // @[package.scala 94:16:@30485.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_103 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_129 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_146 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_153 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_103 <= 1'h0;
    end else begin
      _T_103 <= _T_100;
    end
    if (reset) begin
      _T_129 <= 1'h0;
    end else begin
      _T_129 <= _T_126;
    end
    if (reset) begin
      _T_146 <= 1'h0;
    end else begin
      if (io_parentAck) begin
        _T_146 <= 1'h0;
      end else begin
        if (_T_154) begin
          _T_146 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_153 <= 1'h0;
    end else begin
      _T_153 <= _T_150;
    end
  end
endmodule
module x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1( // @[:@30576.2]
  output  io_in_x406_ready, // @[:@30579.4]
  input   io_sigsIn_datapathEn // @[:@30579.4]
);
  assign io_in_x406_ready = io_sigsIn_datapathEn; // @[sm_x424_inr_UnitPipe.scala 57:18:@30591.4]
endmodule
module x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1( // @[:@30594.2]
  input         clock, // @[:@30595.4]
  input         reset, // @[:@30596.4]
  input         io_in_x404_ready, // @[:@30597.4]
  output        io_in_x404_valid, // @[:@30597.4]
  output [63:0] io_in_x404_bits_addr, // @[:@30597.4]
  output [31:0] io_in_x404_bits_size, // @[:@30597.4]
  output        io_in_x406_ready, // @[:@30597.4]
  input         io_in_x406_valid, // @[:@30597.4]
  input  [63:0] io_in_x219_outdram_number, // @[:@30597.4]
  output [20:0] io_in_x223_outbuf_0_rPort_0_ofs_0, // @[:@30597.4]
  output        io_in_x223_outbuf_0_rPort_0_en_0, // @[:@30597.4]
  output        io_in_x223_outbuf_0_rPort_0_backpressure, // @[:@30597.4]
  input  [31:0] io_in_x223_outbuf_0_rPort_0_output_0, // @[:@30597.4]
  input         io_in_x405_ready, // @[:@30597.4]
  output        io_in_x405_valid, // @[:@30597.4]
  output [31:0] io_in_x405_bits_wdata_0, // @[:@30597.4]
  output        io_in_x405_bits_wstrb, // @[:@30597.4]
  input         io_sigsIn_smEnableOuts_0, // @[:@30597.4]
  input         io_sigsIn_smEnableOuts_1, // @[:@30597.4]
  input         io_sigsIn_smEnableOuts_2, // @[:@30597.4]
  input         io_sigsIn_smChildAcks_0, // @[:@30597.4]
  input         io_sigsIn_smChildAcks_1, // @[:@30597.4]
  input         io_sigsIn_smChildAcks_2, // @[:@30597.4]
  output        io_sigsOut_smDoneIn_0, // @[:@30597.4]
  output        io_sigsOut_smDoneIn_1, // @[:@30597.4]
  output        io_sigsOut_smDoneIn_2, // @[:@30597.4]
  output        io_sigsOut_smCtrCopyDone_0, // @[:@30597.4]
  output        io_sigsOut_smCtrCopyDone_1, // @[:@30597.4]
  output        io_sigsOut_smCtrCopyDone_2, // @[:@30597.4]
  input         io_rr // @[:@30597.4]
);
  wire  x411_inr_UnitPipe_sm_clock; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_reset; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_io_enable; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_io_done; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_io_doneLatch; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_io_ctrDone; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_io_datapathEn; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_io_ctrInc; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_io_parentAck; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  x411_inr_UnitPipe_sm_io_backpressure; // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@30721.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@30721.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@30721.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@30721.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@30721.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@30729.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@30729.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@30729.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@30729.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@30729.4]
  wire  x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_valid; // @[sm_x411_inr_UnitPipe.scala 69:24:@30759.4]
  wire [63:0] x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_bits_addr; // @[sm_x411_inr_UnitPipe.scala 69:24:@30759.4]
  wire [31:0] x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_bits_size; // @[sm_x411_inr_UnitPipe.scala 69:24:@30759.4]
  wire [63:0] x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x219_outdram_number; // @[sm_x411_inr_UnitPipe.scala 69:24:@30759.4]
  wire  x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_sigsIn_backpressure; // @[sm_x411_inr_UnitPipe.scala 69:24:@30759.4]
  wire  x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x411_inr_UnitPipe.scala 69:24:@30759.4]
  wire  x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_rr; // @[sm_x411_inr_UnitPipe.scala 69:24:@30759.4]
  wire  x413_ctrchain_clock; // @[SpatialBlocks.scala 37:22:@30827.4]
  wire  x413_ctrchain_reset; // @[SpatialBlocks.scala 37:22:@30827.4]
  wire  x413_ctrchain_io_input_reset; // @[SpatialBlocks.scala 37:22:@30827.4]
  wire  x413_ctrchain_io_input_enable; // @[SpatialBlocks.scala 37:22:@30827.4]
  wire [22:0] x413_ctrchain_io_output_counts_0; // @[SpatialBlocks.scala 37:22:@30827.4]
  wire  x413_ctrchain_io_output_oobs_0; // @[SpatialBlocks.scala 37:22:@30827.4]
  wire  x413_ctrchain_io_output_done; // @[SpatialBlocks.scala 37:22:@30827.4]
  wire  x420_inr_Foreach_sm_clock; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_reset; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_enable; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_done; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_doneLatch; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_ctrDone; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_datapathEn; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_ctrInc; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_ctrRst; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_parentAck; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_backpressure; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  x420_inr_Foreach_sm_io_break; // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@30908.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@30948.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@30948.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@30948.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@30948.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@30948.4]
  wire  RetimeWrapper_4_clock; // @[package.scala 93:22:@30956.4]
  wire  RetimeWrapper_4_reset; // @[package.scala 93:22:@30956.4]
  wire  RetimeWrapper_4_io_flow; // @[package.scala 93:22:@30956.4]
  wire  RetimeWrapper_4_io_in; // @[package.scala 93:22:@30956.4]
  wire  RetimeWrapper_4_io_out; // @[package.scala 93:22:@30956.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_clock; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_reset; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire [20:0] x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_en_0; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire [31:0] x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_output_0; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_valid; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire [31:0] x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_bits_wdata_0; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_bits_wstrb; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_backpressure; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_datapathEn; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_break; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire [31:0] x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_rr; // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
  wire  x424_inr_UnitPipe_sm_clock; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  x424_inr_UnitPipe_sm_reset; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  x424_inr_UnitPipe_sm_io_enable; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  x424_inr_UnitPipe_sm_io_done; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  x424_inr_UnitPipe_sm_io_doneLatch; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  x424_inr_UnitPipe_sm_io_ctrDone; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  x424_inr_UnitPipe_sm_io_datapathEn; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  x424_inr_UnitPipe_sm_io_ctrInc; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  x424_inr_UnitPipe_sm_io_parentAck; // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
  wire  RetimeWrapper_5_clock; // @[package.scala 93:22:@31168.4]
  wire  RetimeWrapper_5_reset; // @[package.scala 93:22:@31168.4]
  wire  RetimeWrapper_5_io_flow; // @[package.scala 93:22:@31168.4]
  wire  RetimeWrapper_5_io_in; // @[package.scala 93:22:@31168.4]
  wire  RetimeWrapper_5_io_out; // @[package.scala 93:22:@31168.4]
  wire  RetimeWrapper_6_clock; // @[package.scala 93:22:@31176.4]
  wire  RetimeWrapper_6_reset; // @[package.scala 93:22:@31176.4]
  wire  RetimeWrapper_6_io_flow; // @[package.scala 93:22:@31176.4]
  wire  RetimeWrapper_6_io_in; // @[package.scala 93:22:@31176.4]
  wire  RetimeWrapper_6_io_out; // @[package.scala 93:22:@31176.4]
  wire  x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1_io_in_x406_ready; // @[sm_x424_inr_UnitPipe.scala 60:24:@31206.4]
  wire  x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1_io_sigsIn_datapathEn; // @[sm_x424_inr_UnitPipe.scala 60:24:@31206.4]
  wire  _T_359; // @[package.scala 100:49:@30692.4]
  reg  _T_362; // @[package.scala 48:56:@30693.4]
  reg [31:0] _RAND_0;
  wire  _T_375; // @[package.scala 96:25:@30726.4 package.scala 96:25:@30727.4]
  wire  _T_381; // @[package.scala 96:25:@30734.4 package.scala 96:25:@30735.4]
  wire  _T_384; // @[SpatialBlocks.scala 138:93:@30737.4]
  wire  _T_454; // @[package.scala 96:25:@30913.4 package.scala 96:25:@30914.4]
  wire  _T_468; // @[package.scala 96:25:@30953.4 package.scala 96:25:@30954.4]
  wire  _T_474; // @[package.scala 96:25:@30961.4 package.scala 96:25:@30962.4]
  wire  _T_477; // @[SpatialBlocks.scala 138:93:@30964.4]
  wire  _T_479; // @[SpatialBlocks.scala 157:36:@30973.4]
  wire  _T_480; // @[SpatialBlocks.scala 157:78:@30974.4]
  wire  _T_547; // @[package.scala 100:49:@31139.4]
  reg  _T_550; // @[package.scala 48:56:@31140.4]
  reg [31:0] _RAND_1;
  wire  x424_inr_UnitPipe_sigsIn_forwardpressure; // @[sm_x425_outr_UnitPipe.scala 101:55:@31146.4]
  wire  _T_563; // @[package.scala 96:25:@31173.4 package.scala 96:25:@31174.4]
  wire  _T_569; // @[package.scala 96:25:@31181.4 package.scala 96:25:@31182.4]
  wire  _T_572; // @[SpatialBlocks.scala 138:93:@31184.4]
  wire  x424_inr_UnitPipe_sigsIn_baseEn; // @[SpatialBlocks.scala 138:90:@31185.4]
  x411_inr_UnitPipe_sm x411_inr_UnitPipe_sm ( // @[sm_x411_inr_UnitPipe.scala 33:18:@30664.4]
    .clock(x411_inr_UnitPipe_sm_clock),
    .reset(x411_inr_UnitPipe_sm_reset),
    .io_enable(x411_inr_UnitPipe_sm_io_enable),
    .io_done(x411_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x411_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x411_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x411_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x411_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x411_inr_UnitPipe_sm_io_parentAck),
    .io_backpressure(x411_inr_UnitPipe_sm_io_backpressure)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@30721.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@30729.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1 x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1 ( // @[sm_x411_inr_UnitPipe.scala 69:24:@30759.4]
    .io_in_x404_valid(x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_valid),
    .io_in_x404_bits_addr(x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_bits_addr),
    .io_in_x404_bits_size(x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_bits_size),
    .io_in_x219_outdram_number(x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x219_outdram_number),
    .io_sigsIn_backpressure(x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_sigsIn_datapathEn),
    .io_rr(x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_rr)
  );
  x413_ctrchain x413_ctrchain ( // @[SpatialBlocks.scala 37:22:@30827.4]
    .clock(x413_ctrchain_clock),
    .reset(x413_ctrchain_reset),
    .io_input_reset(x413_ctrchain_io_input_reset),
    .io_input_enable(x413_ctrchain_io_input_enable),
    .io_output_counts_0(x413_ctrchain_io_output_counts_0),
    .io_output_oobs_0(x413_ctrchain_io_output_oobs_0),
    .io_output_done(x413_ctrchain_io_output_done)
  );
  x420_inr_Foreach_sm x420_inr_Foreach_sm ( // @[sm_x420_inr_Foreach.scala 33:18:@30880.4]
    .clock(x420_inr_Foreach_sm_clock),
    .reset(x420_inr_Foreach_sm_reset),
    .io_enable(x420_inr_Foreach_sm_io_enable),
    .io_done(x420_inr_Foreach_sm_io_done),
    .io_doneLatch(x420_inr_Foreach_sm_io_doneLatch),
    .io_ctrDone(x420_inr_Foreach_sm_io_ctrDone),
    .io_datapathEn(x420_inr_Foreach_sm_io_datapathEn),
    .io_ctrInc(x420_inr_Foreach_sm_io_ctrInc),
    .io_ctrRst(x420_inr_Foreach_sm_io_ctrRst),
    .io_parentAck(x420_inr_Foreach_sm_io_parentAck),
    .io_backpressure(x420_inr_Foreach_sm_io_backpressure),
    .io_break(x420_inr_Foreach_sm_io_break)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@30908.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@30948.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  RetimeWrapper RetimeWrapper_4 ( // @[package.scala 93:22:@30956.4]
    .clock(RetimeWrapper_4_clock),
    .reset(RetimeWrapper_4_reset),
    .io_flow(RetimeWrapper_4_io_flow),
    .io_in(RetimeWrapper_4_io_in),
    .io_out(RetimeWrapper_4_io_out)
  );
  x420_inr_Foreach_kernelx420_inr_Foreach_concrete1 x420_inr_Foreach_kernelx420_inr_Foreach_concrete1 ( // @[sm_x420_inr_Foreach.scala 78:24:@30991.4]
    .clock(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_clock),
    .reset(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_reset),
    .io_in_x223_outbuf_0_rPort_0_ofs_0(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0),
    .io_in_x223_outbuf_0_rPort_0_en_0(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_en_0),
    .io_in_x223_outbuf_0_rPort_0_backpressure(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure),
    .io_in_x223_outbuf_0_rPort_0_output_0(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_output_0),
    .io_in_x405_valid(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_valid),
    .io_in_x405_bits_wdata_0(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_bits_wdata_0),
    .io_in_x405_bits_wstrb(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_bits_wstrb),
    .io_sigsIn_backpressure(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_backpressure),
    .io_sigsIn_datapathEn(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_datapathEn),
    .io_sigsIn_break(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_break),
    .io_sigsIn_cchainOutputs_0_counts_0(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0),
    .io_sigsIn_cchainOutputs_0_oobs_0(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0),
    .io_rr(x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_rr)
  );
  x424_inr_UnitPipe_sm x424_inr_UnitPipe_sm ( // @[sm_x424_inr_UnitPipe.scala 32:18:@31111.4]
    .clock(x424_inr_UnitPipe_sm_clock),
    .reset(x424_inr_UnitPipe_sm_reset),
    .io_enable(x424_inr_UnitPipe_sm_io_enable),
    .io_done(x424_inr_UnitPipe_sm_io_done),
    .io_doneLatch(x424_inr_UnitPipe_sm_io_doneLatch),
    .io_ctrDone(x424_inr_UnitPipe_sm_io_ctrDone),
    .io_datapathEn(x424_inr_UnitPipe_sm_io_datapathEn),
    .io_ctrInc(x424_inr_UnitPipe_sm_io_ctrInc),
    .io_parentAck(x424_inr_UnitPipe_sm_io_parentAck)
  );
  RetimeWrapper RetimeWrapper_5 ( // @[package.scala 93:22:@31168.4]
    .clock(RetimeWrapper_5_clock),
    .reset(RetimeWrapper_5_reset),
    .io_flow(RetimeWrapper_5_io_flow),
    .io_in(RetimeWrapper_5_io_in),
    .io_out(RetimeWrapper_5_io_out)
  );
  RetimeWrapper RetimeWrapper_6 ( // @[package.scala 93:22:@31176.4]
    .clock(RetimeWrapper_6_clock),
    .reset(RetimeWrapper_6_reset),
    .io_flow(RetimeWrapper_6_io_flow),
    .io_in(RetimeWrapper_6_io_in),
    .io_out(RetimeWrapper_6_io_out)
  );
  x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1 x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1 ( // @[sm_x424_inr_UnitPipe.scala 60:24:@31206.4]
    .io_in_x406_ready(x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1_io_in_x406_ready),
    .io_sigsIn_datapathEn(x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1_io_sigsIn_datapathEn)
  );
  assign _T_359 = x411_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@30692.4]
  assign _T_375 = RetimeWrapper_io_out; // @[package.scala 96:25:@30726.4 package.scala 96:25:@30727.4]
  assign _T_381 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@30734.4 package.scala 96:25:@30735.4]
  assign _T_384 = ~ _T_381; // @[SpatialBlocks.scala 138:93:@30737.4]
  assign _T_454 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@30913.4 package.scala 96:25:@30914.4]
  assign _T_468 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@30953.4 package.scala 96:25:@30954.4]
  assign _T_474 = RetimeWrapper_4_io_out; // @[package.scala 96:25:@30961.4 package.scala 96:25:@30962.4]
  assign _T_477 = ~ _T_474; // @[SpatialBlocks.scala 138:93:@30964.4]
  assign _T_479 = x420_inr_Foreach_sm_io_datapathEn; // @[SpatialBlocks.scala 157:36:@30973.4]
  assign _T_480 = ~ x420_inr_Foreach_sm_io_ctrDone; // @[SpatialBlocks.scala 157:78:@30974.4]
  assign _T_547 = x424_inr_UnitPipe_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@31139.4]
  assign x424_inr_UnitPipe_sigsIn_forwardpressure = io_in_x406_valid | x424_inr_UnitPipe_sm_io_doneLatch; // @[sm_x425_outr_UnitPipe.scala 101:55:@31146.4]
  assign _T_563 = RetimeWrapper_5_io_out; // @[package.scala 96:25:@31173.4 package.scala 96:25:@31174.4]
  assign _T_569 = RetimeWrapper_6_io_out; // @[package.scala 96:25:@31181.4 package.scala 96:25:@31182.4]
  assign _T_572 = ~ _T_569; // @[SpatialBlocks.scala 138:93:@31184.4]
  assign x424_inr_UnitPipe_sigsIn_baseEn = _T_563 & _T_572; // @[SpatialBlocks.scala 138:90:@31185.4]
  assign io_in_x404_valid = x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_valid; // @[sm_x411_inr_UnitPipe.scala 49:23:@30797.4]
  assign io_in_x404_bits_addr = x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_bits_addr; // @[sm_x411_inr_UnitPipe.scala 49:23:@30796.4]
  assign io_in_x404_bits_size = x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x404_bits_size; // @[sm_x411_inr_UnitPipe.scala 49:23:@30795.4]
  assign io_in_x406_ready = x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1_io_in_x406_ready; // @[sm_x424_inr_UnitPipe.scala 46:23:@31242.4]
  assign io_in_x223_outbuf_0_rPort_0_ofs_0 = x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@31042.4]
  assign io_in_x223_outbuf_0_rPort_0_en_0 = x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@31041.4]
  assign io_in_x223_outbuf_0_rPort_0_backpressure = x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@31040.4]
  assign io_in_x405_valid = x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_valid; // @[sm_x420_inr_Foreach.scala 50:23:@31046.4]
  assign io_in_x405_bits_wdata_0 = x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_bits_wdata_0; // @[sm_x420_inr_Foreach.scala 50:23:@31045.4]
  assign io_in_x405_bits_wstrb = x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x405_bits_wstrb; // @[sm_x420_inr_Foreach.scala 50:23:@31044.4]
  assign io_sigsOut_smDoneIn_0 = x411_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@30744.4]
  assign io_sigsOut_smDoneIn_1 = x420_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 156:53:@30971.4]
  assign io_sigsOut_smDoneIn_2 = x424_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@31191.4]
  assign io_sigsOut_smCtrCopyDone_0 = x411_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@30758.4]
  assign io_sigsOut_smCtrCopyDone_1 = x420_inr_Foreach_sm_io_done; // @[SpatialBlocks.scala 168:125:@30990.4]
  assign io_sigsOut_smCtrCopyDone_2 = x424_inr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 168:125:@31205.4]
  assign x411_inr_UnitPipe_sm_clock = clock; // @[:@30665.4]
  assign x411_inr_UnitPipe_sm_reset = reset; // @[:@30666.4]
  assign x411_inr_UnitPipe_sm_io_enable = _T_375 & _T_384; // @[SpatialBlocks.scala 140:18:@30741.4]
  assign x411_inr_UnitPipe_sm_io_ctrDone = x411_inr_UnitPipe_sm_io_ctrInc & _T_362; // @[sm_x425_outr_UnitPipe.scala 77:39:@30696.4]
  assign x411_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@30743.4]
  assign x411_inr_UnitPipe_sm_io_backpressure = io_in_x404_ready | x411_inr_UnitPipe_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@30715.4]
  assign RetimeWrapper_clock = clock; // @[:@30722.4]
  assign RetimeWrapper_reset = reset; // @[:@30723.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@30725.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@30724.4]
  assign RetimeWrapper_1_clock = clock; // @[:@30730.4]
  assign RetimeWrapper_1_reset = reset; // @[:@30731.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@30733.4]
  assign RetimeWrapper_1_io_in = x411_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@30732.4]
  assign x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_in_x219_outdram_number = io_in_x219_outdram_number; // @[sm_x411_inr_UnitPipe.scala 50:31:@30799.4]
  assign x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_sigsIn_backpressure = io_in_x404_ready | x411_inr_UnitPipe_sm_io_doneLatch; // @[sm_x411_inr_UnitPipe.scala 74:22:@30814.4]
  assign x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x411_inr_UnitPipe_sm_io_datapathEn; // @[sm_x411_inr_UnitPipe.scala 74:22:@30812.4]
  assign x411_inr_UnitPipe_kernelx411_inr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x411_inr_UnitPipe.scala 73:18:@30800.4]
  assign x413_ctrchain_clock = clock; // @[:@30828.4]
  assign x413_ctrchain_reset = reset; // @[:@30829.4]
  assign x413_ctrchain_io_input_reset = x420_inr_Foreach_sm_io_ctrRst; // @[SpatialBlocks.scala 159:100:@30989.4]
  assign x413_ctrchain_io_input_enable = x420_inr_Foreach_sm_io_ctrInc; // @[SpatialBlocks.scala 132:75:@30941.4 SpatialBlocks.scala 159:42:@30988.4]
  assign x420_inr_Foreach_sm_clock = clock; // @[:@30881.4]
  assign x420_inr_Foreach_sm_reset = reset; // @[:@30882.4]
  assign x420_inr_Foreach_sm_io_enable = _T_468 & _T_477; // @[SpatialBlocks.scala 140:18:@30968.4]
  assign x420_inr_Foreach_sm_io_ctrDone = io_rr ? _T_454 : 1'h0; // @[sm_x425_outr_UnitPipe.scala 90:38:@30916.4]
  assign x420_inr_Foreach_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@30970.4]
  assign x420_inr_Foreach_sm_io_backpressure = io_in_x405_ready | x420_inr_Foreach_sm_io_doneLatch; // @[SpatialBlocks.scala 133:24:@30942.4]
  assign x420_inr_Foreach_sm_io_break = 1'h0; // @[sm_x425_outr_UnitPipe.scala 94:36:@30922.4]
  assign RetimeWrapper_2_clock = clock; // @[:@30909.4]
  assign RetimeWrapper_2_reset = reset; // @[:@30910.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@30912.4]
  assign RetimeWrapper_2_io_in = x413_ctrchain_io_output_done; // @[package.scala 94:16:@30911.4]
  assign RetimeWrapper_3_clock = clock; // @[:@30949.4]
  assign RetimeWrapper_3_reset = reset; // @[:@30950.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@30952.4]
  assign RetimeWrapper_3_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@30951.4]
  assign RetimeWrapper_4_clock = clock; // @[:@30957.4]
  assign RetimeWrapper_4_reset = reset; // @[:@30958.4]
  assign RetimeWrapper_4_io_flow = 1'h1; // @[package.scala 95:18:@30960.4]
  assign RetimeWrapper_4_io_in = x420_inr_Foreach_sm_io_done; // @[package.scala 94:16:@30959.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_clock = clock; // @[:@30992.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_reset = reset; // @[:@30993.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_in_x223_outbuf_0_rPort_0_output_0 = io_in_x223_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@31039.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_backpressure = io_in_x405_ready | x420_inr_Foreach_sm_io_doneLatch; // @[sm_x420_inr_Foreach.scala 83:22:@31062.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_datapathEn = _T_479 & _T_480; // @[sm_x420_inr_Foreach.scala 83:22:@31060.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_break = x420_inr_Foreach_sm_io_break; // @[sm_x420_inr_Foreach.scala 83:22:@31058.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_counts_0 = {{9{x413_ctrchain_io_output_counts_0[22]}},x413_ctrchain_io_output_counts_0}; // @[sm_x420_inr_Foreach.scala 83:22:@31053.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_sigsIn_cchainOutputs_0_oobs_0 = x413_ctrchain_io_output_oobs_0; // @[sm_x420_inr_Foreach.scala 83:22:@31052.4]
  assign x420_inr_Foreach_kernelx420_inr_Foreach_concrete1_io_rr = io_rr; // @[sm_x420_inr_Foreach.scala 82:18:@31048.4]
  assign x424_inr_UnitPipe_sm_clock = clock; // @[:@31112.4]
  assign x424_inr_UnitPipe_sm_reset = reset; // @[:@31113.4]
  assign x424_inr_UnitPipe_sm_io_enable = x424_inr_UnitPipe_sigsIn_baseEn & x424_inr_UnitPipe_sigsIn_forwardpressure; // @[SpatialBlocks.scala 140:18:@31188.4]
  assign x424_inr_UnitPipe_sm_io_ctrDone = x424_inr_UnitPipe_sm_io_ctrInc & _T_550; // @[sm_x425_outr_UnitPipe.scala 99:39:@31143.4]
  assign x424_inr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_2; // @[SpatialBlocks.scala 142:21:@31190.4]
  assign RetimeWrapper_5_clock = clock; // @[:@31169.4]
  assign RetimeWrapper_5_reset = reset; // @[:@31170.4]
  assign RetimeWrapper_5_io_flow = 1'h1; // @[package.scala 95:18:@31172.4]
  assign RetimeWrapper_5_io_in = io_sigsIn_smEnableOuts_2; // @[package.scala 94:16:@31171.4]
  assign RetimeWrapper_6_clock = clock; // @[:@31177.4]
  assign RetimeWrapper_6_reset = reset; // @[:@31178.4]
  assign RetimeWrapper_6_io_flow = 1'h1; // @[package.scala 95:18:@31180.4]
  assign RetimeWrapper_6_io_in = x424_inr_UnitPipe_sm_io_done; // @[package.scala 94:16:@31179.4]
  assign x424_inr_UnitPipe_kernelx424_inr_UnitPipe_concrete1_io_sigsIn_datapathEn = x424_inr_UnitPipe_sm_io_datapathEn; // @[sm_x424_inr_UnitPipe.scala 65:22:@31255.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_362 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_550 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_362 <= 1'h0;
    end else begin
      _T_362 <= _T_359;
    end
    if (reset) begin
      _T_550 <= 1'h0;
    end else begin
      _T_550 <= _T_547;
    end
  end
endmodule
module x478_kernelx478_concrete1( // @[:@31271.2]
  input          clock, // @[:@31272.4]
  input          reset, // @[:@31273.4]
  input          io_in_x404_ready, // @[:@31274.4]
  output         io_in_x404_valid, // @[:@31274.4]
  output [63:0]  io_in_x404_bits_addr, // @[:@31274.4]
  output [31:0]  io_in_x404_bits_size, // @[:@31274.4]
  input          io_in_x221_TVALID, // @[:@31274.4]
  output         io_in_x221_TREADY, // @[:@31274.4]
  input  [255:0] io_in_x221_TDATA, // @[:@31274.4]
  input  [7:0]   io_in_x221_TID, // @[:@31274.4]
  input  [7:0]   io_in_x221_TDEST, // @[:@31274.4]
  output         io_in_x406_ready, // @[:@31274.4]
  input          io_in_x406_valid, // @[:@31274.4]
  input  [63:0]  io_in_x219_outdram_number, // @[:@31274.4]
  output [20:0]  io_in_x223_outbuf_0_rPort_0_ofs_0, // @[:@31274.4]
  output         io_in_x223_outbuf_0_rPort_0_en_0, // @[:@31274.4]
  output         io_in_x223_outbuf_0_rPort_0_backpressure, // @[:@31274.4]
  input  [31:0]  io_in_x223_outbuf_0_rPort_0_output_0, // @[:@31274.4]
  input          io_in_x405_ready, // @[:@31274.4]
  output         io_in_x405_valid, // @[:@31274.4]
  output [31:0]  io_in_x405_bits_wdata_0, // @[:@31274.4]
  output         io_in_x405_bits_wstrb, // @[:@31274.4]
  output         io_in_x222_TVALID, // @[:@31274.4]
  input          io_in_x222_TREADY, // @[:@31274.4]
  output [255:0] io_in_x222_TDATA, // @[:@31274.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@31274.4]
  input          io_sigsIn_smEnableOuts_1, // @[:@31274.4]
  input          io_sigsIn_smChildAcks_0, // @[:@31274.4]
  input          io_sigsIn_smChildAcks_1, // @[:@31274.4]
  output         io_sigsOut_smDoneIn_0, // @[:@31274.4]
  output         io_sigsOut_smDoneIn_1, // @[:@31274.4]
  input          io_rr // @[:@31274.4]
);
  wire  x403_outr_UnitPipe_sm_clock; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_reset; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_enable; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_done; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_parentAck; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_childAck_0; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_childAck_1; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  x403_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@31409.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@31409.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@31409.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@31409.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@31409.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@31417.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@31417.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@31417.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@31417.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@31417.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_clock; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_reset; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TVALID; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TREADY; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire [255:0] x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TDATA; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire [7:0] x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TID; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire [7:0] x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TDEST; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TVALID; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TREADY; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire [255:0] x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TDATA; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_rr; // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
  wire  x425_outr_UnitPipe_sm_clock; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_reset; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_enable; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_done; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_parentAck; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_doneIn_0; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_doneIn_1; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_doneIn_2; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_childAck_0; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_childAck_1; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_childAck_2; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_ctrCopyDone_0; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_ctrCopyDone_1; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  x425_outr_UnitPipe_sm_io_ctrCopyDone_2; // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
  wire  RetimeWrapper_2_clock; // @[package.scala 93:22:@31698.4]
  wire  RetimeWrapper_2_reset; // @[package.scala 93:22:@31698.4]
  wire  RetimeWrapper_2_io_flow; // @[package.scala 93:22:@31698.4]
  wire  RetimeWrapper_2_io_in; // @[package.scala 93:22:@31698.4]
  wire  RetimeWrapper_2_io_out; // @[package.scala 93:22:@31698.4]
  wire  RetimeWrapper_3_clock; // @[package.scala 93:22:@31706.4]
  wire  RetimeWrapper_3_reset; // @[package.scala 93:22:@31706.4]
  wire  RetimeWrapper_3_io_flow; // @[package.scala 93:22:@31706.4]
  wire  RetimeWrapper_3_io_in; // @[package.scala 93:22:@31706.4]
  wire  RetimeWrapper_3_io_out; // @[package.scala 93:22:@31706.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_clock; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_reset; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_ready; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_valid; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire [63:0] x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_bits_addr; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire [31:0] x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_bits_size; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x406_ready; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x406_valid; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire [63:0] x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x219_outdram_number; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire [20:0] x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_en_0; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire [31:0] x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_output_0; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_ready; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_valid; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire [31:0] x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_bits_wdata_0; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_bits_wstrb; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_rr; // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
  wire  _T_408; // @[package.scala 96:25:@31414.4 package.scala 96:25:@31415.4]
  wire  _T_414; // @[package.scala 96:25:@31422.4 package.scala 96:25:@31423.4]
  wire  _T_417; // @[SpatialBlocks.scala 138:93:@31425.4]
  wire  _T_508; // @[package.scala 96:25:@31703.4 package.scala 96:25:@31704.4]
  wire  _T_514; // @[package.scala 96:25:@31711.4 package.scala 96:25:@31712.4]
  wire  _T_517; // @[SpatialBlocks.scala 138:93:@31714.4]
  x403_outr_UnitPipe_sm x403_outr_UnitPipe_sm ( // @[sm_x403_outr_UnitPipe.scala 32:18:@31347.4]
    .clock(x403_outr_UnitPipe_sm_clock),
    .reset(x403_outr_UnitPipe_sm_reset),
    .io_enable(x403_outr_UnitPipe_sm_io_enable),
    .io_done(x403_outr_UnitPipe_sm_io_done),
    .io_parentAck(x403_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x403_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x403_outr_UnitPipe_sm_io_doneIn_1),
    .io_enableOut_0(x403_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x403_outr_UnitPipe_sm_io_enableOut_1),
    .io_childAck_0(x403_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x403_outr_UnitPipe_sm_io_childAck_1),
    .io_ctrCopyDone_0(x403_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x403_outr_UnitPipe_sm_io_ctrCopyDone_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@31409.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@31417.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1 x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1 ( // @[sm_x403_outr_UnitPipe.scala 87:24:@31448.4]
    .clock(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_clock),
    .reset(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_reset),
    .io_in_x221_TVALID(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TVALID),
    .io_in_x221_TREADY(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TREADY),
    .io_in_x221_TDATA(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TDATA),
    .io_in_x221_TID(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TID),
    .io_in_x221_TDEST(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TDEST),
    .io_in_x222_TVALID(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TVALID),
    .io_in_x222_TREADY(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TREADY),
    .io_in_x222_TDATA(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TDATA),
    .io_sigsIn_smEnableOuts_0(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smCtrCopyDone_0(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_rr(x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_rr)
  );
  x425_outr_UnitPipe_sm x425_outr_UnitPipe_sm ( // @[sm_x425_outr_UnitPipe.scala 36:18:@31626.4]
    .clock(x425_outr_UnitPipe_sm_clock),
    .reset(x425_outr_UnitPipe_sm_reset),
    .io_enable(x425_outr_UnitPipe_sm_io_enable),
    .io_done(x425_outr_UnitPipe_sm_io_done),
    .io_parentAck(x425_outr_UnitPipe_sm_io_parentAck),
    .io_doneIn_0(x425_outr_UnitPipe_sm_io_doneIn_0),
    .io_doneIn_1(x425_outr_UnitPipe_sm_io_doneIn_1),
    .io_doneIn_2(x425_outr_UnitPipe_sm_io_doneIn_2),
    .io_enableOut_0(x425_outr_UnitPipe_sm_io_enableOut_0),
    .io_enableOut_1(x425_outr_UnitPipe_sm_io_enableOut_1),
    .io_enableOut_2(x425_outr_UnitPipe_sm_io_enableOut_2),
    .io_childAck_0(x425_outr_UnitPipe_sm_io_childAck_0),
    .io_childAck_1(x425_outr_UnitPipe_sm_io_childAck_1),
    .io_childAck_2(x425_outr_UnitPipe_sm_io_childAck_2),
    .io_ctrCopyDone_0(x425_outr_UnitPipe_sm_io_ctrCopyDone_0),
    .io_ctrCopyDone_1(x425_outr_UnitPipe_sm_io_ctrCopyDone_1),
    .io_ctrCopyDone_2(x425_outr_UnitPipe_sm_io_ctrCopyDone_2)
  );
  RetimeWrapper RetimeWrapper_2 ( // @[package.scala 93:22:@31698.4]
    .clock(RetimeWrapper_2_clock),
    .reset(RetimeWrapper_2_reset),
    .io_flow(RetimeWrapper_2_io_flow),
    .io_in(RetimeWrapper_2_io_in),
    .io_out(RetimeWrapper_2_io_out)
  );
  RetimeWrapper RetimeWrapper_3 ( // @[package.scala 93:22:@31706.4]
    .clock(RetimeWrapper_3_clock),
    .reset(RetimeWrapper_3_reset),
    .io_flow(RetimeWrapper_3_io_flow),
    .io_in(RetimeWrapper_3_io_in),
    .io_out(RetimeWrapper_3_io_out)
  );
  x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1 x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1 ( // @[sm_x425_outr_UnitPipe.scala 108:24:@31738.4]
    .clock(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_clock),
    .reset(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_reset),
    .io_in_x404_ready(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_ready),
    .io_in_x404_valid(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_valid),
    .io_in_x404_bits_addr(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_bits_addr),
    .io_in_x404_bits_size(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_bits_size),
    .io_in_x406_ready(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x406_ready),
    .io_in_x406_valid(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x406_valid),
    .io_in_x219_outdram_number(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x219_outdram_number),
    .io_in_x223_outbuf_0_rPort_0_ofs_0(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0),
    .io_in_x223_outbuf_0_rPort_0_en_0(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_en_0),
    .io_in_x223_outbuf_0_rPort_0_backpressure(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure),
    .io_in_x223_outbuf_0_rPort_0_output_0(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_output_0),
    .io_in_x405_ready(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_ready),
    .io_in_x405_valid(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_valid),
    .io_in_x405_bits_wdata_0(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_bits_wdata_0),
    .io_in_x405_bits_wstrb(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_bits_wstrb),
    .io_sigsIn_smEnableOuts_0(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smEnableOuts_2(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2),
    .io_sigsIn_smChildAcks_0(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsIn_smChildAcks_2(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2),
    .io_sigsOut_smDoneIn_0(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1),
    .io_sigsOut_smDoneIn_2(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2),
    .io_sigsOut_smCtrCopyDone_0(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0),
    .io_sigsOut_smCtrCopyDone_1(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1),
    .io_sigsOut_smCtrCopyDone_2(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2),
    .io_rr(x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_rr)
  );
  assign _T_408 = RetimeWrapper_io_out; // @[package.scala 96:25:@31414.4 package.scala 96:25:@31415.4]
  assign _T_414 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@31422.4 package.scala 96:25:@31423.4]
  assign _T_417 = ~ _T_414; // @[SpatialBlocks.scala 138:93:@31425.4]
  assign _T_508 = RetimeWrapper_2_io_out; // @[package.scala 96:25:@31703.4 package.scala 96:25:@31704.4]
  assign _T_514 = RetimeWrapper_3_io_out; // @[package.scala 96:25:@31711.4 package.scala 96:25:@31712.4]
  assign _T_517 = ~ _T_514; // @[SpatialBlocks.scala 138:93:@31714.4]
  assign io_in_x404_valid = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_valid; // @[sm_x425_outr_UnitPipe.scala 58:23:@31820.4]
  assign io_in_x404_bits_addr = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_bits_addr; // @[sm_x425_outr_UnitPipe.scala 58:23:@31819.4]
  assign io_in_x404_bits_size = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_bits_size; // @[sm_x425_outr_UnitPipe.scala 58:23:@31818.4]
  assign io_in_x221_TREADY = x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TREADY; // @[sm_x403_outr_UnitPipe.scala 48:23:@31516.4]
  assign io_in_x406_ready = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x406_ready; // @[sm_x425_outr_UnitPipe.scala 59:23:@31824.4]
  assign io_in_x223_outbuf_0_rPort_0_ofs_0 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@31829.4]
  assign io_in_x223_outbuf_0_rPort_0_en_0 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@31828.4]
  assign io_in_x223_outbuf_0_rPort_0_backpressure = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@31827.4]
  assign io_in_x405_valid = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_valid; // @[sm_x425_outr_UnitPipe.scala 62:23:@31833.4]
  assign io_in_x405_bits_wdata_0 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_bits_wdata_0; // @[sm_x425_outr_UnitPipe.scala 62:23:@31832.4]
  assign io_in_x405_bits_wstrb = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_bits_wstrb; // @[sm_x425_outr_UnitPipe.scala 62:23:@31831.4]
  assign io_in_x222_TVALID = x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TVALID; // @[sm_x403_outr_UnitPipe.scala 49:23:@31526.4]
  assign io_in_x222_TDATA = x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TDATA; // @[sm_x403_outr_UnitPipe.scala 49:23:@31524.4]
  assign io_sigsOut_smDoneIn_0 = x403_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@31432.4]
  assign io_sigsOut_smDoneIn_1 = x425_outr_UnitPipe_sm_io_done; // @[SpatialBlocks.scala 156:53:@31721.4]
  assign x403_outr_UnitPipe_sm_clock = clock; // @[:@31348.4]
  assign x403_outr_UnitPipe_sm_reset = reset; // @[:@31349.4]
  assign x403_outr_UnitPipe_sm_io_enable = _T_408 & _T_417; // @[SpatialBlocks.scala 140:18:@31429.4]
  assign x403_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@31431.4]
  assign x403_outr_UnitPipe_sm_io_doneIn_0 = x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@31399.4]
  assign x403_outr_UnitPipe_sm_io_doneIn_1 = x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@31400.4]
  assign x403_outr_UnitPipe_sm_io_ctrCopyDone_0 = x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@31446.4]
  assign x403_outr_UnitPipe_sm_io_ctrCopyDone_1 = x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@31447.4]
  assign RetimeWrapper_clock = clock; // @[:@31410.4]
  assign RetimeWrapper_reset = reset; // @[:@31411.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@31413.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@31412.4]
  assign RetimeWrapper_1_clock = clock; // @[:@31418.4]
  assign RetimeWrapper_1_reset = reset; // @[:@31419.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@31421.4]
  assign RetimeWrapper_1_io_in = x403_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@31420.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_clock = clock; // @[:@31449.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_reset = reset; // @[:@31450.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TVALID = io_in_x221_TVALID; // @[sm_x403_outr_UnitPipe.scala 48:23:@31517.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TDATA = io_in_x221_TDATA; // @[sm_x403_outr_UnitPipe.scala 48:23:@31515.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TID = io_in_x221_TID; // @[sm_x403_outr_UnitPipe.scala 48:23:@31511.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x221_TDEST = io_in_x221_TDEST; // @[sm_x403_outr_UnitPipe.scala 48:23:@31510.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_in_x222_TREADY = io_in_x222_TREADY; // @[sm_x403_outr_UnitPipe.scala 49:23:@31525.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x403_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x403_outr_UnitPipe.scala 92:22:@31542.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x403_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x403_outr_UnitPipe.scala 92:22:@31543.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x403_outr_UnitPipe_sm_io_childAck_0; // @[sm_x403_outr_UnitPipe.scala 92:22:@31538.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x403_outr_UnitPipe_sm_io_childAck_1; // @[sm_x403_outr_UnitPipe.scala 92:22:@31539.4]
  assign x403_outr_UnitPipe_kernelx403_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x403_outr_UnitPipe.scala 91:18:@31527.4]
  assign x425_outr_UnitPipe_sm_clock = clock; // @[:@31627.4]
  assign x425_outr_UnitPipe_sm_reset = reset; // @[:@31628.4]
  assign x425_outr_UnitPipe_sm_io_enable = _T_508 & _T_517; // @[SpatialBlocks.scala 140:18:@31718.4]
  assign x425_outr_UnitPipe_sm_io_parentAck = io_sigsIn_smChildAcks_1; // @[SpatialBlocks.scala 142:21:@31720.4]
  assign x425_outr_UnitPipe_sm_io_doneIn_0 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@31686.4]
  assign x425_outr_UnitPipe_sm_io_doneIn_1 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@31687.4]
  assign x425_outr_UnitPipe_sm_io_doneIn_2 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smDoneIn_2; // @[SpatialBlocks.scala 130:67:@31688.4]
  assign x425_outr_UnitPipe_sm_io_ctrCopyDone_0 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_0; // @[SpatialBlocks.scala 161:90:@31735.4]
  assign x425_outr_UnitPipe_sm_io_ctrCopyDone_1 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_1; // @[SpatialBlocks.scala 161:90:@31736.4]
  assign x425_outr_UnitPipe_sm_io_ctrCopyDone_2 = x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsOut_smCtrCopyDone_2; // @[SpatialBlocks.scala 161:90:@31737.4]
  assign RetimeWrapper_2_clock = clock; // @[:@31699.4]
  assign RetimeWrapper_2_reset = reset; // @[:@31700.4]
  assign RetimeWrapper_2_io_flow = 1'h1; // @[package.scala 95:18:@31702.4]
  assign RetimeWrapper_2_io_in = io_sigsIn_smEnableOuts_1; // @[package.scala 94:16:@31701.4]
  assign RetimeWrapper_3_clock = clock; // @[:@31707.4]
  assign RetimeWrapper_3_reset = reset; // @[:@31708.4]
  assign RetimeWrapper_3_io_flow = 1'h1; // @[package.scala 95:18:@31710.4]
  assign RetimeWrapper_3_io_in = x425_outr_UnitPipe_sm_io_done; // @[package.scala 94:16:@31709.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_clock = clock; // @[:@31739.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_reset = reset; // @[:@31740.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x404_ready = io_in_x404_ready; // @[sm_x425_outr_UnitPipe.scala 58:23:@31821.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x406_valid = io_in_x406_valid; // @[sm_x425_outr_UnitPipe.scala 59:23:@31823.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x219_outdram_number = io_in_x219_outdram_number; // @[sm_x425_outr_UnitPipe.scala 60:31:@31825.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x223_outbuf_0_rPort_0_output_0 = io_in_x223_outbuf_0_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@31826.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_in_x405_ready = io_in_x405_ready; // @[sm_x425_outr_UnitPipe.scala 62:23:@31834.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_0 = x425_outr_UnitPipe_sm_io_enableOut_0; // @[sm_x425_outr_UnitPipe.scala 113:22:@31857.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_1 = x425_outr_UnitPipe_sm_io_enableOut_1; // @[sm_x425_outr_UnitPipe.scala 113:22:@31858.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smEnableOuts_2 = x425_outr_UnitPipe_sm_io_enableOut_2; // @[sm_x425_outr_UnitPipe.scala 113:22:@31859.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_0 = x425_outr_UnitPipe_sm_io_childAck_0; // @[sm_x425_outr_UnitPipe.scala 113:22:@31851.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_1 = x425_outr_UnitPipe_sm_io_childAck_1; // @[sm_x425_outr_UnitPipe.scala 113:22:@31852.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_sigsIn_smChildAcks_2 = x425_outr_UnitPipe_sm_io_childAck_2; // @[sm_x425_outr_UnitPipe.scala 113:22:@31853.4]
  assign x425_outr_UnitPipe_kernelx425_outr_UnitPipe_concrete1_io_rr = io_rr; // @[sm_x425_outr_UnitPipe.scala 112:18:@31835.4]
endmodule
module RootController_kernelRootController_concrete1( // @[:@31887.2]
  input          clock, // @[:@31888.4]
  input          reset, // @[:@31889.4]
  input          io_in_x404_ready, // @[:@31890.4]
  output         io_in_x404_valid, // @[:@31890.4]
  output [63:0]  io_in_x404_bits_addr, // @[:@31890.4]
  output [31:0]  io_in_x404_bits_size, // @[:@31890.4]
  input          io_in_x221_TVALID, // @[:@31890.4]
  output         io_in_x221_TREADY, // @[:@31890.4]
  input  [255:0] io_in_x221_TDATA, // @[:@31890.4]
  input  [7:0]   io_in_x221_TID, // @[:@31890.4]
  input  [7:0]   io_in_x221_TDEST, // @[:@31890.4]
  output         io_in_x406_ready, // @[:@31890.4]
  input          io_in_x406_valid, // @[:@31890.4]
  input  [63:0]  io_in_x219_outdram_number, // @[:@31890.4]
  input          io_in_x405_ready, // @[:@31890.4]
  output         io_in_x405_valid, // @[:@31890.4]
  output [31:0]  io_in_x405_bits_wdata_0, // @[:@31890.4]
  output         io_in_x405_bits_wstrb, // @[:@31890.4]
  output         io_in_x222_TVALID, // @[:@31890.4]
  input          io_in_x222_TREADY, // @[:@31890.4]
  output [255:0] io_in_x222_TDATA, // @[:@31890.4]
  input          io_sigsIn_smEnableOuts_0, // @[:@31890.4]
  input          io_sigsIn_smChildAcks_0, // @[:@31890.4]
  output         io_sigsOut_smDoneIn_0, // @[:@31890.4]
  input          io_rr // @[:@31890.4]
);
  wire  x223_outbuf_0_clock; // @[m_x223_outbuf_0.scala 27:17:@31900.4]
  wire  x223_outbuf_0_reset; // @[m_x223_outbuf_0.scala 27:17:@31900.4]
  wire [20:0] x223_outbuf_0_io_rPort_0_ofs_0; // @[m_x223_outbuf_0.scala 27:17:@31900.4]
  wire  x223_outbuf_0_io_rPort_0_en_0; // @[m_x223_outbuf_0.scala 27:17:@31900.4]
  wire  x223_outbuf_0_io_rPort_0_backpressure; // @[m_x223_outbuf_0.scala 27:17:@31900.4]
  wire [31:0] x223_outbuf_0_io_rPort_0_output_0; // @[m_x223_outbuf_0.scala 27:17:@31900.4]
  wire  x478_sm_clock; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_reset; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_enable; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_done; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_ctrDone; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_ctrInc; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_parentAck; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_doneIn_0; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_doneIn_1; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_enableOut_0; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_enableOut_1; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_childAck_0; // @[sm_x478.scala 37:18:@31958.4]
  wire  x478_sm_io_childAck_1; // @[sm_x478.scala 37:18:@31958.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32025.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32025.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32025.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32025.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32025.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32033.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32033.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32033.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32033.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32033.4]
  wire  x478_kernelx478_concrete1_clock; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_reset; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x404_ready; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x404_valid; // @[sm_x478.scala 102:24:@32062.4]
  wire [63:0] x478_kernelx478_concrete1_io_in_x404_bits_addr; // @[sm_x478.scala 102:24:@32062.4]
  wire [31:0] x478_kernelx478_concrete1_io_in_x404_bits_size; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x221_TVALID; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x221_TREADY; // @[sm_x478.scala 102:24:@32062.4]
  wire [255:0] x478_kernelx478_concrete1_io_in_x221_TDATA; // @[sm_x478.scala 102:24:@32062.4]
  wire [7:0] x478_kernelx478_concrete1_io_in_x221_TID; // @[sm_x478.scala 102:24:@32062.4]
  wire [7:0] x478_kernelx478_concrete1_io_in_x221_TDEST; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x406_ready; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x406_valid; // @[sm_x478.scala 102:24:@32062.4]
  wire [63:0] x478_kernelx478_concrete1_io_in_x219_outdram_number; // @[sm_x478.scala 102:24:@32062.4]
  wire [20:0] x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_en_0; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure; // @[sm_x478.scala 102:24:@32062.4]
  wire [31:0] x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_output_0; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x405_ready; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x405_valid; // @[sm_x478.scala 102:24:@32062.4]
  wire [31:0] x478_kernelx478_concrete1_io_in_x405_bits_wdata_0; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x405_bits_wstrb; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x222_TVALID; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_in_x222_TREADY; // @[sm_x478.scala 102:24:@32062.4]
  wire [255:0] x478_kernelx478_concrete1_io_in_x222_TDATA; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_sigsIn_smEnableOuts_1; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_sigsIn_smChildAcks_0; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_sigsIn_smChildAcks_1; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_sigsOut_smDoneIn_0; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_sigsOut_smDoneIn_1; // @[sm_x478.scala 102:24:@32062.4]
  wire  x478_kernelx478_concrete1_io_rr; // @[sm_x478.scala 102:24:@32062.4]
  wire  _T_266; // @[package.scala 100:49:@31991.4]
  reg  _T_269; // @[package.scala 48:56:@31992.4]
  reg [31:0] _RAND_0;
  wire  _T_283; // @[package.scala 96:25:@32030.4 package.scala 96:25:@32031.4]
  wire  _T_289; // @[package.scala 96:25:@32038.4 package.scala 96:25:@32039.4]
  wire  _T_292; // @[SpatialBlocks.scala 138:93:@32041.4]
  x223_outbuf_0 x223_outbuf_0 ( // @[m_x223_outbuf_0.scala 27:17:@31900.4]
    .clock(x223_outbuf_0_clock),
    .reset(x223_outbuf_0_reset),
    .io_rPort_0_ofs_0(x223_outbuf_0_io_rPort_0_ofs_0),
    .io_rPort_0_en_0(x223_outbuf_0_io_rPort_0_en_0),
    .io_rPort_0_backpressure(x223_outbuf_0_io_rPort_0_backpressure),
    .io_rPort_0_output_0(x223_outbuf_0_io_rPort_0_output_0)
  );
  x478_sm x478_sm ( // @[sm_x478.scala 37:18:@31958.4]
    .clock(x478_sm_clock),
    .reset(x478_sm_reset),
    .io_enable(x478_sm_io_enable),
    .io_done(x478_sm_io_done),
    .io_ctrDone(x478_sm_io_ctrDone),
    .io_ctrInc(x478_sm_io_ctrInc),
    .io_parentAck(x478_sm_io_parentAck),
    .io_doneIn_0(x478_sm_io_doneIn_0),
    .io_doneIn_1(x478_sm_io_doneIn_1),
    .io_enableOut_0(x478_sm_io_enableOut_0),
    .io_enableOut_1(x478_sm_io_enableOut_1),
    .io_childAck_0(x478_sm_io_childAck_0),
    .io_childAck_1(x478_sm_io_childAck_1)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32025.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32033.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  x478_kernelx478_concrete1 x478_kernelx478_concrete1 ( // @[sm_x478.scala 102:24:@32062.4]
    .clock(x478_kernelx478_concrete1_clock),
    .reset(x478_kernelx478_concrete1_reset),
    .io_in_x404_ready(x478_kernelx478_concrete1_io_in_x404_ready),
    .io_in_x404_valid(x478_kernelx478_concrete1_io_in_x404_valid),
    .io_in_x404_bits_addr(x478_kernelx478_concrete1_io_in_x404_bits_addr),
    .io_in_x404_bits_size(x478_kernelx478_concrete1_io_in_x404_bits_size),
    .io_in_x221_TVALID(x478_kernelx478_concrete1_io_in_x221_TVALID),
    .io_in_x221_TREADY(x478_kernelx478_concrete1_io_in_x221_TREADY),
    .io_in_x221_TDATA(x478_kernelx478_concrete1_io_in_x221_TDATA),
    .io_in_x221_TID(x478_kernelx478_concrete1_io_in_x221_TID),
    .io_in_x221_TDEST(x478_kernelx478_concrete1_io_in_x221_TDEST),
    .io_in_x406_ready(x478_kernelx478_concrete1_io_in_x406_ready),
    .io_in_x406_valid(x478_kernelx478_concrete1_io_in_x406_valid),
    .io_in_x219_outdram_number(x478_kernelx478_concrete1_io_in_x219_outdram_number),
    .io_in_x223_outbuf_0_rPort_0_ofs_0(x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0),
    .io_in_x223_outbuf_0_rPort_0_en_0(x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_en_0),
    .io_in_x223_outbuf_0_rPort_0_backpressure(x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure),
    .io_in_x223_outbuf_0_rPort_0_output_0(x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_output_0),
    .io_in_x405_ready(x478_kernelx478_concrete1_io_in_x405_ready),
    .io_in_x405_valid(x478_kernelx478_concrete1_io_in_x405_valid),
    .io_in_x405_bits_wdata_0(x478_kernelx478_concrete1_io_in_x405_bits_wdata_0),
    .io_in_x405_bits_wstrb(x478_kernelx478_concrete1_io_in_x405_bits_wstrb),
    .io_in_x222_TVALID(x478_kernelx478_concrete1_io_in_x222_TVALID),
    .io_in_x222_TREADY(x478_kernelx478_concrete1_io_in_x222_TREADY),
    .io_in_x222_TDATA(x478_kernelx478_concrete1_io_in_x222_TDATA),
    .io_sigsIn_smEnableOuts_0(x478_kernelx478_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smEnableOuts_1(x478_kernelx478_concrete1_io_sigsIn_smEnableOuts_1),
    .io_sigsIn_smChildAcks_0(x478_kernelx478_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsIn_smChildAcks_1(x478_kernelx478_concrete1_io_sigsIn_smChildAcks_1),
    .io_sigsOut_smDoneIn_0(x478_kernelx478_concrete1_io_sigsOut_smDoneIn_0),
    .io_sigsOut_smDoneIn_1(x478_kernelx478_concrete1_io_sigsOut_smDoneIn_1),
    .io_rr(x478_kernelx478_concrete1_io_rr)
  );
  assign _T_266 = x478_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@31991.4]
  assign _T_283 = RetimeWrapper_io_out; // @[package.scala 96:25:@32030.4 package.scala 96:25:@32031.4]
  assign _T_289 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@32038.4 package.scala 96:25:@32039.4]
  assign _T_292 = ~ _T_289; // @[SpatialBlocks.scala 138:93:@32041.4]
  assign io_in_x404_valid = x478_kernelx478_concrete1_io_in_x404_valid; // @[sm_x478.scala 63:23:@32143.4]
  assign io_in_x404_bits_addr = x478_kernelx478_concrete1_io_in_x404_bits_addr; // @[sm_x478.scala 63:23:@32142.4]
  assign io_in_x404_bits_size = x478_kernelx478_concrete1_io_in_x404_bits_size; // @[sm_x478.scala 63:23:@32141.4]
  assign io_in_x221_TREADY = x478_kernelx478_concrete1_io_in_x221_TREADY; // @[sm_x478.scala 64:23:@32152.4]
  assign io_in_x406_ready = x478_kernelx478_concrete1_io_in_x406_ready; // @[sm_x478.scala 65:23:@32156.4]
  assign io_in_x405_valid = x478_kernelx478_concrete1_io_in_x405_valid; // @[sm_x478.scala 68:23:@32165.4]
  assign io_in_x405_bits_wdata_0 = x478_kernelx478_concrete1_io_in_x405_bits_wdata_0; // @[sm_x478.scala 68:23:@32164.4]
  assign io_in_x405_bits_wstrb = x478_kernelx478_concrete1_io_in_x405_bits_wstrb; // @[sm_x478.scala 68:23:@32163.4]
  assign io_in_x222_TVALID = x478_kernelx478_concrete1_io_in_x222_TVALID; // @[sm_x478.scala 69:23:@32175.4]
  assign io_in_x222_TDATA = x478_kernelx478_concrete1_io_in_x222_TDATA; // @[sm_x478.scala 69:23:@32173.4]
  assign io_sigsOut_smDoneIn_0 = x478_sm_io_done; // @[SpatialBlocks.scala 156:53:@32048.4]
  assign x223_outbuf_0_clock = clock; // @[:@31901.4]
  assign x223_outbuf_0_reset = reset; // @[:@31902.4]
  assign x223_outbuf_0_io_rPort_0_ofs_0 = x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_ofs_0; // @[MemInterfaceType.scala 66:44:@32161.4]
  assign x223_outbuf_0_io_rPort_0_en_0 = x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_en_0; // @[MemInterfaceType.scala 66:44:@32160.4]
  assign x223_outbuf_0_io_rPort_0_backpressure = x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_backpressure; // @[MemInterfaceType.scala 66:44:@32159.4]
  assign x478_sm_clock = clock; // @[:@31959.4]
  assign x478_sm_reset = reset; // @[:@31960.4]
  assign x478_sm_io_enable = _T_283 & _T_292; // @[SpatialBlocks.scala 140:18:@32045.4]
  assign x478_sm_io_ctrDone = x478_sm_io_ctrInc & _T_269; // @[sm_RootController.scala 82:26:@31995.4]
  assign x478_sm_io_parentAck = io_sigsIn_smChildAcks_0; // @[SpatialBlocks.scala 142:21:@32047.4]
  assign x478_sm_io_doneIn_0 = x478_kernelx478_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@32015.4]
  assign x478_sm_io_doneIn_1 = x478_kernelx478_concrete1_io_sigsOut_smDoneIn_1; // @[SpatialBlocks.scala 130:67:@32016.4]
  assign RetimeWrapper_clock = clock; // @[:@32026.4]
  assign RetimeWrapper_reset = reset; // @[:@32027.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32029.4]
  assign RetimeWrapper_io_in = io_sigsIn_smEnableOuts_0; // @[package.scala 94:16:@32028.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32034.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32035.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32037.4]
  assign RetimeWrapper_1_io_in = x478_sm_io_done; // @[package.scala 94:16:@32036.4]
  assign x478_kernelx478_concrete1_clock = clock; // @[:@32063.4]
  assign x478_kernelx478_concrete1_reset = reset; // @[:@32064.4]
  assign x478_kernelx478_concrete1_io_in_x404_ready = io_in_x404_ready; // @[sm_x478.scala 63:23:@32144.4]
  assign x478_kernelx478_concrete1_io_in_x221_TVALID = io_in_x221_TVALID; // @[sm_x478.scala 64:23:@32153.4]
  assign x478_kernelx478_concrete1_io_in_x221_TDATA = io_in_x221_TDATA; // @[sm_x478.scala 64:23:@32151.4]
  assign x478_kernelx478_concrete1_io_in_x221_TID = io_in_x221_TID; // @[sm_x478.scala 64:23:@32147.4]
  assign x478_kernelx478_concrete1_io_in_x221_TDEST = io_in_x221_TDEST; // @[sm_x478.scala 64:23:@32146.4]
  assign x478_kernelx478_concrete1_io_in_x406_valid = io_in_x406_valid; // @[sm_x478.scala 65:23:@32155.4]
  assign x478_kernelx478_concrete1_io_in_x219_outdram_number = io_in_x219_outdram_number; // @[sm_x478.scala 66:31:@32157.4]
  assign x478_kernelx478_concrete1_io_in_x223_outbuf_0_rPort_0_output_0 = x223_outbuf_0_io_rPort_0_output_0; // @[MemInterfaceType.scala 66:44:@32158.4]
  assign x478_kernelx478_concrete1_io_in_x405_ready = io_in_x405_ready; // @[sm_x478.scala 68:23:@32166.4]
  assign x478_kernelx478_concrete1_io_in_x222_TREADY = io_in_x222_TREADY; // @[sm_x478.scala 69:23:@32174.4]
  assign x478_kernelx478_concrete1_io_sigsIn_smEnableOuts_0 = x478_sm_io_enableOut_0; // @[sm_x478.scala 107:22:@32186.4]
  assign x478_kernelx478_concrete1_io_sigsIn_smEnableOuts_1 = x478_sm_io_enableOut_1; // @[sm_x478.scala 107:22:@32187.4]
  assign x478_kernelx478_concrete1_io_sigsIn_smChildAcks_0 = x478_sm_io_childAck_0; // @[sm_x478.scala 107:22:@32182.4]
  assign x478_kernelx478_concrete1_io_sigsIn_smChildAcks_1 = x478_sm_io_childAck_1; // @[sm_x478.scala 107:22:@32183.4]
  assign x478_kernelx478_concrete1_io_rr = io_rr; // @[sm_x478.scala 106:18:@32176.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_269 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_269 <= 1'h0;
    end else begin
      _T_269 <= _T_266;
    end
  end
endmodule
module AccelUnit( // @[:@32209.2]
  input          clock, // @[:@32210.4]
  input          reset, // @[:@32211.4]
  input          io_enable, // @[:@32212.4]
  output         io_done, // @[:@32212.4]
  input          io_reset, // @[:@32212.4]
  input          io_memStreams_loads_0_cmd_ready, // @[:@32212.4]
  output         io_memStreams_loads_0_cmd_valid, // @[:@32212.4]
  output [63:0]  io_memStreams_loads_0_cmd_bits_addr, // @[:@32212.4]
  output [31:0]  io_memStreams_loads_0_cmd_bits_size, // @[:@32212.4]
  output         io_memStreams_loads_0_data_ready, // @[:@32212.4]
  input          io_memStreams_loads_0_data_valid, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_0, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_1, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_2, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_3, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_4, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_5, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_6, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_7, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_8, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_9, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_10, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_11, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_12, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_13, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_14, // @[:@32212.4]
  input  [31:0]  io_memStreams_loads_0_data_bits_rdata_15, // @[:@32212.4]
  input          io_memStreams_stores_0_cmd_ready, // @[:@32212.4]
  output         io_memStreams_stores_0_cmd_valid, // @[:@32212.4]
  output [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@32212.4]
  output [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@32212.4]
  input          io_memStreams_stores_0_data_ready, // @[:@32212.4]
  output         io_memStreams_stores_0_data_valid, // @[:@32212.4]
  output [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@32212.4]
  output         io_memStreams_stores_0_data_bits_wstrb, // @[:@32212.4]
  output         io_memStreams_stores_0_wresp_ready, // @[:@32212.4]
  input          io_memStreams_stores_0_wresp_valid, // @[:@32212.4]
  input          io_memStreams_stores_0_wresp_bits, // @[:@32212.4]
  input          io_memStreams_gathers_0_cmd_ready, // @[:@32212.4]
  output         io_memStreams_gathers_0_cmd_valid, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_0, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_1, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_2, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_3, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_4, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_5, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_6, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_7, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_8, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_9, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_10, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_11, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_12, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_13, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_14, // @[:@32212.4]
  output [63:0]  io_memStreams_gathers_0_cmd_bits_addr_15, // @[:@32212.4]
  output         io_memStreams_gathers_0_data_ready, // @[:@32212.4]
  input          io_memStreams_gathers_0_data_valid, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_0, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_1, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_2, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_3, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_4, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_5, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_6, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_7, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_8, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_9, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_10, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_11, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_12, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_13, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_14, // @[:@32212.4]
  input  [31:0]  io_memStreams_gathers_0_data_bits_15, // @[:@32212.4]
  input          io_memStreams_scatters_0_cmd_ready, // @[:@32212.4]
  output         io_memStreams_scatters_0_cmd_valid, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_0, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_1, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_2, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_3, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_4, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_5, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_6, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_7, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_8, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_9, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_10, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_11, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_12, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_13, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_14, // @[:@32212.4]
  output [63:0]  io_memStreams_scatters_0_cmd_bits_addr_addr_15, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_0, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_1, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_2, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_3, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_4, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_5, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_6, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_7, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_8, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_9, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_10, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_11, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_12, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_13, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_14, // @[:@32212.4]
  output [31:0]  io_memStreams_scatters_0_cmd_bits_wdata_15, // @[:@32212.4]
  output         io_memStreams_scatters_0_wresp_ready, // @[:@32212.4]
  input          io_memStreams_scatters_0_wresp_valid, // @[:@32212.4]
  input          io_memStreams_scatters_0_wresp_bits, // @[:@32212.4]
  input          io_axiStreamsIn_0_TVALID, // @[:@32212.4]
  output         io_axiStreamsIn_0_TREADY, // @[:@32212.4]
  input  [255:0] io_axiStreamsIn_0_TDATA, // @[:@32212.4]
  input  [31:0]  io_axiStreamsIn_0_TSTRB, // @[:@32212.4]
  input  [31:0]  io_axiStreamsIn_0_TKEEP, // @[:@32212.4]
  input          io_axiStreamsIn_0_TLAST, // @[:@32212.4]
  input  [7:0]   io_axiStreamsIn_0_TID, // @[:@32212.4]
  input  [7:0]   io_axiStreamsIn_0_TDEST, // @[:@32212.4]
  input  [31:0]  io_axiStreamsIn_0_TUSER, // @[:@32212.4]
  output         io_axiStreamsOut_0_TVALID, // @[:@32212.4]
  input          io_axiStreamsOut_0_TREADY, // @[:@32212.4]
  output [255:0] io_axiStreamsOut_0_TDATA, // @[:@32212.4]
  output [31:0]  io_axiStreamsOut_0_TSTRB, // @[:@32212.4]
  output [31:0]  io_axiStreamsOut_0_TKEEP, // @[:@32212.4]
  output         io_axiStreamsOut_0_TLAST, // @[:@32212.4]
  output [7:0]   io_axiStreamsOut_0_TID, // @[:@32212.4]
  output [7:0]   io_axiStreamsOut_0_TDEST, // @[:@32212.4]
  output [31:0]  io_axiStreamsOut_0_TUSER, // @[:@32212.4]
  output         io_heap_0_req_valid, // @[:@32212.4]
  output         io_heap_0_req_bits_allocDealloc, // @[:@32212.4]
  output [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@32212.4]
  input          io_heap_0_resp_valid, // @[:@32212.4]
  input          io_heap_0_resp_bits_allocDealloc, // @[:@32212.4]
  input  [63:0]  io_heap_0_resp_bits_sizeAddr, // @[:@32212.4]
  input  [63:0]  io_argIns_0, // @[:@32212.4]
  input  [63:0]  io_argIns_1, // @[:@32212.4]
  input          io_argOuts_0_port_ready, // @[:@32212.4]
  output         io_argOuts_0_port_valid, // @[:@32212.4]
  output [63:0]  io_argOuts_0_port_bits, // @[:@32212.4]
  input  [63:0]  io_argOuts_0_echo // @[:@32212.4]
);
  wire  SingleCounter_clock; // @[Main.scala 40:32:@32360.4]
  wire  SingleCounter_reset; // @[Main.scala 40:32:@32360.4]
  wire  SingleCounter_io_input_reset; // @[Main.scala 40:32:@32360.4]
  wire  SingleCounter_io_output_done; // @[Main.scala 40:32:@32360.4]
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@32378.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@32378.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@32378.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@32378.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@32378.4]
  wire  SRFF_clock; // @[Main.scala 44:28:@32387.4]
  wire  SRFF_reset; // @[Main.scala 44:28:@32387.4]
  wire  SRFF_io_input_set; // @[Main.scala 44:28:@32387.4]
  wire  SRFF_io_input_reset; // @[Main.scala 44:28:@32387.4]
  wire  SRFF_io_input_asyn_reset; // @[Main.scala 44:28:@32387.4]
  wire  SRFF_io_output; // @[Main.scala 44:28:@32387.4]
  wire  RootController_sm_clock; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_reset; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_enable; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_done; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_rst; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_ctrDone; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_ctrInc; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_parentAck; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_doneIn_0; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_enableOut_0; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RootController_sm_io_childAck_0; // @[sm_RootController.scala 36:18:@32426.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@32458.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@32458.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@32458.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@32458.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@32458.4]
  wire  RootController_kernelRootController_concrete1_clock; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_reset; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x404_ready; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x404_valid; // @[sm_RootController.scala 91:24:@32520.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x404_bits_addr; // @[sm_RootController.scala 91:24:@32520.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x404_bits_size; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x221_TVALID; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x221_TREADY; // @[sm_RootController.scala 91:24:@32520.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x221_TDATA; // @[sm_RootController.scala 91:24:@32520.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x221_TID; // @[sm_RootController.scala 91:24:@32520.4]
  wire [7:0] RootController_kernelRootController_concrete1_io_in_x221_TDEST; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x406_ready; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x406_valid; // @[sm_RootController.scala 91:24:@32520.4]
  wire [63:0] RootController_kernelRootController_concrete1_io_in_x219_outdram_number; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x405_ready; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x405_valid; // @[sm_RootController.scala 91:24:@32520.4]
  wire [31:0] RootController_kernelRootController_concrete1_io_in_x405_bits_wdata_0; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x405_bits_wstrb; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x222_TVALID; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_in_x222_TREADY; // @[sm_RootController.scala 91:24:@32520.4]
  wire [255:0] RootController_kernelRootController_concrete1_io_in_x222_TDATA; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[sm_RootController.scala 91:24:@32520.4]
  wire  RootController_kernelRootController_concrete1_io_rr; // @[sm_RootController.scala 91:24:@32520.4]
  wire  _T_599; // @[package.scala 96:25:@32383.4 package.scala 96:25:@32384.4]
  wire  _T_664; // @[Main.scala 46:50:@32454.4]
  wire  _T_665; // @[Main.scala 46:59:@32455.4]
  wire  _T_677; // @[package.scala 100:49:@32475.4]
  reg  _T_680; // @[package.scala 48:56:@32476.4]
  reg [31:0] _RAND_0;
  SingleCounter SingleCounter ( // @[Main.scala 40:32:@32360.4]
    .clock(SingleCounter_clock),
    .reset(SingleCounter_reset),
    .io_input_reset(SingleCounter_io_input_reset),
    .io_output_done(SingleCounter_io_output_done)
  );
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@32378.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  SRFF SRFF ( // @[Main.scala 44:28:@32387.4]
    .clock(SRFF_clock),
    .reset(SRFF_reset),
    .io_input_set(SRFF_io_input_set),
    .io_input_reset(SRFF_io_input_reset),
    .io_input_asyn_reset(SRFF_io_input_asyn_reset),
    .io_output(SRFF_io_output)
  );
  RootController_sm RootController_sm ( // @[sm_RootController.scala 36:18:@32426.4]
    .clock(RootController_sm_clock),
    .reset(RootController_sm_reset),
    .io_enable(RootController_sm_io_enable),
    .io_done(RootController_sm_io_done),
    .io_rst(RootController_sm_io_rst),
    .io_ctrDone(RootController_sm_io_ctrDone),
    .io_ctrInc(RootController_sm_io_ctrInc),
    .io_parentAck(RootController_sm_io_parentAck),
    .io_doneIn_0(RootController_sm_io_doneIn_0),
    .io_enableOut_0(RootController_sm_io_enableOut_0),
    .io_childAck_0(RootController_sm_io_childAck_0)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@32458.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  RootController_kernelRootController_concrete1 RootController_kernelRootController_concrete1 ( // @[sm_RootController.scala 91:24:@32520.4]
    .clock(RootController_kernelRootController_concrete1_clock),
    .reset(RootController_kernelRootController_concrete1_reset),
    .io_in_x404_ready(RootController_kernelRootController_concrete1_io_in_x404_ready),
    .io_in_x404_valid(RootController_kernelRootController_concrete1_io_in_x404_valid),
    .io_in_x404_bits_addr(RootController_kernelRootController_concrete1_io_in_x404_bits_addr),
    .io_in_x404_bits_size(RootController_kernelRootController_concrete1_io_in_x404_bits_size),
    .io_in_x221_TVALID(RootController_kernelRootController_concrete1_io_in_x221_TVALID),
    .io_in_x221_TREADY(RootController_kernelRootController_concrete1_io_in_x221_TREADY),
    .io_in_x221_TDATA(RootController_kernelRootController_concrete1_io_in_x221_TDATA),
    .io_in_x221_TID(RootController_kernelRootController_concrete1_io_in_x221_TID),
    .io_in_x221_TDEST(RootController_kernelRootController_concrete1_io_in_x221_TDEST),
    .io_in_x406_ready(RootController_kernelRootController_concrete1_io_in_x406_ready),
    .io_in_x406_valid(RootController_kernelRootController_concrete1_io_in_x406_valid),
    .io_in_x219_outdram_number(RootController_kernelRootController_concrete1_io_in_x219_outdram_number),
    .io_in_x405_ready(RootController_kernelRootController_concrete1_io_in_x405_ready),
    .io_in_x405_valid(RootController_kernelRootController_concrete1_io_in_x405_valid),
    .io_in_x405_bits_wdata_0(RootController_kernelRootController_concrete1_io_in_x405_bits_wdata_0),
    .io_in_x405_bits_wstrb(RootController_kernelRootController_concrete1_io_in_x405_bits_wstrb),
    .io_in_x222_TVALID(RootController_kernelRootController_concrete1_io_in_x222_TVALID),
    .io_in_x222_TREADY(RootController_kernelRootController_concrete1_io_in_x222_TREADY),
    .io_in_x222_TDATA(RootController_kernelRootController_concrete1_io_in_x222_TDATA),
    .io_sigsIn_smEnableOuts_0(RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0),
    .io_sigsIn_smChildAcks_0(RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0),
    .io_sigsOut_smDoneIn_0(RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0),
    .io_rr(RootController_kernelRootController_concrete1_io_rr)
  );
  assign _T_599 = RetimeWrapper_io_out; // @[package.scala 96:25:@32383.4 package.scala 96:25:@32384.4]
  assign _T_664 = io_enable & _T_599; // @[Main.scala 46:50:@32454.4]
  assign _T_665 = ~ SRFF_io_output; // @[Main.scala 46:59:@32455.4]
  assign _T_677 = RootController_sm_io_ctrInc == 1'h0; // @[package.scala 100:49:@32475.4]
  assign io_done = SRFF_io_output; // @[Main.scala 53:23:@32474.4]
  assign io_memStreams_loads_0_cmd_valid = 1'h0;
  assign io_memStreams_loads_0_cmd_bits_addr = 64'h0;
  assign io_memStreams_loads_0_cmd_bits_size = 32'h0;
  assign io_memStreams_loads_0_data_ready = 1'h0;
  assign io_memStreams_stores_0_cmd_valid = RootController_kernelRootController_concrete1_io_in_x404_valid; // @[sm_RootController.scala 60:23:@32583.4]
  assign io_memStreams_stores_0_cmd_bits_addr = RootController_kernelRootController_concrete1_io_in_x404_bits_addr; // @[sm_RootController.scala 60:23:@32582.4]
  assign io_memStreams_stores_0_cmd_bits_size = RootController_kernelRootController_concrete1_io_in_x404_bits_size; // @[sm_RootController.scala 60:23:@32581.4]
  assign io_memStreams_stores_0_data_valid = RootController_kernelRootController_concrete1_io_in_x405_valid; // @[sm_RootController.scala 64:23:@32600.4]
  assign io_memStreams_stores_0_data_bits_wdata_0 = RootController_kernelRootController_concrete1_io_in_x405_bits_wdata_0; // @[sm_RootController.scala 64:23:@32599.4]
  assign io_memStreams_stores_0_data_bits_wstrb = RootController_kernelRootController_concrete1_io_in_x405_bits_wstrb; // @[sm_RootController.scala 64:23:@32598.4]
  assign io_memStreams_stores_0_wresp_ready = RootController_kernelRootController_concrete1_io_in_x406_ready; // @[sm_RootController.scala 62:23:@32596.4]
  assign io_memStreams_gathers_0_cmd_valid = 1'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_0 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_1 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_2 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_3 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_4 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_5 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_6 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_7 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_8 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_9 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_10 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_11 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_12 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_13 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_14 = 64'h0;
  assign io_memStreams_gathers_0_cmd_bits_addr_15 = 64'h0;
  assign io_memStreams_gathers_0_data_ready = 1'h0;
  assign io_memStreams_scatters_0_cmd_valid = 1'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_0 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_1 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_2 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_3 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_4 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_5 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_6 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_7 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_8 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_9 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_10 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_11 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_12 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_13 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_14 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_addr_addr_15 = 64'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_0 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_1 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_2 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_3 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_4 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_5 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_6 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_7 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_8 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_9 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_10 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_11 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_12 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_13 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_14 = 32'h0;
  assign io_memStreams_scatters_0_cmd_bits_wdata_15 = 32'h0;
  assign io_memStreams_scatters_0_wresp_ready = 1'h0;
  assign io_axiStreamsIn_0_TREADY = RootController_kernelRootController_concrete1_io_in_x221_TREADY; // @[sm_RootController.scala 61:23:@32592.4]
  assign io_axiStreamsOut_0_TVALID = RootController_kernelRootController_concrete1_io_in_x222_TVALID; // @[sm_RootController.scala 65:23:@32610.4]
  assign io_axiStreamsOut_0_TDATA = RootController_kernelRootController_concrete1_io_in_x222_TDATA; // @[sm_RootController.scala 65:23:@32608.4]
  assign io_axiStreamsOut_0_TSTRB = 32'hffffffff; // @[sm_RootController.scala 65:23:@32607.4]
  assign io_axiStreamsOut_0_TKEEP = 32'hffffffff; // @[sm_RootController.scala 65:23:@32606.4]
  assign io_axiStreamsOut_0_TLAST = 1'h0; // @[sm_RootController.scala 65:23:@32605.4]
  assign io_axiStreamsOut_0_TID = 8'h0; // @[sm_RootController.scala 65:23:@32604.4]
  assign io_axiStreamsOut_0_TDEST = 8'h0; // @[sm_RootController.scala 65:23:@32603.4]
  assign io_axiStreamsOut_0_TUSER = 32'h4; // @[sm_RootController.scala 65:23:@32602.4]
  assign io_heap_0_req_valid = 1'h0;
  assign io_heap_0_req_bits_allocDealloc = 1'h0;
  assign io_heap_0_req_bits_sizeAddr = 64'h0;
  assign io_argOuts_0_port_valid = 1'h0;
  assign io_argOuts_0_port_bits = 64'h0;
  assign SingleCounter_clock = clock; // @[:@32361.4]
  assign SingleCounter_reset = reset; // @[:@32362.4]
  assign SingleCounter_io_input_reset = reset; // @[Main.scala 41:79:@32376.4]
  assign RetimeWrapper_clock = clock; // @[:@32379.4]
  assign RetimeWrapper_reset = reset; // @[:@32380.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@32382.4]
  assign RetimeWrapper_io_in = SingleCounter_io_output_done; // @[package.scala 94:16:@32381.4]
  assign SRFF_clock = clock; // @[:@32388.4]
  assign SRFF_reset = reset; // @[:@32389.4]
  assign SRFF_io_input_set = RootController_sm_io_done; // @[Main.scala 62:29:@32638.4]
  assign SRFF_io_input_reset = RetimeWrapper_1_io_out; // @[Main.scala 51:31:@32472.4]
  assign SRFF_io_input_asyn_reset = RetimeWrapper_1_io_out; // @[Main.scala 52:36:@32473.4]
  assign RootController_sm_clock = clock; // @[:@32427.4]
  assign RootController_sm_reset = reset; // @[:@32428.4]
  assign RootController_sm_io_enable = _T_664 & _T_665; // @[Main.scala 50:33:@32471.4 SpatialBlocks.scala 140:18:@32505.4]
  assign RootController_sm_io_rst = RetimeWrapper_1_io_out; // @[SpatialBlocks.scala 134:15:@32499.4]
  assign RootController_sm_io_ctrDone = RootController_sm_io_ctrInc & _T_680; // @[Main.scala 54:34:@32479.4]
  assign RootController_sm_io_parentAck = 1'h0; // @[Main.scala 49:36:@32467.4 SpatialBlocks.scala 142:21:@32507.4]
  assign RootController_sm_io_doneIn_0 = RootController_kernelRootController_concrete1_io_sigsOut_smDoneIn_0; // @[SpatialBlocks.scala 130:67:@32496.4]
  assign RetimeWrapper_1_clock = clock; // @[:@32459.4]
  assign RetimeWrapper_1_reset = reset; // @[:@32460.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@32462.4]
  assign RetimeWrapper_1_io_in = reset | io_reset; // @[package.scala 94:16:@32461.4]
  assign RootController_kernelRootController_concrete1_clock = clock; // @[:@32521.4]
  assign RootController_kernelRootController_concrete1_reset = reset; // @[:@32522.4]
  assign RootController_kernelRootController_concrete1_io_in_x404_ready = io_memStreams_stores_0_cmd_ready; // @[sm_RootController.scala 60:23:@32584.4]
  assign RootController_kernelRootController_concrete1_io_in_x221_TVALID = io_axiStreamsIn_0_TVALID; // @[sm_RootController.scala 61:23:@32593.4]
  assign RootController_kernelRootController_concrete1_io_in_x221_TDATA = io_axiStreamsIn_0_TDATA; // @[sm_RootController.scala 61:23:@32591.4]
  assign RootController_kernelRootController_concrete1_io_in_x221_TID = io_axiStreamsIn_0_TID; // @[sm_RootController.scala 61:23:@32587.4]
  assign RootController_kernelRootController_concrete1_io_in_x221_TDEST = io_axiStreamsIn_0_TDEST; // @[sm_RootController.scala 61:23:@32586.4]
  assign RootController_kernelRootController_concrete1_io_in_x406_valid = io_memStreams_stores_0_wresp_valid; // @[sm_RootController.scala 62:23:@32595.4]
  assign RootController_kernelRootController_concrete1_io_in_x219_outdram_number = io_argIns_1; // @[sm_RootController.scala 63:31:@32597.4]
  assign RootController_kernelRootController_concrete1_io_in_x405_ready = io_memStreams_stores_0_data_ready; // @[sm_RootController.scala 64:23:@32601.4]
  assign RootController_kernelRootController_concrete1_io_in_x222_TREADY = io_axiStreamsOut_0_TREADY; // @[sm_RootController.scala 65:23:@32609.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smEnableOuts_0 = RootController_sm_io_enableOut_0; // @[sm_RootController.scala 96:22:@32619.4]
  assign RootController_kernelRootController_concrete1_io_sigsIn_smChildAcks_0 = RootController_sm_io_childAck_0; // @[sm_RootController.scala 96:22:@32617.4]
  assign RootController_kernelRootController_concrete1_io_rr = RetimeWrapper_io_out; // @[sm_RootController.scala 95:18:@32611.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_680 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_680 <= 1'h0;
    end else begin
      _T_680 <= _T_677;
    end
  end
endmodule
module Counter( // @[:@32640.2]
  input        clock, // @[:@32641.4]
  input        reset, // @[:@32642.4]
  input        io_enable, // @[:@32643.4]
  output [5:0] io_out, // @[:@32643.4]
  output [5:0] io_next // @[:@32643.4]
);
  reg [5:0] count; // @[Counter.scala 15:22:@32645.4]
  reg [31:0] _RAND_0;
  wire [6:0] _T_17; // @[Counter.scala 17:24:@32646.4]
  wire [5:0] newCount; // @[Counter.scala 17:24:@32647.4]
  wire [5:0] _GEN_0; // @[Counter.scala 21:26:@32652.6]
  assign _T_17 = count + 6'h1; // @[Counter.scala 17:24:@32646.4]
  assign newCount = count + 6'h1; // @[Counter.scala 17:24:@32647.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@32652.6]
  assign io_out = count; // @[Counter.scala 25:10:@32655.4]
  assign io_next = count + 6'h1; // @[Counter.scala 26:11:@32656.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 6'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module SRAM_17( // @[:@32692.2]
  input         clock, // @[:@32693.4]
  input         reset, // @[:@32694.4]
  input  [5:0]  io_raddr, // @[:@32695.4]
  input         io_wen, // @[:@32695.4]
  input  [5:0]  io_waddr, // @[:@32695.4]
  input  [63:0] io_wdata_addr, // @[:@32695.4]
  input  [31:0] io_wdata_size, // @[:@32695.4]
  output [63:0] io_rdata_addr, // @[:@32695.4]
  output [31:0] io_rdata_size // @[:@32695.4]
);
  wire [95:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@32697.4]
  wire [95:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@32697.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@32697.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@32697.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@32697.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@32697.4]
  wire [5:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@32697.4]
  wire [5:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@32697.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@32697.4]
  wire [95:0] _T_17; // @[SRAM.scala 175:38:@32711.4]
  wire  _T_20; // @[SRAM.scala 182:49:@32716.4]
  wire  _T_21; // @[SRAM.scala 182:37:@32717.4]
  reg  _T_24; // @[SRAM.scala 182:29:@32718.4]
  reg [31:0] _RAND_0;
  reg [95:0] _T_28; // @[SRAM.scala 183:29:@32721.4]
  reg [95:0] _RAND_1;
  wire [95:0] _T_29; // @[SRAM.scala 184:22:@32723.4]
  SRAMVerilogAWS #(.DWIDTH(96), .WORDS(64), .AWIDTH(6)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@32697.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_17 = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:38:@32711.4]
  assign _T_20 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@32716.4]
  assign _T_21 = io_wen & _T_20; // @[SRAM.scala 182:37:@32717.4]
  assign _T_29 = _T_24 ? _T_28 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:22:@32723.4]
  assign io_rdata_addr = _T_29[95:32]; // @[SRAM.scala 184:16:@32732.4]
  assign io_rdata_size = _T_29[31:0]; // @[SRAM.scala 184:16:@32731.4]
  assign SRAMVerilogAWS_wdata = {io_wdata_addr,io_wdata_size}; // @[SRAM.scala 175:20:@32712.4]
  assign SRAMVerilogAWS_backpressure = 1'h1; // @[SRAM.scala 176:27:@32713.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@32709.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@32715.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@32714.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@32710.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@32708.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@32707.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_24 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  _T_28 = _RAND_1[95:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_24 <= 1'h0;
    end else begin
      _T_24 <= _T_21;
    end
    if (reset) begin
      _T_28 <= 96'h0;
    end else begin
      _T_28 <= _T_17;
    end
  end
endmodule
module FIFO( // @[:@32734.2]
  input         clock, // @[:@32735.4]
  input         reset, // @[:@32736.4]
  output        io_in_ready, // @[:@32737.4]
  input         io_in_valid, // @[:@32737.4]
  input  [63:0] io_in_bits_addr, // @[:@32737.4]
  input  [31:0] io_in_bits_size, // @[:@32737.4]
  input         io_out_ready, // @[:@32737.4]
  output        io_out_valid, // @[:@32737.4]
  output [63:0] io_out_bits_addr, // @[:@32737.4]
  output [31:0] io_out_bits_size // @[:@32737.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@33133.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@33133.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@33133.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@33133.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@33133.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@33143.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@33143.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@33143.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@33143.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@33143.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@33158.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@33158.4]
  wire [5:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@33158.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@33158.4]
  wire [5:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@33158.4]
  wire [63:0] SRAM_io_wdata_addr; // @[FIFO.scala 73:19:@33158.4]
  wire [31:0] SRAM_io_wdata_size; // @[FIFO.scala 73:19:@33158.4]
  wire [63:0] SRAM_io_rdata_addr; // @[FIFO.scala 73:19:@33158.4]
  wire [31:0] SRAM_io_rdata_size; // @[FIFO.scala 73:19:@33158.4]
  wire  writeEn; // @[FIFO.scala 30:29:@33131.4]
  wire  readEn; // @[FIFO.scala 31:29:@33132.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@33153.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@33154.4]
  wire  _T_824; // @[FIFO.scala 45:27:@33155.4]
  wire  empty; // @[FIFO.scala 45:24:@33156.4]
  wire  full; // @[FIFO.scala 46:23:@33157.4]
  wire  _T_827; // @[FIFO.scala 83:17:@33170.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@33171.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@33133.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@33143.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_17 SRAM ( // @[FIFO.scala 73:19:@33158.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata_addr(SRAM_io_wdata_addr),
    .io_wdata_size(SRAM_io_wdata_size),
    .io_rdata_addr(SRAM_io_rdata_addr),
    .io_rdata_size(SRAM_io_rdata_size)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@33131.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@33132.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@33154.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@33155.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@33156.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@33157.4]
  assign _T_827 = writeEn != readEn; // @[FIFO.scala 83:17:@33170.4]
  assign _GEN_0 = _T_827 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@33171.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@33177.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@33175.4]
  assign io_out_bits_addr = SRAM_io_rdata_addr; // @[FIFO.scala 79:17:@33168.4]
  assign io_out_bits_size = SRAM_io_rdata_size; // @[FIFO.scala 79:17:@33167.4]
  assign enqCounter_clock = clock; // @[:@33134.4]
  assign enqCounter_reset = reset; // @[:@33135.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@33141.4]
  assign deqCounter_clock = clock; // @[:@33144.4]
  assign deqCounter_reset = reset; // @[:@33145.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@33151.4]
  assign SRAM_clock = clock; // @[:@33159.4]
  assign SRAM_reset = reset; // @[:@33160.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@33162.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@33163.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@33164.4]
  assign SRAM_io_wdata_addr = io_in_bits_addr; // @[FIFO.scala 78:16:@33166.4]
  assign SRAM_io_wdata_size = io_in_bits_size; // @[FIFO.scala 78:16:@33165.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_827) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module Counter_2( // @[:@33179.2]
  input        clock, // @[:@33180.4]
  input        reset, // @[:@33181.4]
  input        io_enable, // @[:@33182.4]
  output [3:0] io_out // @[:@33182.4]
);
  reg [3:0] count; // @[Counter.scala 15:22:@33184.4]
  reg [31:0] _RAND_0;
  wire [4:0] _T_17; // @[Counter.scala 17:24:@33185.4]
  wire [3:0] newCount; // @[Counter.scala 17:24:@33186.4]
  wire [3:0] _GEN_0; // @[Counter.scala 21:26:@33191.6]
  assign _T_17 = count + 4'h1; // @[Counter.scala 17:24:@33185.4]
  assign newCount = count + 4'h1; // @[Counter.scala 17:24:@33186.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@33191.6]
  assign io_out = count; // @[Counter.scala 25:10:@33194.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_enable) begin
        count <= newCount;
      end
    end
  end
endmodule
module Counter_4( // @[:@33215.2]
  input        clock, // @[:@33216.4]
  input        reset, // @[:@33217.4]
  input        io_reset, // @[:@33218.4]
  input        io_enable, // @[:@33218.4]
  input  [1:0] io_stride, // @[:@33218.4]
  output [1:0] io_out, // @[:@33218.4]
  output [1:0] io_next // @[:@33218.4]
);
  reg [1:0] count; // @[Counter.scala 15:22:@33220.4]
  reg [31:0] _RAND_0;
  wire [2:0] _T_17; // @[Counter.scala 17:24:@33221.4]
  wire [1:0] newCount; // @[Counter.scala 17:24:@33222.4]
  wire [1:0] _GEN_0; // @[Counter.scala 21:26:@33227.6]
  wire [1:0] _GEN_1; // @[Counter.scala 19:18:@33223.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@33221.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@33222.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@33227.6]
  assign _GEN_1 = io_reset ? 2'h0 : _GEN_0; // @[Counter.scala 19:18:@33223.4]
  assign io_out = count; // @[Counter.scala 25:10:@33230.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@33231.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 2'h0;
    end else begin
      if (io_reset) begin
        count <= 2'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module SRAM_18( // @[:@33267.2]
  input         clock, // @[:@33268.4]
  input         reset, // @[:@33269.4]
  input  [1:0]  io_raddr, // @[:@33270.4]
  input         io_wen, // @[:@33270.4]
  input  [1:0]  io_waddr, // @[:@33270.4]
  input  [31:0] io_wdata, // @[:@33270.4]
  output [31:0] io_rdata, // @[:@33270.4]
  input         io_backpressure // @[:@33270.4]
);
  wire [31:0] SRAMVerilogAWS_rdata; // @[SRAM.scala 169:30:@33272.4]
  wire [31:0] SRAMVerilogAWS_wdata; // @[SRAM.scala 169:30:@33272.4]
  wire  SRAMVerilogAWS_backpressure; // @[SRAM.scala 169:30:@33272.4]
  wire  SRAMVerilogAWS_wen; // @[SRAM.scala 169:30:@33272.4]
  wire  SRAMVerilogAWS_waddrEn; // @[SRAM.scala 169:30:@33272.4]
  wire  SRAMVerilogAWS_raddrEn; // @[SRAM.scala 169:30:@33272.4]
  wire [1:0] SRAMVerilogAWS_waddr; // @[SRAM.scala 169:30:@33272.4]
  wire [1:0] SRAMVerilogAWS_raddr; // @[SRAM.scala 169:30:@33272.4]
  wire  SRAMVerilogAWS_clk; // @[SRAM.scala 169:30:@33272.4]
  wire  _T_19; // @[SRAM.scala 182:49:@33290.4]
  wire  _T_20; // @[SRAM.scala 182:37:@33291.4]
  reg  _T_23; // @[SRAM.scala 182:29:@33292.4]
  reg [31:0] _RAND_0;
  reg [31:0] _T_26; // @[SRAM.scala 183:29:@33294.4]
  reg [31:0] _RAND_1;
  SRAMVerilogAWS #(.DWIDTH(32), .WORDS(4), .AWIDTH(2)) SRAMVerilogAWS ( // @[SRAM.scala 169:30:@33272.4]
    .rdata(SRAMVerilogAWS_rdata),
    .wdata(SRAMVerilogAWS_wdata),
    .backpressure(SRAMVerilogAWS_backpressure),
    .wen(SRAMVerilogAWS_wen),
    .waddrEn(SRAMVerilogAWS_waddrEn),
    .raddrEn(SRAMVerilogAWS_raddrEn),
    .waddr(SRAMVerilogAWS_waddr),
    .raddr(SRAMVerilogAWS_raddr),
    .clk(SRAMVerilogAWS_clk)
  );
  assign _T_19 = io_raddr == io_waddr; // @[SRAM.scala 182:49:@33290.4]
  assign _T_20 = io_wen & _T_19; // @[SRAM.scala 182:37:@33291.4]
  assign io_rdata = _T_23 ? _T_26 : SRAMVerilogAWS_rdata; // @[SRAM.scala 184:16:@33299.4]
  assign SRAMVerilogAWS_wdata = io_wdata; // @[SRAM.scala 175:20:@33286.4]
  assign SRAMVerilogAWS_backpressure = io_backpressure; // @[SRAM.scala 176:27:@33287.4]
  assign SRAMVerilogAWS_wen = io_wen; // @[SRAM.scala 173:18:@33284.4]
  assign SRAMVerilogAWS_waddrEn = 1'h1; // @[SRAM.scala 178:22:@33289.4]
  assign SRAMVerilogAWS_raddrEn = 1'h1; // @[SRAM.scala 177:22:@33288.4]
  assign SRAMVerilogAWS_waddr = io_waddr; // @[SRAM.scala 174:20:@33285.4]
  assign SRAMVerilogAWS_raddr = io_raddr; // @[SRAM.scala 172:20:@33283.4]
  assign SRAMVerilogAWS_clk = clock; // @[SRAM.scala 171:18:@33282.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_23 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_26 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _T_20;
    end
    if (reset) begin
      _T_26 <= 32'h0;
    end else begin
      _T_26 <= io_wdata;
    end
  end
endmodule
module FIFO_1( // @[:@33301.2]
  input         clock, // @[:@33302.4]
  input         reset, // @[:@33303.4]
  output        io_in_ready, // @[:@33304.4]
  input         io_in_valid, // @[:@33304.4]
  input  [31:0] io_in_bits, // @[:@33304.4]
  input         io_out_ready, // @[:@33304.4]
  output        io_out_valid, // @[:@33304.4]
  output [31:0] io_out_bits // @[:@33304.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@33330.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@33330.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@33330.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@33330.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@33330.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@33330.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@33330.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@33340.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@33340.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@33340.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@33340.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@33340.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@33340.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@33340.4]
  wire  SRAM_clock; // @[FIFO.scala 73:19:@33355.4]
  wire  SRAM_reset; // @[FIFO.scala 73:19:@33355.4]
  wire [1:0] SRAM_io_raddr; // @[FIFO.scala 73:19:@33355.4]
  wire  SRAM_io_wen; // @[FIFO.scala 73:19:@33355.4]
  wire [1:0] SRAM_io_waddr; // @[FIFO.scala 73:19:@33355.4]
  wire [31:0] SRAM_io_wdata; // @[FIFO.scala 73:19:@33355.4]
  wire [31:0] SRAM_io_rdata; // @[FIFO.scala 73:19:@33355.4]
  wire  SRAM_io_backpressure; // @[FIFO.scala 73:19:@33355.4]
  wire  writeEn; // @[FIFO.scala 30:29:@33328.4]
  wire  readEn; // @[FIFO.scala 31:29:@33329.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@33350.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@33351.4]
  wire  _T_104; // @[FIFO.scala 45:27:@33352.4]
  wire  empty; // @[FIFO.scala 45:24:@33353.4]
  wire  full; // @[FIFO.scala 46:23:@33354.4]
  wire  _T_107; // @[FIFO.scala 83:17:@33365.4]
  wire  _GEN_0; // @[FIFO.scala 83:29:@33366.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@33330.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@33340.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  SRAM_18 SRAM ( // @[FIFO.scala 73:19:@33355.4]
    .clock(SRAM_clock),
    .reset(SRAM_reset),
    .io_raddr(SRAM_io_raddr),
    .io_wen(SRAM_io_wen),
    .io_waddr(SRAM_io_waddr),
    .io_wdata(SRAM_io_wdata),
    .io_rdata(SRAM_io_rdata),
    .io_backpressure(SRAM_io_backpressure)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@33328.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@33329.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@33351.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@33352.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@33353.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@33354.4]
  assign _T_107 = writeEn != readEn; // @[FIFO.scala 83:17:@33365.4]
  assign _GEN_0 = _T_107 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@33366.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@33372.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@33370.4]
  assign io_out_bits = SRAM_io_rdata; // @[FIFO.scala 79:17:@33363.4]
  assign enqCounter_clock = clock; // @[:@33331.4]
  assign enqCounter_reset = reset; // @[:@33332.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@33338.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@33339.4]
  assign deqCounter_clock = clock; // @[:@33341.4]
  assign deqCounter_reset = reset; // @[:@33342.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@33348.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@33349.4]
  assign SRAM_clock = clock; // @[:@33356.4]
  assign SRAM_reset = reset; // @[:@33357.4]
  assign SRAM_io_raddr = readEn ? deqCounter_io_next : deqCounter_io_out; // @[FIFO.scala 75:16:@33359.4]
  assign SRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 76:14:@33360.4]
  assign SRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 77:16:@33361.4]
  assign SRAM_io_wdata = io_in_bits; // @[FIFO.scala 78:16:@33362.4]
  assign SRAM_io_backpressure = 1'h1; // @[FIFO.scala 80:23:@33364.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_107) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec( // @[:@35759.2]
  input         clock, // @[:@35760.4]
  input         reset, // @[:@35761.4]
  output        io_in_ready, // @[:@35762.4]
  input         io_in_valid, // @[:@35762.4]
  input  [31:0] io_in_bits_0, // @[:@35762.4]
  input         io_out_ready, // @[:@35762.4]
  output        io_out_valid, // @[:@35762.4]
  output [31:0] io_out_bits_0, // @[:@35762.4]
  output [31:0] io_out_bits_1, // @[:@35762.4]
  output [31:0] io_out_bits_2, // @[:@35762.4]
  output [31:0] io_out_bits_3, // @[:@35762.4]
  output [31:0] io_out_bits_4, // @[:@35762.4]
  output [31:0] io_out_bits_5, // @[:@35762.4]
  output [31:0] io_out_bits_6, // @[:@35762.4]
  output [31:0] io_out_bits_7, // @[:@35762.4]
  output [31:0] io_out_bits_8, // @[:@35762.4]
  output [31:0] io_out_bits_9, // @[:@35762.4]
  output [31:0] io_out_bits_10, // @[:@35762.4]
  output [31:0] io_out_bits_11, // @[:@35762.4]
  output [31:0] io_out_bits_12, // @[:@35762.4]
  output [31:0] io_out_bits_13, // @[:@35762.4]
  output [31:0] io_out_bits_14, // @[:@35762.4]
  output [31:0] io_out_bits_15 // @[:@35762.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@35766.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@35766.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@35766.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@35766.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@35777.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@35777.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@35777.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@35777.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@35790.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@35790.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@35790.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@35790.4]
  wire [31:0] fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@35790.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@35790.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@35790.4]
  wire [31:0] fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@35790.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@35825.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@35825.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@35825.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@35825.4]
  wire [31:0] fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@35825.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@35825.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@35825.4]
  wire [31:0] fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@35825.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@35860.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@35860.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@35860.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@35860.4]
  wire [31:0] fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@35860.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@35860.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@35860.4]
  wire [31:0] fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@35860.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@35895.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@35895.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@35895.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@35895.4]
  wire [31:0] fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@35895.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@35895.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@35895.4]
  wire [31:0] fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@35895.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@35930.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@35930.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@35930.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@35930.4]
  wire [31:0] fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@35930.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@35930.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@35930.4]
  wire [31:0] fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@35930.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@35965.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@35965.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@35965.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@35965.4]
  wire [31:0] fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@35965.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@35965.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@35965.4]
  wire [31:0] fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@35965.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@36000.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@36000.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@36000.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@36000.4]
  wire [31:0] fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@36000.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@36000.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@36000.4]
  wire [31:0] fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@36000.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@36035.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@36035.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@36035.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@36035.4]
  wire [31:0] fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@36035.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@36035.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@36035.4]
  wire [31:0] fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@36035.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@36070.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@36070.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@36070.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@36070.4]
  wire [31:0] fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@36070.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@36070.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@36070.4]
  wire [31:0] fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@36070.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@36105.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@36105.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@36105.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@36105.4]
  wire [31:0] fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@36105.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@36105.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@36105.4]
  wire [31:0] fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@36105.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@36140.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@36140.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@36140.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@36140.4]
  wire [31:0] fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@36140.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@36140.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@36140.4]
  wire [31:0] fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@36140.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@36175.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@36175.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@36175.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@36175.4]
  wire [31:0] fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@36175.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@36175.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@36175.4]
  wire [31:0] fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@36175.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@36210.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@36210.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@36210.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@36210.4]
  wire [31:0] fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@36210.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@36210.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@36210.4]
  wire [31:0] fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@36210.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@36245.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@36245.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@36245.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@36245.4]
  wire [31:0] fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@36245.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@36245.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@36245.4]
  wire [31:0] fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@36245.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@36280.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@36280.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@36280.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@36280.4]
  wire [31:0] fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@36280.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@36280.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@36280.4]
  wire [31:0] fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@36280.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@36315.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@36315.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@36315.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@36315.4]
  wire [31:0] fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@36315.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@36315.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@36315.4]
  wire [31:0] fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@36315.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@35765.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@35788.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@35815.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@35850.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@35885.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@35920.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@35955.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@35990.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@36025.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@36060.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@36095.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@36130.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@36165.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@36200.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@36235.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@36270.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@36305.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@36340.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36351.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36352.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36353.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36354.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36355.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36356.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36357.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36358.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36359.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36360.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36361.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36362.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36363.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36364.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36365.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@36382.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36366.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@36401.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@36402.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@36403.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@36404.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@36405.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@36406.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@36407.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@36408.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@36409.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@36410.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@36411.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@36412.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@36413.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@36414.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@35766.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@35777.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_1 fifos_0 ( // @[FIFOVec.scala 40:19:@35790.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_1 fifos_1 ( // @[FIFOVec.scala 40:19:@35825.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_1 fifos_2 ( // @[FIFOVec.scala 40:19:@35860.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_1 fifos_3 ( // @[FIFOVec.scala 40:19:@35895.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_1 fifos_4 ( // @[FIFOVec.scala 40:19:@35930.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_1 fifos_5 ( // @[FIFOVec.scala 40:19:@35965.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_1 fifos_6 ( // @[FIFOVec.scala 40:19:@36000.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_1 fifos_7 ( // @[FIFOVec.scala 40:19:@36035.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_1 fifos_8 ( // @[FIFOVec.scala 40:19:@36070.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_1 fifos_9 ( // @[FIFOVec.scala 40:19:@36105.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_1 fifos_10 ( // @[FIFOVec.scala 40:19:@36140.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_1 fifos_11 ( // @[FIFOVec.scala 40:19:@36175.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_1 fifos_12 ( // @[FIFOVec.scala 40:19:@36210.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_1 fifos_13 ( // @[FIFOVec.scala 40:19:@36245.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_1 fifos_14 ( // @[FIFOVec.scala 40:19:@36280.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_1 fifos_15 ( // @[FIFOVec.scala 40:19:@36315.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@35765.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@35788.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@35815.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@35850.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@35885.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@35920.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@35955.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@35990.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@36025.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@36060.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@36095.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@36130.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@36165.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@36200.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@36235.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@36270.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@36305.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@36340.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36351.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36352.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36353.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36354.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36355.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36356.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36357.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36358.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36359.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36360.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36361.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36362.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36363.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36364.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36365.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@36382.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@36350.4 FIFOVec.scala 49:42:@36366.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@36401.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@36402.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@36403.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@36404.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@36405.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@36406.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@36407.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@36408.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@36409.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@36410.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@36411.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@36412.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@36413.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@36414.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@36383.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@36417.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@36725.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@36726.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@36727.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@36728.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@36729.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@36730.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@36731.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@36732.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@36733.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@36734.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@36735.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@36736.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@36737.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@36738.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@36739.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@36740.4]
  assign enqCounter_clock = clock; // @[:@35767.4]
  assign enqCounter_reset = reset; // @[:@35768.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@35775.4]
  assign deqCounter_clock = clock; // @[:@35778.4]
  assign deqCounter_reset = reset; // @[:@35779.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@35786.4]
  assign fifos_0_clock = clock; // @[:@35791.4]
  assign fifos_0_reset = reset; // @[:@35792.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@35818.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@35820.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@35824.4]
  assign fifos_1_clock = clock; // @[:@35826.4]
  assign fifos_1_reset = reset; // @[:@35827.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@35853.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@35855.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@35859.4]
  assign fifos_2_clock = clock; // @[:@35861.4]
  assign fifos_2_reset = reset; // @[:@35862.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@35888.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@35890.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@35894.4]
  assign fifos_3_clock = clock; // @[:@35896.4]
  assign fifos_3_reset = reset; // @[:@35897.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@35923.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@35925.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@35929.4]
  assign fifos_4_clock = clock; // @[:@35931.4]
  assign fifos_4_reset = reset; // @[:@35932.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@35958.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@35960.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@35964.4]
  assign fifos_5_clock = clock; // @[:@35966.4]
  assign fifos_5_reset = reset; // @[:@35967.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@35993.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@35995.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@35999.4]
  assign fifos_6_clock = clock; // @[:@36001.4]
  assign fifos_6_reset = reset; // @[:@36002.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@36028.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36030.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36034.4]
  assign fifos_7_clock = clock; // @[:@36036.4]
  assign fifos_7_reset = reset; // @[:@36037.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@36063.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36065.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36069.4]
  assign fifos_8_clock = clock; // @[:@36071.4]
  assign fifos_8_reset = reset; // @[:@36072.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@36098.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36100.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36104.4]
  assign fifos_9_clock = clock; // @[:@36106.4]
  assign fifos_9_reset = reset; // @[:@36107.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@36133.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36135.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36139.4]
  assign fifos_10_clock = clock; // @[:@36141.4]
  assign fifos_10_reset = reset; // @[:@36142.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@36168.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36170.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36174.4]
  assign fifos_11_clock = clock; // @[:@36176.4]
  assign fifos_11_reset = reset; // @[:@36177.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@36203.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36205.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36209.4]
  assign fifos_12_clock = clock; // @[:@36211.4]
  assign fifos_12_reset = reset; // @[:@36212.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@36238.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36240.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36244.4]
  assign fifos_13_clock = clock; // @[:@36246.4]
  assign fifos_13_reset = reset; // @[:@36247.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@36273.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36275.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36279.4]
  assign fifos_14_clock = clock; // @[:@36281.4]
  assign fifos_14_reset = reset; // @[:@36282.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@36308.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36310.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36314.4]
  assign fifos_15_clock = clock; // @[:@36316.4]
  assign fifos_15_reset = reset; // @[:@36317.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@36343.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@36345.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@36349.4]
endmodule
module FFRAM( // @[:@36814.2]
  input        clock, // @[:@36815.4]
  input        reset, // @[:@36816.4]
  input  [1:0] io_raddr, // @[:@36817.4]
  input        io_wen, // @[:@36817.4]
  input  [1:0] io_waddr, // @[:@36817.4]
  input        io_wdata, // @[:@36817.4]
  output       io_rdata, // @[:@36817.4]
  input        io_banks_0_wdata_valid, // @[:@36817.4]
  input        io_banks_0_wdata_bits, // @[:@36817.4]
  input        io_banks_1_wdata_valid, // @[:@36817.4]
  input        io_banks_1_wdata_bits, // @[:@36817.4]
  input        io_banks_2_wdata_valid, // @[:@36817.4]
  input        io_banks_2_wdata_bits, // @[:@36817.4]
  input        io_banks_3_wdata_valid, // @[:@36817.4]
  input        io_banks_3_wdata_bits // @[:@36817.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@36821.4]
  reg [31:0] _RAND_0;
  wire  _T_88; // @[SRAM.scala 148:37:@36822.4]
  wire  _T_89; // @[SRAM.scala 148:25:@36823.4]
  wire  _T_90; // @[SRAM.scala 148:15:@36824.4]
  wire  _T_91; // @[SRAM.scala 149:15:@36826.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@36825.4]
  reg  regs_1; // @[SRAM.scala 145:20:@36832.4]
  reg [31:0] _RAND_1;
  wire  _T_97; // @[SRAM.scala 148:37:@36833.4]
  wire  _T_98; // @[SRAM.scala 148:25:@36834.4]
  wire  _T_99; // @[SRAM.scala 148:15:@36835.4]
  wire  _T_100; // @[SRAM.scala 149:15:@36837.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@36836.4]
  reg  regs_2; // @[SRAM.scala 145:20:@36843.4]
  reg [31:0] _RAND_2;
  wire  _T_106; // @[SRAM.scala 148:37:@36844.4]
  wire  _T_107; // @[SRAM.scala 148:25:@36845.4]
  wire  _T_108; // @[SRAM.scala 148:15:@36846.4]
  wire  _T_109; // @[SRAM.scala 149:15:@36848.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@36847.4]
  reg  regs_3; // @[SRAM.scala 145:20:@36854.4]
  reg [31:0] _RAND_3;
  wire  _T_115; // @[SRAM.scala 148:37:@36855.4]
  wire  _T_116; // @[SRAM.scala 148:25:@36856.4]
  wire  _T_117; // @[SRAM.scala 148:15:@36857.4]
  wire  _T_118; // @[SRAM.scala 149:15:@36859.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@36858.4]
  wire  _GEN_5; // @[SRAM.scala 155:12:@36868.4]
  wire  _GEN_6; // @[SRAM.scala 155:12:@36868.4]
  assign _T_88 = io_waddr == 2'h0; // @[SRAM.scala 148:37:@36822.4]
  assign _T_89 = io_wen & _T_88; // @[SRAM.scala 148:25:@36823.4]
  assign _T_90 = io_banks_0_wdata_valid | _T_89; // @[SRAM.scala 148:15:@36824.4]
  assign _T_91 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@36826.6]
  assign _GEN_0 = _T_90 ? _T_91 : regs_0; // @[SRAM.scala 148:48:@36825.4]
  assign _T_97 = io_waddr == 2'h1; // @[SRAM.scala 148:37:@36833.4]
  assign _T_98 = io_wen & _T_97; // @[SRAM.scala 148:25:@36834.4]
  assign _T_99 = io_banks_1_wdata_valid | _T_98; // @[SRAM.scala 148:15:@36835.4]
  assign _T_100 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@36837.6]
  assign _GEN_1 = _T_99 ? _T_100 : regs_1; // @[SRAM.scala 148:48:@36836.4]
  assign _T_106 = io_waddr == 2'h2; // @[SRAM.scala 148:37:@36844.4]
  assign _T_107 = io_wen & _T_106; // @[SRAM.scala 148:25:@36845.4]
  assign _T_108 = io_banks_2_wdata_valid | _T_107; // @[SRAM.scala 148:15:@36846.4]
  assign _T_109 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@36848.6]
  assign _GEN_2 = _T_108 ? _T_109 : regs_2; // @[SRAM.scala 148:48:@36847.4]
  assign _T_115 = io_waddr == 2'h3; // @[SRAM.scala 148:37:@36855.4]
  assign _T_116 = io_wen & _T_115; // @[SRAM.scala 148:25:@36856.4]
  assign _T_117 = io_banks_3_wdata_valid | _T_116; // @[SRAM.scala 148:15:@36857.4]
  assign _T_118 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@36859.6]
  assign _GEN_3 = _T_117 ? _T_118 : regs_3; // @[SRAM.scala 148:48:@36858.4]
  assign _GEN_5 = 2'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@36868.4]
  assign _GEN_6 = 2'h2 == io_raddr ? regs_2 : _GEN_5; // @[SRAM.scala 155:12:@36868.4]
  assign io_rdata = 2'h3 == io_raddr ? regs_3 : _GEN_6; // @[SRAM.scala 155:12:@36868.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_90) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_99) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_108) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_117) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_17( // @[:@36870.2]
  input   clock, // @[:@36871.4]
  input   reset, // @[:@36872.4]
  output  io_in_ready, // @[:@36873.4]
  input   io_in_valid, // @[:@36873.4]
  input   io_in_bits, // @[:@36873.4]
  input   io_out_ready, // @[:@36873.4]
  output  io_out_valid, // @[:@36873.4]
  output  io_out_bits // @[:@36873.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@36899.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@36899.4]
  wire  enqCounter_io_reset; // @[FIFO.scala 34:26:@36899.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@36899.4]
  wire [1:0] enqCounter_io_stride; // @[FIFO.scala 34:26:@36899.4]
  wire [1:0] enqCounter_io_out; // @[FIFO.scala 34:26:@36899.4]
  wire [1:0] enqCounter_io_next; // @[FIFO.scala 34:26:@36899.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@36909.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@36909.4]
  wire  deqCounter_io_reset; // @[FIFO.scala 38:26:@36909.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@36909.4]
  wire [1:0] deqCounter_io_stride; // @[FIFO.scala 38:26:@36909.4]
  wire [1:0] deqCounter_io_out; // @[FIFO.scala 38:26:@36909.4]
  wire [1:0] deqCounter_io_next; // @[FIFO.scala 38:26:@36909.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@36924.4]
  wire [1:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@36924.4]
  wire [1:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@36924.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@36924.4]
  wire  writeEn; // @[FIFO.scala 30:29:@36897.4]
  wire  readEn; // @[FIFO.scala 31:29:@36898.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@36919.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@36920.4]
  wire  _T_104; // @[FIFO.scala 45:27:@36921.4]
  wire  empty; // @[FIFO.scala 45:24:@36922.4]
  wire  full; // @[FIFO.scala 46:23:@36923.4]
  wire  _T_157; // @[FIFO.scala 83:17:@37010.4]
  wire  _GEN_4; // @[FIFO.scala 83:29:@37011.4]
  Counter_4 enqCounter ( // @[FIFO.scala 34:26:@36899.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_reset(enqCounter_io_reset),
    .io_enable(enqCounter_io_enable),
    .io_stride(enqCounter_io_stride),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter_4 deqCounter ( // @[FIFO.scala 38:26:@36909.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_reset(deqCounter_io_reset),
    .io_enable(deqCounter_io_enable),
    .io_stride(deqCounter_io_stride),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM FFRAM ( // @[FIFO.scala 49:19:@36924.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@36897.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@36898.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@36920.4]
  assign _T_104 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@36921.4]
  assign empty = ptrMatch & _T_104; // @[FIFO.scala 45:24:@36922.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@36923.4]
  assign _T_157 = writeEn != readEn; // @[FIFO.scala 83:17:@37010.4]
  assign _GEN_4 = _T_157 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@37011.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@37017.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@37015.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@36949.4]
  assign enqCounter_clock = clock; // @[:@36900.4]
  assign enqCounter_reset = reset; // @[:@36901.4]
  assign enqCounter_io_reset = 1'h0;
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@36907.4]
  assign enqCounter_io_stride = 2'h1; // @[FIFO.scala 37:24:@36908.4]
  assign deqCounter_clock = clock; // @[:@36910.4]
  assign deqCounter_reset = reset; // @[:@36911.4]
  assign deqCounter_io_reset = 1'h0;
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@36917.4]
  assign deqCounter_io_stride = 2'h1; // @[FIFO.scala 41:24:@36918.4]
  assign FFRAM_clock = clock; // @[:@36925.4]
  assign FFRAM_reset = reset; // @[:@36926.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@36945.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@36946.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@36947.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@36948.4]
  assign FFRAM_io_banks_0_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@36951.4]
  assign FFRAM_io_banks_0_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@36950.4]
  assign FFRAM_io_banks_1_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@36954.4]
  assign FFRAM_io_banks_1_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@36953.4]
  assign FFRAM_io_banks_2_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@36957.4]
  assign FFRAM_io_banks_2_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@36956.4]
  assign FFRAM_io_banks_3_wdata_valid = 1'h0; // @[FIFO.scala 59:15:@36960.4]
  assign FFRAM_io_banks_3_wdata_bits = 1'h0; // @[FIFO.scala 59:15:@36959.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_157) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module FIFOVec_1( // @[:@40634.2]
  input   clock, // @[:@40635.4]
  input   reset, // @[:@40636.4]
  output  io_in_ready, // @[:@40637.4]
  input   io_in_valid, // @[:@40637.4]
  input   io_in_bits_0, // @[:@40637.4]
  input   io_out_ready, // @[:@40637.4]
  output  io_out_valid, // @[:@40637.4]
  output  io_out_bits_0, // @[:@40637.4]
  output  io_out_bits_1, // @[:@40637.4]
  output  io_out_bits_2, // @[:@40637.4]
  output  io_out_bits_3, // @[:@40637.4]
  output  io_out_bits_4, // @[:@40637.4]
  output  io_out_bits_5, // @[:@40637.4]
  output  io_out_bits_6, // @[:@40637.4]
  output  io_out_bits_7, // @[:@40637.4]
  output  io_out_bits_8, // @[:@40637.4]
  output  io_out_bits_9, // @[:@40637.4]
  output  io_out_bits_10, // @[:@40637.4]
  output  io_out_bits_11, // @[:@40637.4]
  output  io_out_bits_12, // @[:@40637.4]
  output  io_out_bits_13, // @[:@40637.4]
  output  io_out_bits_14, // @[:@40637.4]
  output  io_out_bits_15 // @[:@40637.4]
);
  wire  enqCounter_clock; // @[FIFOVec.scala 24:26:@40641.4]
  wire  enqCounter_reset; // @[FIFOVec.scala 24:26:@40641.4]
  wire  enqCounter_io_enable; // @[FIFOVec.scala 24:26:@40641.4]
  wire [3:0] enqCounter_io_out; // @[FIFOVec.scala 24:26:@40641.4]
  wire  deqCounter_clock; // @[FIFOVec.scala 28:26:@40652.4]
  wire  deqCounter_reset; // @[FIFOVec.scala 28:26:@40652.4]
  wire  deqCounter_io_enable; // @[FIFOVec.scala 28:26:@40652.4]
  wire [3:0] deqCounter_io_out; // @[FIFOVec.scala 28:26:@40652.4]
  wire  fifos_0_clock; // @[FIFOVec.scala 40:19:@40665.4]
  wire  fifos_0_reset; // @[FIFOVec.scala 40:19:@40665.4]
  wire  fifos_0_io_in_ready; // @[FIFOVec.scala 40:19:@40665.4]
  wire  fifos_0_io_in_valid; // @[FIFOVec.scala 40:19:@40665.4]
  wire  fifos_0_io_in_bits; // @[FIFOVec.scala 40:19:@40665.4]
  wire  fifos_0_io_out_ready; // @[FIFOVec.scala 40:19:@40665.4]
  wire  fifos_0_io_out_valid; // @[FIFOVec.scala 40:19:@40665.4]
  wire  fifos_0_io_out_bits; // @[FIFOVec.scala 40:19:@40665.4]
  wire  fifos_1_clock; // @[FIFOVec.scala 40:19:@40700.4]
  wire  fifos_1_reset; // @[FIFOVec.scala 40:19:@40700.4]
  wire  fifos_1_io_in_ready; // @[FIFOVec.scala 40:19:@40700.4]
  wire  fifos_1_io_in_valid; // @[FIFOVec.scala 40:19:@40700.4]
  wire  fifos_1_io_in_bits; // @[FIFOVec.scala 40:19:@40700.4]
  wire  fifos_1_io_out_ready; // @[FIFOVec.scala 40:19:@40700.4]
  wire  fifos_1_io_out_valid; // @[FIFOVec.scala 40:19:@40700.4]
  wire  fifos_1_io_out_bits; // @[FIFOVec.scala 40:19:@40700.4]
  wire  fifos_2_clock; // @[FIFOVec.scala 40:19:@40735.4]
  wire  fifos_2_reset; // @[FIFOVec.scala 40:19:@40735.4]
  wire  fifos_2_io_in_ready; // @[FIFOVec.scala 40:19:@40735.4]
  wire  fifos_2_io_in_valid; // @[FIFOVec.scala 40:19:@40735.4]
  wire  fifos_2_io_in_bits; // @[FIFOVec.scala 40:19:@40735.4]
  wire  fifos_2_io_out_ready; // @[FIFOVec.scala 40:19:@40735.4]
  wire  fifos_2_io_out_valid; // @[FIFOVec.scala 40:19:@40735.4]
  wire  fifos_2_io_out_bits; // @[FIFOVec.scala 40:19:@40735.4]
  wire  fifos_3_clock; // @[FIFOVec.scala 40:19:@40770.4]
  wire  fifos_3_reset; // @[FIFOVec.scala 40:19:@40770.4]
  wire  fifos_3_io_in_ready; // @[FIFOVec.scala 40:19:@40770.4]
  wire  fifos_3_io_in_valid; // @[FIFOVec.scala 40:19:@40770.4]
  wire  fifos_3_io_in_bits; // @[FIFOVec.scala 40:19:@40770.4]
  wire  fifos_3_io_out_ready; // @[FIFOVec.scala 40:19:@40770.4]
  wire  fifos_3_io_out_valid; // @[FIFOVec.scala 40:19:@40770.4]
  wire  fifos_3_io_out_bits; // @[FIFOVec.scala 40:19:@40770.4]
  wire  fifos_4_clock; // @[FIFOVec.scala 40:19:@40805.4]
  wire  fifos_4_reset; // @[FIFOVec.scala 40:19:@40805.4]
  wire  fifos_4_io_in_ready; // @[FIFOVec.scala 40:19:@40805.4]
  wire  fifos_4_io_in_valid; // @[FIFOVec.scala 40:19:@40805.4]
  wire  fifos_4_io_in_bits; // @[FIFOVec.scala 40:19:@40805.4]
  wire  fifos_4_io_out_ready; // @[FIFOVec.scala 40:19:@40805.4]
  wire  fifos_4_io_out_valid; // @[FIFOVec.scala 40:19:@40805.4]
  wire  fifos_4_io_out_bits; // @[FIFOVec.scala 40:19:@40805.4]
  wire  fifos_5_clock; // @[FIFOVec.scala 40:19:@40840.4]
  wire  fifos_5_reset; // @[FIFOVec.scala 40:19:@40840.4]
  wire  fifos_5_io_in_ready; // @[FIFOVec.scala 40:19:@40840.4]
  wire  fifos_5_io_in_valid; // @[FIFOVec.scala 40:19:@40840.4]
  wire  fifos_5_io_in_bits; // @[FIFOVec.scala 40:19:@40840.4]
  wire  fifos_5_io_out_ready; // @[FIFOVec.scala 40:19:@40840.4]
  wire  fifos_5_io_out_valid; // @[FIFOVec.scala 40:19:@40840.4]
  wire  fifos_5_io_out_bits; // @[FIFOVec.scala 40:19:@40840.4]
  wire  fifos_6_clock; // @[FIFOVec.scala 40:19:@40875.4]
  wire  fifos_6_reset; // @[FIFOVec.scala 40:19:@40875.4]
  wire  fifos_6_io_in_ready; // @[FIFOVec.scala 40:19:@40875.4]
  wire  fifos_6_io_in_valid; // @[FIFOVec.scala 40:19:@40875.4]
  wire  fifos_6_io_in_bits; // @[FIFOVec.scala 40:19:@40875.4]
  wire  fifos_6_io_out_ready; // @[FIFOVec.scala 40:19:@40875.4]
  wire  fifos_6_io_out_valid; // @[FIFOVec.scala 40:19:@40875.4]
  wire  fifos_6_io_out_bits; // @[FIFOVec.scala 40:19:@40875.4]
  wire  fifos_7_clock; // @[FIFOVec.scala 40:19:@40910.4]
  wire  fifos_7_reset; // @[FIFOVec.scala 40:19:@40910.4]
  wire  fifos_7_io_in_ready; // @[FIFOVec.scala 40:19:@40910.4]
  wire  fifos_7_io_in_valid; // @[FIFOVec.scala 40:19:@40910.4]
  wire  fifos_7_io_in_bits; // @[FIFOVec.scala 40:19:@40910.4]
  wire  fifos_7_io_out_ready; // @[FIFOVec.scala 40:19:@40910.4]
  wire  fifos_7_io_out_valid; // @[FIFOVec.scala 40:19:@40910.4]
  wire  fifos_7_io_out_bits; // @[FIFOVec.scala 40:19:@40910.4]
  wire  fifos_8_clock; // @[FIFOVec.scala 40:19:@40945.4]
  wire  fifos_8_reset; // @[FIFOVec.scala 40:19:@40945.4]
  wire  fifos_8_io_in_ready; // @[FIFOVec.scala 40:19:@40945.4]
  wire  fifos_8_io_in_valid; // @[FIFOVec.scala 40:19:@40945.4]
  wire  fifos_8_io_in_bits; // @[FIFOVec.scala 40:19:@40945.4]
  wire  fifos_8_io_out_ready; // @[FIFOVec.scala 40:19:@40945.4]
  wire  fifos_8_io_out_valid; // @[FIFOVec.scala 40:19:@40945.4]
  wire  fifos_8_io_out_bits; // @[FIFOVec.scala 40:19:@40945.4]
  wire  fifos_9_clock; // @[FIFOVec.scala 40:19:@40980.4]
  wire  fifos_9_reset; // @[FIFOVec.scala 40:19:@40980.4]
  wire  fifos_9_io_in_ready; // @[FIFOVec.scala 40:19:@40980.4]
  wire  fifos_9_io_in_valid; // @[FIFOVec.scala 40:19:@40980.4]
  wire  fifos_9_io_in_bits; // @[FIFOVec.scala 40:19:@40980.4]
  wire  fifos_9_io_out_ready; // @[FIFOVec.scala 40:19:@40980.4]
  wire  fifos_9_io_out_valid; // @[FIFOVec.scala 40:19:@40980.4]
  wire  fifos_9_io_out_bits; // @[FIFOVec.scala 40:19:@40980.4]
  wire  fifos_10_clock; // @[FIFOVec.scala 40:19:@41015.4]
  wire  fifos_10_reset; // @[FIFOVec.scala 40:19:@41015.4]
  wire  fifos_10_io_in_ready; // @[FIFOVec.scala 40:19:@41015.4]
  wire  fifos_10_io_in_valid; // @[FIFOVec.scala 40:19:@41015.4]
  wire  fifos_10_io_in_bits; // @[FIFOVec.scala 40:19:@41015.4]
  wire  fifos_10_io_out_ready; // @[FIFOVec.scala 40:19:@41015.4]
  wire  fifos_10_io_out_valid; // @[FIFOVec.scala 40:19:@41015.4]
  wire  fifos_10_io_out_bits; // @[FIFOVec.scala 40:19:@41015.4]
  wire  fifos_11_clock; // @[FIFOVec.scala 40:19:@41050.4]
  wire  fifos_11_reset; // @[FIFOVec.scala 40:19:@41050.4]
  wire  fifos_11_io_in_ready; // @[FIFOVec.scala 40:19:@41050.4]
  wire  fifos_11_io_in_valid; // @[FIFOVec.scala 40:19:@41050.4]
  wire  fifos_11_io_in_bits; // @[FIFOVec.scala 40:19:@41050.4]
  wire  fifos_11_io_out_ready; // @[FIFOVec.scala 40:19:@41050.4]
  wire  fifos_11_io_out_valid; // @[FIFOVec.scala 40:19:@41050.4]
  wire  fifos_11_io_out_bits; // @[FIFOVec.scala 40:19:@41050.4]
  wire  fifos_12_clock; // @[FIFOVec.scala 40:19:@41085.4]
  wire  fifos_12_reset; // @[FIFOVec.scala 40:19:@41085.4]
  wire  fifos_12_io_in_ready; // @[FIFOVec.scala 40:19:@41085.4]
  wire  fifos_12_io_in_valid; // @[FIFOVec.scala 40:19:@41085.4]
  wire  fifos_12_io_in_bits; // @[FIFOVec.scala 40:19:@41085.4]
  wire  fifos_12_io_out_ready; // @[FIFOVec.scala 40:19:@41085.4]
  wire  fifos_12_io_out_valid; // @[FIFOVec.scala 40:19:@41085.4]
  wire  fifos_12_io_out_bits; // @[FIFOVec.scala 40:19:@41085.4]
  wire  fifos_13_clock; // @[FIFOVec.scala 40:19:@41120.4]
  wire  fifos_13_reset; // @[FIFOVec.scala 40:19:@41120.4]
  wire  fifos_13_io_in_ready; // @[FIFOVec.scala 40:19:@41120.4]
  wire  fifos_13_io_in_valid; // @[FIFOVec.scala 40:19:@41120.4]
  wire  fifos_13_io_in_bits; // @[FIFOVec.scala 40:19:@41120.4]
  wire  fifos_13_io_out_ready; // @[FIFOVec.scala 40:19:@41120.4]
  wire  fifos_13_io_out_valid; // @[FIFOVec.scala 40:19:@41120.4]
  wire  fifos_13_io_out_bits; // @[FIFOVec.scala 40:19:@41120.4]
  wire  fifos_14_clock; // @[FIFOVec.scala 40:19:@41155.4]
  wire  fifos_14_reset; // @[FIFOVec.scala 40:19:@41155.4]
  wire  fifos_14_io_in_ready; // @[FIFOVec.scala 40:19:@41155.4]
  wire  fifos_14_io_in_valid; // @[FIFOVec.scala 40:19:@41155.4]
  wire  fifos_14_io_in_bits; // @[FIFOVec.scala 40:19:@41155.4]
  wire  fifos_14_io_out_ready; // @[FIFOVec.scala 40:19:@41155.4]
  wire  fifos_14_io_out_valid; // @[FIFOVec.scala 40:19:@41155.4]
  wire  fifos_14_io_out_bits; // @[FIFOVec.scala 40:19:@41155.4]
  wire  fifos_15_clock; // @[FIFOVec.scala 40:19:@41190.4]
  wire  fifos_15_reset; // @[FIFOVec.scala 40:19:@41190.4]
  wire  fifos_15_io_in_ready; // @[FIFOVec.scala 40:19:@41190.4]
  wire  fifos_15_io_in_valid; // @[FIFOVec.scala 40:19:@41190.4]
  wire  fifos_15_io_in_bits; // @[FIFOVec.scala 40:19:@41190.4]
  wire  fifos_15_io_out_ready; // @[FIFOVec.scala 40:19:@41190.4]
  wire  fifos_15_io_out_valid; // @[FIFOVec.scala 40:19:@41190.4]
  wire  fifos_15_io_out_bits; // @[FIFOVec.scala 40:19:@41190.4]
  wire  writeEn; // @[FIFOVec.scala 21:29:@40640.4]
  wire [15:0] enqDecoder; // @[OneHot.scala 45:35:@40663.4]
  wire  _T_149; // @[FIFOVec.scala 42:49:@40690.4]
  wire  _T_158; // @[FIFOVec.scala 42:49:@40725.4]
  wire  _T_167; // @[FIFOVec.scala 42:49:@40760.4]
  wire  _T_176; // @[FIFOVec.scala 42:49:@40795.4]
  wire  _T_185; // @[FIFOVec.scala 42:49:@40830.4]
  wire  _T_194; // @[FIFOVec.scala 42:49:@40865.4]
  wire  _T_203; // @[FIFOVec.scala 42:49:@40900.4]
  wire  _T_212; // @[FIFOVec.scala 42:49:@40935.4]
  wire  _T_221; // @[FIFOVec.scala 42:49:@40970.4]
  wire  _T_230; // @[FIFOVec.scala 42:49:@41005.4]
  wire  _T_239; // @[FIFOVec.scala 42:49:@41040.4]
  wire  _T_248; // @[FIFOVec.scala 42:49:@41075.4]
  wire  _T_257; // @[FIFOVec.scala 42:49:@41110.4]
  wire  _T_266; // @[FIFOVec.scala 42:49:@41145.4]
  wire  _T_275; // @[FIFOVec.scala 42:49:@41180.4]
  wire  _T_284; // @[FIFOVec.scala 42:49:@41215.4]
  wire  _T_296_0; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41226.4]
  wire  _T_296_1; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41227.4]
  wire  _GEN_1; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_2; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41228.4]
  wire  _GEN_2; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_3; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41229.4]
  wire  _GEN_3; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_4; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41230.4]
  wire  _GEN_4; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_5; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41231.4]
  wire  _GEN_5; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_6; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41232.4]
  wire  _GEN_6; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_7; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41233.4]
  wire  _GEN_7; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_8; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41234.4]
  wire  _GEN_8; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_9; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41235.4]
  wire  _GEN_9; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_10; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41236.4]
  wire  _GEN_10; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_11; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41237.4]
  wire  _GEN_11; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_12; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41238.4]
  wire  _GEN_12; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_13; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41239.4]
  wire  _GEN_13; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_14; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41240.4]
  wire  _GEN_14; // @[FIFOVec.scala 49:21:@41257.4]
  wire  _T_296_15; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41241.4]
  wire  _T_355; // @[FIFOVec.scala 51:93:@41276.4]
  wire  _T_356; // @[FIFOVec.scala 51:93:@41277.4]
  wire  _T_357; // @[FIFOVec.scala 51:93:@41278.4]
  wire  _T_358; // @[FIFOVec.scala 51:93:@41279.4]
  wire  _T_359; // @[FIFOVec.scala 51:93:@41280.4]
  wire  _T_360; // @[FIFOVec.scala 51:93:@41281.4]
  wire  _T_361; // @[FIFOVec.scala 51:93:@41282.4]
  wire  _T_362; // @[FIFOVec.scala 51:93:@41283.4]
  wire  _T_363; // @[FIFOVec.scala 51:93:@41284.4]
  wire  _T_364; // @[FIFOVec.scala 51:93:@41285.4]
  wire  _T_365; // @[FIFOVec.scala 51:93:@41286.4]
  wire  _T_366; // @[FIFOVec.scala 51:93:@41287.4]
  wire  _T_367; // @[FIFOVec.scala 51:93:@41288.4]
  wire  _T_368; // @[FIFOVec.scala 51:93:@41289.4]
  Counter_2 enqCounter ( // @[FIFOVec.scala 24:26:@40641.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out)
  );
  Counter_2 deqCounter ( // @[FIFOVec.scala 28:26:@40652.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out)
  );
  FIFO_17 fifos_0 ( // @[FIFOVec.scala 40:19:@40665.4]
    .clock(fifos_0_clock),
    .reset(fifos_0_reset),
    .io_in_ready(fifos_0_io_in_ready),
    .io_in_valid(fifos_0_io_in_valid),
    .io_in_bits(fifos_0_io_in_bits),
    .io_out_ready(fifos_0_io_out_ready),
    .io_out_valid(fifos_0_io_out_valid),
    .io_out_bits(fifos_0_io_out_bits)
  );
  FIFO_17 fifos_1 ( // @[FIFOVec.scala 40:19:@40700.4]
    .clock(fifos_1_clock),
    .reset(fifos_1_reset),
    .io_in_ready(fifos_1_io_in_ready),
    .io_in_valid(fifos_1_io_in_valid),
    .io_in_bits(fifos_1_io_in_bits),
    .io_out_ready(fifos_1_io_out_ready),
    .io_out_valid(fifos_1_io_out_valid),
    .io_out_bits(fifos_1_io_out_bits)
  );
  FIFO_17 fifos_2 ( // @[FIFOVec.scala 40:19:@40735.4]
    .clock(fifos_2_clock),
    .reset(fifos_2_reset),
    .io_in_ready(fifos_2_io_in_ready),
    .io_in_valid(fifos_2_io_in_valid),
    .io_in_bits(fifos_2_io_in_bits),
    .io_out_ready(fifos_2_io_out_ready),
    .io_out_valid(fifos_2_io_out_valid),
    .io_out_bits(fifos_2_io_out_bits)
  );
  FIFO_17 fifos_3 ( // @[FIFOVec.scala 40:19:@40770.4]
    .clock(fifos_3_clock),
    .reset(fifos_3_reset),
    .io_in_ready(fifos_3_io_in_ready),
    .io_in_valid(fifos_3_io_in_valid),
    .io_in_bits(fifos_3_io_in_bits),
    .io_out_ready(fifos_3_io_out_ready),
    .io_out_valid(fifos_3_io_out_valid),
    .io_out_bits(fifos_3_io_out_bits)
  );
  FIFO_17 fifos_4 ( // @[FIFOVec.scala 40:19:@40805.4]
    .clock(fifos_4_clock),
    .reset(fifos_4_reset),
    .io_in_ready(fifos_4_io_in_ready),
    .io_in_valid(fifos_4_io_in_valid),
    .io_in_bits(fifos_4_io_in_bits),
    .io_out_ready(fifos_4_io_out_ready),
    .io_out_valid(fifos_4_io_out_valid),
    .io_out_bits(fifos_4_io_out_bits)
  );
  FIFO_17 fifos_5 ( // @[FIFOVec.scala 40:19:@40840.4]
    .clock(fifos_5_clock),
    .reset(fifos_5_reset),
    .io_in_ready(fifos_5_io_in_ready),
    .io_in_valid(fifos_5_io_in_valid),
    .io_in_bits(fifos_5_io_in_bits),
    .io_out_ready(fifos_5_io_out_ready),
    .io_out_valid(fifos_5_io_out_valid),
    .io_out_bits(fifos_5_io_out_bits)
  );
  FIFO_17 fifos_6 ( // @[FIFOVec.scala 40:19:@40875.4]
    .clock(fifos_6_clock),
    .reset(fifos_6_reset),
    .io_in_ready(fifos_6_io_in_ready),
    .io_in_valid(fifos_6_io_in_valid),
    .io_in_bits(fifos_6_io_in_bits),
    .io_out_ready(fifos_6_io_out_ready),
    .io_out_valid(fifos_6_io_out_valid),
    .io_out_bits(fifos_6_io_out_bits)
  );
  FIFO_17 fifos_7 ( // @[FIFOVec.scala 40:19:@40910.4]
    .clock(fifos_7_clock),
    .reset(fifos_7_reset),
    .io_in_ready(fifos_7_io_in_ready),
    .io_in_valid(fifos_7_io_in_valid),
    .io_in_bits(fifos_7_io_in_bits),
    .io_out_ready(fifos_7_io_out_ready),
    .io_out_valid(fifos_7_io_out_valid),
    .io_out_bits(fifos_7_io_out_bits)
  );
  FIFO_17 fifos_8 ( // @[FIFOVec.scala 40:19:@40945.4]
    .clock(fifos_8_clock),
    .reset(fifos_8_reset),
    .io_in_ready(fifos_8_io_in_ready),
    .io_in_valid(fifos_8_io_in_valid),
    .io_in_bits(fifos_8_io_in_bits),
    .io_out_ready(fifos_8_io_out_ready),
    .io_out_valid(fifos_8_io_out_valid),
    .io_out_bits(fifos_8_io_out_bits)
  );
  FIFO_17 fifos_9 ( // @[FIFOVec.scala 40:19:@40980.4]
    .clock(fifos_9_clock),
    .reset(fifos_9_reset),
    .io_in_ready(fifos_9_io_in_ready),
    .io_in_valid(fifos_9_io_in_valid),
    .io_in_bits(fifos_9_io_in_bits),
    .io_out_ready(fifos_9_io_out_ready),
    .io_out_valid(fifos_9_io_out_valid),
    .io_out_bits(fifos_9_io_out_bits)
  );
  FIFO_17 fifos_10 ( // @[FIFOVec.scala 40:19:@41015.4]
    .clock(fifos_10_clock),
    .reset(fifos_10_reset),
    .io_in_ready(fifos_10_io_in_ready),
    .io_in_valid(fifos_10_io_in_valid),
    .io_in_bits(fifos_10_io_in_bits),
    .io_out_ready(fifos_10_io_out_ready),
    .io_out_valid(fifos_10_io_out_valid),
    .io_out_bits(fifos_10_io_out_bits)
  );
  FIFO_17 fifos_11 ( // @[FIFOVec.scala 40:19:@41050.4]
    .clock(fifos_11_clock),
    .reset(fifos_11_reset),
    .io_in_ready(fifos_11_io_in_ready),
    .io_in_valid(fifos_11_io_in_valid),
    .io_in_bits(fifos_11_io_in_bits),
    .io_out_ready(fifos_11_io_out_ready),
    .io_out_valid(fifos_11_io_out_valid),
    .io_out_bits(fifos_11_io_out_bits)
  );
  FIFO_17 fifos_12 ( // @[FIFOVec.scala 40:19:@41085.4]
    .clock(fifos_12_clock),
    .reset(fifos_12_reset),
    .io_in_ready(fifos_12_io_in_ready),
    .io_in_valid(fifos_12_io_in_valid),
    .io_in_bits(fifos_12_io_in_bits),
    .io_out_ready(fifos_12_io_out_ready),
    .io_out_valid(fifos_12_io_out_valid),
    .io_out_bits(fifos_12_io_out_bits)
  );
  FIFO_17 fifos_13 ( // @[FIFOVec.scala 40:19:@41120.4]
    .clock(fifos_13_clock),
    .reset(fifos_13_reset),
    .io_in_ready(fifos_13_io_in_ready),
    .io_in_valid(fifos_13_io_in_valid),
    .io_in_bits(fifos_13_io_in_bits),
    .io_out_ready(fifos_13_io_out_ready),
    .io_out_valid(fifos_13_io_out_valid),
    .io_out_bits(fifos_13_io_out_bits)
  );
  FIFO_17 fifos_14 ( // @[FIFOVec.scala 40:19:@41155.4]
    .clock(fifos_14_clock),
    .reset(fifos_14_reset),
    .io_in_ready(fifos_14_io_in_ready),
    .io_in_valid(fifos_14_io_in_valid),
    .io_in_bits(fifos_14_io_in_bits),
    .io_out_ready(fifos_14_io_out_ready),
    .io_out_valid(fifos_14_io_out_valid),
    .io_out_bits(fifos_14_io_out_bits)
  );
  FIFO_17 fifos_15 ( // @[FIFOVec.scala 40:19:@41190.4]
    .clock(fifos_15_clock),
    .reset(fifos_15_reset),
    .io_in_ready(fifos_15_io_in_ready),
    .io_in_valid(fifos_15_io_in_valid),
    .io_in_bits(fifos_15_io_in_bits),
    .io_out_ready(fifos_15_io_out_ready),
    .io_out_valid(fifos_15_io_out_valid),
    .io_out_bits(fifos_15_io_out_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFOVec.scala 21:29:@40640.4]
  assign enqDecoder = 16'h1 << enqCounter_io_out; // @[OneHot.scala 45:35:@40663.4]
  assign _T_149 = enqDecoder[0]; // @[FIFOVec.scala 42:49:@40690.4]
  assign _T_158 = enqDecoder[1]; // @[FIFOVec.scala 42:49:@40725.4]
  assign _T_167 = enqDecoder[2]; // @[FIFOVec.scala 42:49:@40760.4]
  assign _T_176 = enqDecoder[3]; // @[FIFOVec.scala 42:49:@40795.4]
  assign _T_185 = enqDecoder[4]; // @[FIFOVec.scala 42:49:@40830.4]
  assign _T_194 = enqDecoder[5]; // @[FIFOVec.scala 42:49:@40865.4]
  assign _T_203 = enqDecoder[6]; // @[FIFOVec.scala 42:49:@40900.4]
  assign _T_212 = enqDecoder[7]; // @[FIFOVec.scala 42:49:@40935.4]
  assign _T_221 = enqDecoder[8]; // @[FIFOVec.scala 42:49:@40970.4]
  assign _T_230 = enqDecoder[9]; // @[FIFOVec.scala 42:49:@41005.4]
  assign _T_239 = enqDecoder[10]; // @[FIFOVec.scala 42:49:@41040.4]
  assign _T_248 = enqDecoder[11]; // @[FIFOVec.scala 42:49:@41075.4]
  assign _T_257 = enqDecoder[12]; // @[FIFOVec.scala 42:49:@41110.4]
  assign _T_266 = enqDecoder[13]; // @[FIFOVec.scala 42:49:@41145.4]
  assign _T_275 = enqDecoder[14]; // @[FIFOVec.scala 42:49:@41180.4]
  assign _T_284 = enqDecoder[15]; // @[FIFOVec.scala 42:49:@41215.4]
  assign _T_296_0 = fifos_0_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41226.4]
  assign _T_296_1 = fifos_1_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41227.4]
  assign _GEN_1 = 4'h1 == enqCounter_io_out ? _T_296_1 : _T_296_0; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_2 = fifos_2_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41228.4]
  assign _GEN_2 = 4'h2 == enqCounter_io_out ? _T_296_2 : _GEN_1; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_3 = fifos_3_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41229.4]
  assign _GEN_3 = 4'h3 == enqCounter_io_out ? _T_296_3 : _GEN_2; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_4 = fifos_4_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41230.4]
  assign _GEN_4 = 4'h4 == enqCounter_io_out ? _T_296_4 : _GEN_3; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_5 = fifos_5_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41231.4]
  assign _GEN_5 = 4'h5 == enqCounter_io_out ? _T_296_5 : _GEN_4; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_6 = fifos_6_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41232.4]
  assign _GEN_6 = 4'h6 == enqCounter_io_out ? _T_296_6 : _GEN_5; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_7 = fifos_7_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41233.4]
  assign _GEN_7 = 4'h7 == enqCounter_io_out ? _T_296_7 : _GEN_6; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_8 = fifos_8_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41234.4]
  assign _GEN_8 = 4'h8 == enqCounter_io_out ? _T_296_8 : _GEN_7; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_9 = fifos_9_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41235.4]
  assign _GEN_9 = 4'h9 == enqCounter_io_out ? _T_296_9 : _GEN_8; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_10 = fifos_10_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41236.4]
  assign _GEN_10 = 4'ha == enqCounter_io_out ? _T_296_10 : _GEN_9; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_11 = fifos_11_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41237.4]
  assign _GEN_11 = 4'hb == enqCounter_io_out ? _T_296_11 : _GEN_10; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_12 = fifos_12_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41238.4]
  assign _GEN_12 = 4'hc == enqCounter_io_out ? _T_296_12 : _GEN_11; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_13 = fifos_13_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41239.4]
  assign _GEN_13 = 4'hd == enqCounter_io_out ? _T_296_13 : _GEN_12; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_14 = fifos_14_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41240.4]
  assign _GEN_14 = 4'he == enqCounter_io_out ? _T_296_14 : _GEN_13; // @[FIFOVec.scala 49:21:@41257.4]
  assign _T_296_15 = fifos_15_io_in_ready; // @[FIFOVec.scala 49:42:@41225.4 FIFOVec.scala 49:42:@41241.4]
  assign _T_355 = fifos_0_io_out_valid & fifos_1_io_out_valid; // @[FIFOVec.scala 51:93:@41276.4]
  assign _T_356 = _T_355 & fifos_2_io_out_valid; // @[FIFOVec.scala 51:93:@41277.4]
  assign _T_357 = _T_356 & fifos_3_io_out_valid; // @[FIFOVec.scala 51:93:@41278.4]
  assign _T_358 = _T_357 & fifos_4_io_out_valid; // @[FIFOVec.scala 51:93:@41279.4]
  assign _T_359 = _T_358 & fifos_5_io_out_valid; // @[FIFOVec.scala 51:93:@41280.4]
  assign _T_360 = _T_359 & fifos_6_io_out_valid; // @[FIFOVec.scala 51:93:@41281.4]
  assign _T_361 = _T_360 & fifos_7_io_out_valid; // @[FIFOVec.scala 51:93:@41282.4]
  assign _T_362 = _T_361 & fifos_8_io_out_valid; // @[FIFOVec.scala 51:93:@41283.4]
  assign _T_363 = _T_362 & fifos_9_io_out_valid; // @[FIFOVec.scala 51:93:@41284.4]
  assign _T_364 = _T_363 & fifos_10_io_out_valid; // @[FIFOVec.scala 51:93:@41285.4]
  assign _T_365 = _T_364 & fifos_11_io_out_valid; // @[FIFOVec.scala 51:93:@41286.4]
  assign _T_366 = _T_365 & fifos_12_io_out_valid; // @[FIFOVec.scala 51:93:@41287.4]
  assign _T_367 = _T_366 & fifos_13_io_out_valid; // @[FIFOVec.scala 51:93:@41288.4]
  assign _T_368 = _T_367 & fifos_14_io_out_valid; // @[FIFOVec.scala 51:93:@41289.4]
  assign io_in_ready = 4'hf == enqCounter_io_out ? _T_296_15 : _GEN_14; // @[FIFOVec.scala 49:15:@41258.4]
  assign io_out_valid = _T_368 & fifos_15_io_out_valid; // @[FIFOVec.scala 51:16:@41292.4]
  assign io_out_bits_0 = fifos_0_io_out_bits; // @[FIFOVec.scala 53:15:@41600.4]
  assign io_out_bits_1 = fifos_1_io_out_bits; // @[FIFOVec.scala 53:15:@41601.4]
  assign io_out_bits_2 = fifos_2_io_out_bits; // @[FIFOVec.scala 53:15:@41602.4]
  assign io_out_bits_3 = fifos_3_io_out_bits; // @[FIFOVec.scala 53:15:@41603.4]
  assign io_out_bits_4 = fifos_4_io_out_bits; // @[FIFOVec.scala 53:15:@41604.4]
  assign io_out_bits_5 = fifos_5_io_out_bits; // @[FIFOVec.scala 53:15:@41605.4]
  assign io_out_bits_6 = fifos_6_io_out_bits; // @[FIFOVec.scala 53:15:@41606.4]
  assign io_out_bits_7 = fifos_7_io_out_bits; // @[FIFOVec.scala 53:15:@41607.4]
  assign io_out_bits_8 = fifos_8_io_out_bits; // @[FIFOVec.scala 53:15:@41608.4]
  assign io_out_bits_9 = fifos_9_io_out_bits; // @[FIFOVec.scala 53:15:@41609.4]
  assign io_out_bits_10 = fifos_10_io_out_bits; // @[FIFOVec.scala 53:15:@41610.4]
  assign io_out_bits_11 = fifos_11_io_out_bits; // @[FIFOVec.scala 53:15:@41611.4]
  assign io_out_bits_12 = fifos_12_io_out_bits; // @[FIFOVec.scala 53:15:@41612.4]
  assign io_out_bits_13 = fifos_13_io_out_bits; // @[FIFOVec.scala 53:15:@41613.4]
  assign io_out_bits_14 = fifos_14_io_out_bits; // @[FIFOVec.scala 53:15:@41614.4]
  assign io_out_bits_15 = fifos_15_io_out_bits; // @[FIFOVec.scala 53:15:@41615.4]
  assign enqCounter_clock = clock; // @[:@40642.4]
  assign enqCounter_reset = reset; // @[:@40643.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFOVec.scala 26:24:@40650.4]
  assign deqCounter_clock = clock; // @[:@40653.4]
  assign deqCounter_reset = reset; // @[:@40654.4]
  assign deqCounter_io_enable = 1'h0; // @[FIFOVec.scala 30:24:@40661.4]
  assign fifos_0_clock = clock; // @[:@40666.4]
  assign fifos_0_reset = reset; // @[:@40667.4]
  assign fifos_0_io_in_valid = _T_149 & writeEn; // @[FIFOVec.scala 42:19:@40693.4]
  assign fifos_0_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40695.4]
  assign fifos_0_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40699.4]
  assign fifos_1_clock = clock; // @[:@40701.4]
  assign fifos_1_reset = reset; // @[:@40702.4]
  assign fifos_1_io_in_valid = _T_158 & writeEn; // @[FIFOVec.scala 42:19:@40728.4]
  assign fifos_1_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40730.4]
  assign fifos_1_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40734.4]
  assign fifos_2_clock = clock; // @[:@40736.4]
  assign fifos_2_reset = reset; // @[:@40737.4]
  assign fifos_2_io_in_valid = _T_167 & writeEn; // @[FIFOVec.scala 42:19:@40763.4]
  assign fifos_2_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40765.4]
  assign fifos_2_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40769.4]
  assign fifos_3_clock = clock; // @[:@40771.4]
  assign fifos_3_reset = reset; // @[:@40772.4]
  assign fifos_3_io_in_valid = _T_176 & writeEn; // @[FIFOVec.scala 42:19:@40798.4]
  assign fifos_3_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40800.4]
  assign fifos_3_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40804.4]
  assign fifos_4_clock = clock; // @[:@40806.4]
  assign fifos_4_reset = reset; // @[:@40807.4]
  assign fifos_4_io_in_valid = _T_185 & writeEn; // @[FIFOVec.scala 42:19:@40833.4]
  assign fifos_4_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40835.4]
  assign fifos_4_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40839.4]
  assign fifos_5_clock = clock; // @[:@40841.4]
  assign fifos_5_reset = reset; // @[:@40842.4]
  assign fifos_5_io_in_valid = _T_194 & writeEn; // @[FIFOVec.scala 42:19:@40868.4]
  assign fifos_5_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40870.4]
  assign fifos_5_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40874.4]
  assign fifos_6_clock = clock; // @[:@40876.4]
  assign fifos_6_reset = reset; // @[:@40877.4]
  assign fifos_6_io_in_valid = _T_203 & writeEn; // @[FIFOVec.scala 42:19:@40903.4]
  assign fifos_6_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40905.4]
  assign fifos_6_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40909.4]
  assign fifos_7_clock = clock; // @[:@40911.4]
  assign fifos_7_reset = reset; // @[:@40912.4]
  assign fifos_7_io_in_valid = _T_212 & writeEn; // @[FIFOVec.scala 42:19:@40938.4]
  assign fifos_7_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40940.4]
  assign fifos_7_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40944.4]
  assign fifos_8_clock = clock; // @[:@40946.4]
  assign fifos_8_reset = reset; // @[:@40947.4]
  assign fifos_8_io_in_valid = _T_221 & writeEn; // @[FIFOVec.scala 42:19:@40973.4]
  assign fifos_8_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@40975.4]
  assign fifos_8_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@40979.4]
  assign fifos_9_clock = clock; // @[:@40981.4]
  assign fifos_9_reset = reset; // @[:@40982.4]
  assign fifos_9_io_in_valid = _T_230 & writeEn; // @[FIFOVec.scala 42:19:@41008.4]
  assign fifos_9_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41010.4]
  assign fifos_9_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41014.4]
  assign fifos_10_clock = clock; // @[:@41016.4]
  assign fifos_10_reset = reset; // @[:@41017.4]
  assign fifos_10_io_in_valid = _T_239 & writeEn; // @[FIFOVec.scala 42:19:@41043.4]
  assign fifos_10_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41045.4]
  assign fifos_10_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41049.4]
  assign fifos_11_clock = clock; // @[:@41051.4]
  assign fifos_11_reset = reset; // @[:@41052.4]
  assign fifos_11_io_in_valid = _T_248 & writeEn; // @[FIFOVec.scala 42:19:@41078.4]
  assign fifos_11_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41080.4]
  assign fifos_11_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41084.4]
  assign fifos_12_clock = clock; // @[:@41086.4]
  assign fifos_12_reset = reset; // @[:@41087.4]
  assign fifos_12_io_in_valid = _T_257 & writeEn; // @[FIFOVec.scala 42:19:@41113.4]
  assign fifos_12_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41115.4]
  assign fifos_12_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41119.4]
  assign fifos_13_clock = clock; // @[:@41121.4]
  assign fifos_13_reset = reset; // @[:@41122.4]
  assign fifos_13_io_in_valid = _T_266 & writeEn; // @[FIFOVec.scala 42:19:@41148.4]
  assign fifos_13_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41150.4]
  assign fifos_13_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41154.4]
  assign fifos_14_clock = clock; // @[:@41156.4]
  assign fifos_14_reset = reset; // @[:@41157.4]
  assign fifos_14_io_in_valid = _T_275 & writeEn; // @[FIFOVec.scala 42:19:@41183.4]
  assign fifos_14_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41185.4]
  assign fifos_14_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41189.4]
  assign fifos_15_clock = clock; // @[:@41191.4]
  assign fifos_15_reset = reset; // @[:@41192.4]
  assign fifos_15_io_in_valid = _T_284 & writeEn; // @[FIFOVec.scala 42:19:@41218.4]
  assign fifos_15_io_in_bits = io_in_bits_0; // @[FIFOVec.scala 43:18:@41220.4]
  assign fifos_15_io_out_ready = io_out_valid & io_out_ready; // @[FIFOVec.scala 44:20:@41224.4]
endmodule
module FIFOWidthConvert( // @[:@41617.2]
  input         clock, // @[:@41618.4]
  input         reset, // @[:@41619.4]
  output        io_in_ready, // @[:@41620.4]
  input         io_in_valid, // @[:@41620.4]
  input  [31:0] io_in_bits_data_0, // @[:@41620.4]
  input         io_in_bits_strobe, // @[:@41620.4]
  input         io_out_ready, // @[:@41620.4]
  output        io_out_valid, // @[:@41620.4]
  output [31:0] io_out_bits_data_0, // @[:@41620.4]
  output [31:0] io_out_bits_data_1, // @[:@41620.4]
  output [31:0] io_out_bits_data_2, // @[:@41620.4]
  output [31:0] io_out_bits_data_3, // @[:@41620.4]
  output [31:0] io_out_bits_data_4, // @[:@41620.4]
  output [31:0] io_out_bits_data_5, // @[:@41620.4]
  output [31:0] io_out_bits_data_6, // @[:@41620.4]
  output [31:0] io_out_bits_data_7, // @[:@41620.4]
  output [31:0] io_out_bits_data_8, // @[:@41620.4]
  output [31:0] io_out_bits_data_9, // @[:@41620.4]
  output [31:0] io_out_bits_data_10, // @[:@41620.4]
  output [31:0] io_out_bits_data_11, // @[:@41620.4]
  output [31:0] io_out_bits_data_12, // @[:@41620.4]
  output [31:0] io_out_bits_data_13, // @[:@41620.4]
  output [31:0] io_out_bits_data_14, // @[:@41620.4]
  output [31:0] io_out_bits_data_15, // @[:@41620.4]
  output [63:0] io_out_bits_strobe // @[:@41620.4]
);
  wire  FIFOVec_clock; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire  FIFOVec_reset; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire  FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire  FIFOVec_io_in_valid; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_in_bits_0; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire  FIFOVec_io_out_ready; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire  FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_0; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_1; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_2; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_3; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_4; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_5; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_6; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_7; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_8; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_9; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_10; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_11; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_12; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_13; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_14; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire [31:0] FIFOVec_io_out_bits_15; // @[FIFOWidthConvert.scala 61:22:@41622.4]
  wire  FIFOVec_1_clock; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_reset; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_in_ready; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_in_valid; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_in_bits_0; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_ready; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_valid; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_0; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_1; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_2; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_3; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_4; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_5; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_6; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_7; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_8; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_9; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_10; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_11; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_12; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_13; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_14; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire  FIFOVec_1_io_out_bits_15; // @[FIFOWidthConvert.scala 62:26:@41663.4]
  wire [319:0] _T_55; // @[Cat.scala 30:58:@41722.4]
  wire [511:0] _T_61; // @[Cat.scala 30:58:@41728.4]
  wire [9:0] _T_108; // @[Cat.scala 30:58:@41786.4]
  wire [15:0] _T_114; // @[Cat.scala 30:58:@41792.4]
  wire  _T_115; // @[FIFOWidthConvert.scala 36:14:@41793.4]
  wire  _T_119; // @[FIFOWidthConvert.scala 36:14:@41797.4]
  wire  _T_123; // @[FIFOWidthConvert.scala 36:14:@41801.4]
  wire  _T_127; // @[FIFOWidthConvert.scala 36:14:@41805.4]
  wire  _T_131; // @[FIFOWidthConvert.scala 36:14:@41809.4]
  wire  _T_135; // @[FIFOWidthConvert.scala 36:14:@41813.4]
  wire  _T_139; // @[FIFOWidthConvert.scala 36:14:@41817.4]
  wire  _T_143; // @[FIFOWidthConvert.scala 36:14:@41821.4]
  wire  _T_147; // @[FIFOWidthConvert.scala 36:14:@41825.4]
  wire  _T_151; // @[FIFOWidthConvert.scala 36:14:@41829.4]
  wire  _T_155; // @[FIFOWidthConvert.scala 36:14:@41833.4]
  wire  _T_159; // @[FIFOWidthConvert.scala 36:14:@41837.4]
  wire  _T_163; // @[FIFOWidthConvert.scala 36:14:@41841.4]
  wire  _T_167; // @[FIFOWidthConvert.scala 36:14:@41845.4]
  wire  _T_171; // @[FIFOWidthConvert.scala 36:14:@41849.4]
  wire  _T_175; // @[FIFOWidthConvert.scala 36:14:@41853.4]
  wire [9:0] _T_257; // @[Cat.scala 30:58:@41930.4]
  wire [18:0] _T_266; // @[Cat.scala 30:58:@41939.4]
  wire [27:0] _T_275; // @[Cat.scala 30:58:@41948.4]
  wire [36:0] _T_284; // @[Cat.scala 30:58:@41957.4]
  wire [45:0] _T_293; // @[Cat.scala 30:58:@41966.4]
  wire [54:0] _T_302; // @[Cat.scala 30:58:@41975.4]
  wire [62:0] _T_310; // @[Cat.scala 30:58:@41983.4]
  FIFOVec FIFOVec ( // @[FIFOWidthConvert.scala 61:22:@41622.4]
    .clock(FIFOVec_clock),
    .reset(FIFOVec_reset),
    .io_in_ready(FIFOVec_io_in_ready),
    .io_in_valid(FIFOVec_io_in_valid),
    .io_in_bits_0(FIFOVec_io_in_bits_0),
    .io_out_ready(FIFOVec_io_out_ready),
    .io_out_valid(FIFOVec_io_out_valid),
    .io_out_bits_0(FIFOVec_io_out_bits_0),
    .io_out_bits_1(FIFOVec_io_out_bits_1),
    .io_out_bits_2(FIFOVec_io_out_bits_2),
    .io_out_bits_3(FIFOVec_io_out_bits_3),
    .io_out_bits_4(FIFOVec_io_out_bits_4),
    .io_out_bits_5(FIFOVec_io_out_bits_5),
    .io_out_bits_6(FIFOVec_io_out_bits_6),
    .io_out_bits_7(FIFOVec_io_out_bits_7),
    .io_out_bits_8(FIFOVec_io_out_bits_8),
    .io_out_bits_9(FIFOVec_io_out_bits_9),
    .io_out_bits_10(FIFOVec_io_out_bits_10),
    .io_out_bits_11(FIFOVec_io_out_bits_11),
    .io_out_bits_12(FIFOVec_io_out_bits_12),
    .io_out_bits_13(FIFOVec_io_out_bits_13),
    .io_out_bits_14(FIFOVec_io_out_bits_14),
    .io_out_bits_15(FIFOVec_io_out_bits_15)
  );
  FIFOVec_1 FIFOVec_1 ( // @[FIFOWidthConvert.scala 62:26:@41663.4]
    .clock(FIFOVec_1_clock),
    .reset(FIFOVec_1_reset),
    .io_in_ready(FIFOVec_1_io_in_ready),
    .io_in_valid(FIFOVec_1_io_in_valid),
    .io_in_bits_0(FIFOVec_1_io_in_bits_0),
    .io_out_ready(FIFOVec_1_io_out_ready),
    .io_out_valid(FIFOVec_1_io_out_valid),
    .io_out_bits_0(FIFOVec_1_io_out_bits_0),
    .io_out_bits_1(FIFOVec_1_io_out_bits_1),
    .io_out_bits_2(FIFOVec_1_io_out_bits_2),
    .io_out_bits_3(FIFOVec_1_io_out_bits_3),
    .io_out_bits_4(FIFOVec_1_io_out_bits_4),
    .io_out_bits_5(FIFOVec_1_io_out_bits_5),
    .io_out_bits_6(FIFOVec_1_io_out_bits_6),
    .io_out_bits_7(FIFOVec_1_io_out_bits_7),
    .io_out_bits_8(FIFOVec_1_io_out_bits_8),
    .io_out_bits_9(FIFOVec_1_io_out_bits_9),
    .io_out_bits_10(FIFOVec_1_io_out_bits_10),
    .io_out_bits_11(FIFOVec_1_io_out_bits_11),
    .io_out_bits_12(FIFOVec_1_io_out_bits_12),
    .io_out_bits_13(FIFOVec_1_io_out_bits_13),
    .io_out_bits_14(FIFOVec_1_io_out_bits_14),
    .io_out_bits_15(FIFOVec_1_io_out_bits_15)
  );
  assign _T_55 = {FIFOVec_io_out_bits_15,FIFOVec_io_out_bits_14,FIFOVec_io_out_bits_13,FIFOVec_io_out_bits_12,FIFOVec_io_out_bits_11,FIFOVec_io_out_bits_10,FIFOVec_io_out_bits_9,FIFOVec_io_out_bits_8,FIFOVec_io_out_bits_7,FIFOVec_io_out_bits_6}; // @[Cat.scala 30:58:@41722.4]
  assign _T_61 = {_T_55,FIFOVec_io_out_bits_5,FIFOVec_io_out_bits_4,FIFOVec_io_out_bits_3,FIFOVec_io_out_bits_2,FIFOVec_io_out_bits_1,FIFOVec_io_out_bits_0}; // @[Cat.scala 30:58:@41728.4]
  assign _T_108 = {FIFOVec_1_io_out_bits_0,FIFOVec_1_io_out_bits_1,FIFOVec_1_io_out_bits_2,FIFOVec_1_io_out_bits_3,FIFOVec_1_io_out_bits_4,FIFOVec_1_io_out_bits_5,FIFOVec_1_io_out_bits_6,FIFOVec_1_io_out_bits_7,FIFOVec_1_io_out_bits_8,FIFOVec_1_io_out_bits_9}; // @[Cat.scala 30:58:@41786.4]
  assign _T_114 = {_T_108,FIFOVec_1_io_out_bits_10,FIFOVec_1_io_out_bits_11,FIFOVec_1_io_out_bits_12,FIFOVec_1_io_out_bits_13,FIFOVec_1_io_out_bits_14,FIFOVec_1_io_out_bits_15}; // @[Cat.scala 30:58:@41792.4]
  assign _T_115 = _T_114[0]; // @[FIFOWidthConvert.scala 36:14:@41793.4]
  assign _T_119 = _T_114[1]; // @[FIFOWidthConvert.scala 36:14:@41797.4]
  assign _T_123 = _T_114[2]; // @[FIFOWidthConvert.scala 36:14:@41801.4]
  assign _T_127 = _T_114[3]; // @[FIFOWidthConvert.scala 36:14:@41805.4]
  assign _T_131 = _T_114[4]; // @[FIFOWidthConvert.scala 36:14:@41809.4]
  assign _T_135 = _T_114[5]; // @[FIFOWidthConvert.scala 36:14:@41813.4]
  assign _T_139 = _T_114[6]; // @[FIFOWidthConvert.scala 36:14:@41817.4]
  assign _T_143 = _T_114[7]; // @[FIFOWidthConvert.scala 36:14:@41821.4]
  assign _T_147 = _T_114[8]; // @[FIFOWidthConvert.scala 36:14:@41825.4]
  assign _T_151 = _T_114[9]; // @[FIFOWidthConvert.scala 36:14:@41829.4]
  assign _T_155 = _T_114[10]; // @[FIFOWidthConvert.scala 36:14:@41833.4]
  assign _T_159 = _T_114[11]; // @[FIFOWidthConvert.scala 36:14:@41837.4]
  assign _T_163 = _T_114[12]; // @[FIFOWidthConvert.scala 36:14:@41841.4]
  assign _T_167 = _T_114[13]; // @[FIFOWidthConvert.scala 36:14:@41845.4]
  assign _T_171 = _T_114[14]; // @[FIFOWidthConvert.scala 36:14:@41849.4]
  assign _T_175 = _T_114[15]; // @[FIFOWidthConvert.scala 36:14:@41853.4]
  assign _T_257 = {_T_175,_T_175,_T_175,_T_175,_T_171,_T_171,_T_171,_T_171,_T_167,_T_167}; // @[Cat.scala 30:58:@41930.4]
  assign _T_266 = {_T_257,_T_167,_T_167,_T_163,_T_163,_T_163,_T_163,_T_159,_T_159,_T_159}; // @[Cat.scala 30:58:@41939.4]
  assign _T_275 = {_T_266,_T_159,_T_155,_T_155,_T_155,_T_155,_T_151,_T_151,_T_151,_T_151}; // @[Cat.scala 30:58:@41948.4]
  assign _T_284 = {_T_275,_T_147,_T_147,_T_147,_T_147,_T_143,_T_143,_T_143,_T_143,_T_139}; // @[Cat.scala 30:58:@41957.4]
  assign _T_293 = {_T_284,_T_139,_T_139,_T_139,_T_135,_T_135,_T_135,_T_135,_T_131,_T_131}; // @[Cat.scala 30:58:@41966.4]
  assign _T_302 = {_T_293,_T_131,_T_131,_T_127,_T_127,_T_127,_T_127,_T_123,_T_123,_T_123}; // @[Cat.scala 30:58:@41975.4]
  assign _T_310 = {_T_302,_T_123,_T_119,_T_119,_T_119,_T_119,_T_115,_T_115,_T_115}; // @[Cat.scala 30:58:@41983.4]
  assign io_in_ready = FIFOVec_io_in_ready; // @[FIFOWidthConvert.scala 71:17:@41712.4]
  assign io_out_valid = FIFOVec_io_out_valid; // @[FIFOWidthConvert.scala 72:18:@41713.4]
  assign io_out_bits_data_0 = _T_61[31:0]; // @[FIFOWidthConvert.scala 73:22:@41762.4]
  assign io_out_bits_data_1 = _T_61[63:32]; // @[FIFOWidthConvert.scala 73:22:@41763.4]
  assign io_out_bits_data_2 = _T_61[95:64]; // @[FIFOWidthConvert.scala 73:22:@41764.4]
  assign io_out_bits_data_3 = _T_61[127:96]; // @[FIFOWidthConvert.scala 73:22:@41765.4]
  assign io_out_bits_data_4 = _T_61[159:128]; // @[FIFOWidthConvert.scala 73:22:@41766.4]
  assign io_out_bits_data_5 = _T_61[191:160]; // @[FIFOWidthConvert.scala 73:22:@41767.4]
  assign io_out_bits_data_6 = _T_61[223:192]; // @[FIFOWidthConvert.scala 73:22:@41768.4]
  assign io_out_bits_data_7 = _T_61[255:224]; // @[FIFOWidthConvert.scala 73:22:@41769.4]
  assign io_out_bits_data_8 = _T_61[287:256]; // @[FIFOWidthConvert.scala 73:22:@41770.4]
  assign io_out_bits_data_9 = _T_61[319:288]; // @[FIFOWidthConvert.scala 73:22:@41771.4]
  assign io_out_bits_data_10 = _T_61[351:320]; // @[FIFOWidthConvert.scala 73:22:@41772.4]
  assign io_out_bits_data_11 = _T_61[383:352]; // @[FIFOWidthConvert.scala 73:22:@41773.4]
  assign io_out_bits_data_12 = _T_61[415:384]; // @[FIFOWidthConvert.scala 73:22:@41774.4]
  assign io_out_bits_data_13 = _T_61[447:416]; // @[FIFOWidthConvert.scala 73:22:@41775.4]
  assign io_out_bits_data_14 = _T_61[479:448]; // @[FIFOWidthConvert.scala 73:22:@41776.4]
  assign io_out_bits_data_15 = _T_61[511:480]; // @[FIFOWidthConvert.scala 73:22:@41777.4]
  assign io_out_bits_strobe = {_T_310,_T_115}; // @[FIFOWidthConvert.scala 74:24:@41985.4]
  assign FIFOVec_clock = clock; // @[:@41623.4]
  assign FIFOVec_reset = reset; // @[:@41624.4]
  assign FIFOVec_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 68:22:@41709.4]
  assign FIFOVec_io_in_bits_0 = io_in_bits_data_0; // @[FIFOWidthConvert.scala 67:24:@41708.4]
  assign FIFOVec_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 75:23:@41986.4]
  assign FIFOVec_1_clock = clock; // @[:@41664.4]
  assign FIFOVec_1_reset = reset; // @[:@41665.4]
  assign FIFOVec_1_io_in_valid = io_in_valid; // @[FIFOWidthConvert.scala 70:26:@41711.4]
  assign FIFOVec_1_io_in_bits_0 = io_in_bits_strobe; // @[FIFOWidthConvert.scala 69:28:@41710.4]
  assign FIFOVec_1_io_out_ready = io_out_ready; // @[FIFOWidthConvert.scala 76:27:@41987.4]
endmodule
module FFRAM_16( // @[:@42025.2]
  input        clock, // @[:@42026.4]
  input        reset, // @[:@42027.4]
  input  [5:0] io_raddr, // @[:@42028.4]
  input        io_wen, // @[:@42028.4]
  input  [5:0] io_waddr, // @[:@42028.4]
  input        io_wdata, // @[:@42028.4]
  output       io_rdata, // @[:@42028.4]
  input        io_banks_0_wdata_valid, // @[:@42028.4]
  input        io_banks_0_wdata_bits, // @[:@42028.4]
  input        io_banks_1_wdata_valid, // @[:@42028.4]
  input        io_banks_1_wdata_bits, // @[:@42028.4]
  input        io_banks_2_wdata_valid, // @[:@42028.4]
  input        io_banks_2_wdata_bits, // @[:@42028.4]
  input        io_banks_3_wdata_valid, // @[:@42028.4]
  input        io_banks_3_wdata_bits, // @[:@42028.4]
  input        io_banks_4_wdata_valid, // @[:@42028.4]
  input        io_banks_4_wdata_bits, // @[:@42028.4]
  input        io_banks_5_wdata_valid, // @[:@42028.4]
  input        io_banks_5_wdata_bits, // @[:@42028.4]
  input        io_banks_6_wdata_valid, // @[:@42028.4]
  input        io_banks_6_wdata_bits, // @[:@42028.4]
  input        io_banks_7_wdata_valid, // @[:@42028.4]
  input        io_banks_7_wdata_bits, // @[:@42028.4]
  input        io_banks_8_wdata_valid, // @[:@42028.4]
  input        io_banks_8_wdata_bits, // @[:@42028.4]
  input        io_banks_9_wdata_valid, // @[:@42028.4]
  input        io_banks_9_wdata_bits, // @[:@42028.4]
  input        io_banks_10_wdata_valid, // @[:@42028.4]
  input        io_banks_10_wdata_bits, // @[:@42028.4]
  input        io_banks_11_wdata_valid, // @[:@42028.4]
  input        io_banks_11_wdata_bits, // @[:@42028.4]
  input        io_banks_12_wdata_valid, // @[:@42028.4]
  input        io_banks_12_wdata_bits, // @[:@42028.4]
  input        io_banks_13_wdata_valid, // @[:@42028.4]
  input        io_banks_13_wdata_bits, // @[:@42028.4]
  input        io_banks_14_wdata_valid, // @[:@42028.4]
  input        io_banks_14_wdata_bits, // @[:@42028.4]
  input        io_banks_15_wdata_valid, // @[:@42028.4]
  input        io_banks_15_wdata_bits, // @[:@42028.4]
  input        io_banks_16_wdata_valid, // @[:@42028.4]
  input        io_banks_16_wdata_bits, // @[:@42028.4]
  input        io_banks_17_wdata_valid, // @[:@42028.4]
  input        io_banks_17_wdata_bits, // @[:@42028.4]
  input        io_banks_18_wdata_valid, // @[:@42028.4]
  input        io_banks_18_wdata_bits, // @[:@42028.4]
  input        io_banks_19_wdata_valid, // @[:@42028.4]
  input        io_banks_19_wdata_bits, // @[:@42028.4]
  input        io_banks_20_wdata_valid, // @[:@42028.4]
  input        io_banks_20_wdata_bits, // @[:@42028.4]
  input        io_banks_21_wdata_valid, // @[:@42028.4]
  input        io_banks_21_wdata_bits, // @[:@42028.4]
  input        io_banks_22_wdata_valid, // @[:@42028.4]
  input        io_banks_22_wdata_bits, // @[:@42028.4]
  input        io_banks_23_wdata_valid, // @[:@42028.4]
  input        io_banks_23_wdata_bits, // @[:@42028.4]
  input        io_banks_24_wdata_valid, // @[:@42028.4]
  input        io_banks_24_wdata_bits, // @[:@42028.4]
  input        io_banks_25_wdata_valid, // @[:@42028.4]
  input        io_banks_25_wdata_bits, // @[:@42028.4]
  input        io_banks_26_wdata_valid, // @[:@42028.4]
  input        io_banks_26_wdata_bits, // @[:@42028.4]
  input        io_banks_27_wdata_valid, // @[:@42028.4]
  input        io_banks_27_wdata_bits, // @[:@42028.4]
  input        io_banks_28_wdata_valid, // @[:@42028.4]
  input        io_banks_28_wdata_bits, // @[:@42028.4]
  input        io_banks_29_wdata_valid, // @[:@42028.4]
  input        io_banks_29_wdata_bits, // @[:@42028.4]
  input        io_banks_30_wdata_valid, // @[:@42028.4]
  input        io_banks_30_wdata_bits, // @[:@42028.4]
  input        io_banks_31_wdata_valid, // @[:@42028.4]
  input        io_banks_31_wdata_bits, // @[:@42028.4]
  input        io_banks_32_wdata_valid, // @[:@42028.4]
  input        io_banks_32_wdata_bits, // @[:@42028.4]
  input        io_banks_33_wdata_valid, // @[:@42028.4]
  input        io_banks_33_wdata_bits, // @[:@42028.4]
  input        io_banks_34_wdata_valid, // @[:@42028.4]
  input        io_banks_34_wdata_bits, // @[:@42028.4]
  input        io_banks_35_wdata_valid, // @[:@42028.4]
  input        io_banks_35_wdata_bits, // @[:@42028.4]
  input        io_banks_36_wdata_valid, // @[:@42028.4]
  input        io_banks_36_wdata_bits, // @[:@42028.4]
  input        io_banks_37_wdata_valid, // @[:@42028.4]
  input        io_banks_37_wdata_bits, // @[:@42028.4]
  input        io_banks_38_wdata_valid, // @[:@42028.4]
  input        io_banks_38_wdata_bits, // @[:@42028.4]
  input        io_banks_39_wdata_valid, // @[:@42028.4]
  input        io_banks_39_wdata_bits, // @[:@42028.4]
  input        io_banks_40_wdata_valid, // @[:@42028.4]
  input        io_banks_40_wdata_bits, // @[:@42028.4]
  input        io_banks_41_wdata_valid, // @[:@42028.4]
  input        io_banks_41_wdata_bits, // @[:@42028.4]
  input        io_banks_42_wdata_valid, // @[:@42028.4]
  input        io_banks_42_wdata_bits, // @[:@42028.4]
  input        io_banks_43_wdata_valid, // @[:@42028.4]
  input        io_banks_43_wdata_bits, // @[:@42028.4]
  input        io_banks_44_wdata_valid, // @[:@42028.4]
  input        io_banks_44_wdata_bits, // @[:@42028.4]
  input        io_banks_45_wdata_valid, // @[:@42028.4]
  input        io_banks_45_wdata_bits, // @[:@42028.4]
  input        io_banks_46_wdata_valid, // @[:@42028.4]
  input        io_banks_46_wdata_bits, // @[:@42028.4]
  input        io_banks_47_wdata_valid, // @[:@42028.4]
  input        io_banks_47_wdata_bits, // @[:@42028.4]
  input        io_banks_48_wdata_valid, // @[:@42028.4]
  input        io_banks_48_wdata_bits, // @[:@42028.4]
  input        io_banks_49_wdata_valid, // @[:@42028.4]
  input        io_banks_49_wdata_bits, // @[:@42028.4]
  input        io_banks_50_wdata_valid, // @[:@42028.4]
  input        io_banks_50_wdata_bits, // @[:@42028.4]
  input        io_banks_51_wdata_valid, // @[:@42028.4]
  input        io_banks_51_wdata_bits, // @[:@42028.4]
  input        io_banks_52_wdata_valid, // @[:@42028.4]
  input        io_banks_52_wdata_bits, // @[:@42028.4]
  input        io_banks_53_wdata_valid, // @[:@42028.4]
  input        io_banks_53_wdata_bits, // @[:@42028.4]
  input        io_banks_54_wdata_valid, // @[:@42028.4]
  input        io_banks_54_wdata_bits, // @[:@42028.4]
  input        io_banks_55_wdata_valid, // @[:@42028.4]
  input        io_banks_55_wdata_bits, // @[:@42028.4]
  input        io_banks_56_wdata_valid, // @[:@42028.4]
  input        io_banks_56_wdata_bits, // @[:@42028.4]
  input        io_banks_57_wdata_valid, // @[:@42028.4]
  input        io_banks_57_wdata_bits, // @[:@42028.4]
  input        io_banks_58_wdata_valid, // @[:@42028.4]
  input        io_banks_58_wdata_bits, // @[:@42028.4]
  input        io_banks_59_wdata_valid, // @[:@42028.4]
  input        io_banks_59_wdata_bits, // @[:@42028.4]
  input        io_banks_60_wdata_valid, // @[:@42028.4]
  input        io_banks_60_wdata_bits, // @[:@42028.4]
  input        io_banks_61_wdata_valid, // @[:@42028.4]
  input        io_banks_61_wdata_bits, // @[:@42028.4]
  input        io_banks_62_wdata_valid, // @[:@42028.4]
  input        io_banks_62_wdata_bits, // @[:@42028.4]
  input        io_banks_63_wdata_valid, // @[:@42028.4]
  input        io_banks_63_wdata_bits // @[:@42028.4]
);
  reg  regs_0; // @[SRAM.scala 145:20:@42032.4]
  reg [31:0] _RAND_0;
  wire  _T_688; // @[SRAM.scala 148:37:@42033.4]
  wire  _T_689; // @[SRAM.scala 148:25:@42034.4]
  wire  _T_690; // @[SRAM.scala 148:15:@42035.4]
  wire  _T_691; // @[SRAM.scala 149:15:@42037.6]
  wire  _GEN_0; // @[SRAM.scala 148:48:@42036.4]
  reg  regs_1; // @[SRAM.scala 145:20:@42043.4]
  reg [31:0] _RAND_1;
  wire  _T_697; // @[SRAM.scala 148:37:@42044.4]
  wire  _T_698; // @[SRAM.scala 148:25:@42045.4]
  wire  _T_699; // @[SRAM.scala 148:15:@42046.4]
  wire  _T_700; // @[SRAM.scala 149:15:@42048.6]
  wire  _GEN_1; // @[SRAM.scala 148:48:@42047.4]
  reg  regs_2; // @[SRAM.scala 145:20:@42054.4]
  reg [31:0] _RAND_2;
  wire  _T_706; // @[SRAM.scala 148:37:@42055.4]
  wire  _T_707; // @[SRAM.scala 148:25:@42056.4]
  wire  _T_708; // @[SRAM.scala 148:15:@42057.4]
  wire  _T_709; // @[SRAM.scala 149:15:@42059.6]
  wire  _GEN_2; // @[SRAM.scala 148:48:@42058.4]
  reg  regs_3; // @[SRAM.scala 145:20:@42065.4]
  reg [31:0] _RAND_3;
  wire  _T_715; // @[SRAM.scala 148:37:@42066.4]
  wire  _T_716; // @[SRAM.scala 148:25:@42067.4]
  wire  _T_717; // @[SRAM.scala 148:15:@42068.4]
  wire  _T_718; // @[SRAM.scala 149:15:@42070.6]
  wire  _GEN_3; // @[SRAM.scala 148:48:@42069.4]
  reg  regs_4; // @[SRAM.scala 145:20:@42076.4]
  reg [31:0] _RAND_4;
  wire  _T_724; // @[SRAM.scala 148:37:@42077.4]
  wire  _T_725; // @[SRAM.scala 148:25:@42078.4]
  wire  _T_726; // @[SRAM.scala 148:15:@42079.4]
  wire  _T_727; // @[SRAM.scala 149:15:@42081.6]
  wire  _GEN_4; // @[SRAM.scala 148:48:@42080.4]
  reg  regs_5; // @[SRAM.scala 145:20:@42087.4]
  reg [31:0] _RAND_5;
  wire  _T_733; // @[SRAM.scala 148:37:@42088.4]
  wire  _T_734; // @[SRAM.scala 148:25:@42089.4]
  wire  _T_735; // @[SRAM.scala 148:15:@42090.4]
  wire  _T_736; // @[SRAM.scala 149:15:@42092.6]
  wire  _GEN_5; // @[SRAM.scala 148:48:@42091.4]
  reg  regs_6; // @[SRAM.scala 145:20:@42098.4]
  reg [31:0] _RAND_6;
  wire  _T_742; // @[SRAM.scala 148:37:@42099.4]
  wire  _T_743; // @[SRAM.scala 148:25:@42100.4]
  wire  _T_744; // @[SRAM.scala 148:15:@42101.4]
  wire  _T_745; // @[SRAM.scala 149:15:@42103.6]
  wire  _GEN_6; // @[SRAM.scala 148:48:@42102.4]
  reg  regs_7; // @[SRAM.scala 145:20:@42109.4]
  reg [31:0] _RAND_7;
  wire  _T_751; // @[SRAM.scala 148:37:@42110.4]
  wire  _T_752; // @[SRAM.scala 148:25:@42111.4]
  wire  _T_753; // @[SRAM.scala 148:15:@42112.4]
  wire  _T_754; // @[SRAM.scala 149:15:@42114.6]
  wire  _GEN_7; // @[SRAM.scala 148:48:@42113.4]
  reg  regs_8; // @[SRAM.scala 145:20:@42120.4]
  reg [31:0] _RAND_8;
  wire  _T_760; // @[SRAM.scala 148:37:@42121.4]
  wire  _T_761; // @[SRAM.scala 148:25:@42122.4]
  wire  _T_762; // @[SRAM.scala 148:15:@42123.4]
  wire  _T_763; // @[SRAM.scala 149:15:@42125.6]
  wire  _GEN_8; // @[SRAM.scala 148:48:@42124.4]
  reg  regs_9; // @[SRAM.scala 145:20:@42131.4]
  reg [31:0] _RAND_9;
  wire  _T_769; // @[SRAM.scala 148:37:@42132.4]
  wire  _T_770; // @[SRAM.scala 148:25:@42133.4]
  wire  _T_771; // @[SRAM.scala 148:15:@42134.4]
  wire  _T_772; // @[SRAM.scala 149:15:@42136.6]
  wire  _GEN_9; // @[SRAM.scala 148:48:@42135.4]
  reg  regs_10; // @[SRAM.scala 145:20:@42142.4]
  reg [31:0] _RAND_10;
  wire  _T_778; // @[SRAM.scala 148:37:@42143.4]
  wire  _T_779; // @[SRAM.scala 148:25:@42144.4]
  wire  _T_780; // @[SRAM.scala 148:15:@42145.4]
  wire  _T_781; // @[SRAM.scala 149:15:@42147.6]
  wire  _GEN_10; // @[SRAM.scala 148:48:@42146.4]
  reg  regs_11; // @[SRAM.scala 145:20:@42153.4]
  reg [31:0] _RAND_11;
  wire  _T_787; // @[SRAM.scala 148:37:@42154.4]
  wire  _T_788; // @[SRAM.scala 148:25:@42155.4]
  wire  _T_789; // @[SRAM.scala 148:15:@42156.4]
  wire  _T_790; // @[SRAM.scala 149:15:@42158.6]
  wire  _GEN_11; // @[SRAM.scala 148:48:@42157.4]
  reg  regs_12; // @[SRAM.scala 145:20:@42164.4]
  reg [31:0] _RAND_12;
  wire  _T_796; // @[SRAM.scala 148:37:@42165.4]
  wire  _T_797; // @[SRAM.scala 148:25:@42166.4]
  wire  _T_798; // @[SRAM.scala 148:15:@42167.4]
  wire  _T_799; // @[SRAM.scala 149:15:@42169.6]
  wire  _GEN_12; // @[SRAM.scala 148:48:@42168.4]
  reg  regs_13; // @[SRAM.scala 145:20:@42175.4]
  reg [31:0] _RAND_13;
  wire  _T_805; // @[SRAM.scala 148:37:@42176.4]
  wire  _T_806; // @[SRAM.scala 148:25:@42177.4]
  wire  _T_807; // @[SRAM.scala 148:15:@42178.4]
  wire  _T_808; // @[SRAM.scala 149:15:@42180.6]
  wire  _GEN_13; // @[SRAM.scala 148:48:@42179.4]
  reg  regs_14; // @[SRAM.scala 145:20:@42186.4]
  reg [31:0] _RAND_14;
  wire  _T_814; // @[SRAM.scala 148:37:@42187.4]
  wire  _T_815; // @[SRAM.scala 148:25:@42188.4]
  wire  _T_816; // @[SRAM.scala 148:15:@42189.4]
  wire  _T_817; // @[SRAM.scala 149:15:@42191.6]
  wire  _GEN_14; // @[SRAM.scala 148:48:@42190.4]
  reg  regs_15; // @[SRAM.scala 145:20:@42197.4]
  reg [31:0] _RAND_15;
  wire  _T_823; // @[SRAM.scala 148:37:@42198.4]
  wire  _T_824; // @[SRAM.scala 148:25:@42199.4]
  wire  _T_825; // @[SRAM.scala 148:15:@42200.4]
  wire  _T_826; // @[SRAM.scala 149:15:@42202.6]
  wire  _GEN_15; // @[SRAM.scala 148:48:@42201.4]
  reg  regs_16; // @[SRAM.scala 145:20:@42208.4]
  reg [31:0] _RAND_16;
  wire  _T_832; // @[SRAM.scala 148:37:@42209.4]
  wire  _T_833; // @[SRAM.scala 148:25:@42210.4]
  wire  _T_834; // @[SRAM.scala 148:15:@42211.4]
  wire  _T_835; // @[SRAM.scala 149:15:@42213.6]
  wire  _GEN_16; // @[SRAM.scala 148:48:@42212.4]
  reg  regs_17; // @[SRAM.scala 145:20:@42219.4]
  reg [31:0] _RAND_17;
  wire  _T_841; // @[SRAM.scala 148:37:@42220.4]
  wire  _T_842; // @[SRAM.scala 148:25:@42221.4]
  wire  _T_843; // @[SRAM.scala 148:15:@42222.4]
  wire  _T_844; // @[SRAM.scala 149:15:@42224.6]
  wire  _GEN_17; // @[SRAM.scala 148:48:@42223.4]
  reg  regs_18; // @[SRAM.scala 145:20:@42230.4]
  reg [31:0] _RAND_18;
  wire  _T_850; // @[SRAM.scala 148:37:@42231.4]
  wire  _T_851; // @[SRAM.scala 148:25:@42232.4]
  wire  _T_852; // @[SRAM.scala 148:15:@42233.4]
  wire  _T_853; // @[SRAM.scala 149:15:@42235.6]
  wire  _GEN_18; // @[SRAM.scala 148:48:@42234.4]
  reg  regs_19; // @[SRAM.scala 145:20:@42241.4]
  reg [31:0] _RAND_19;
  wire  _T_859; // @[SRAM.scala 148:37:@42242.4]
  wire  _T_860; // @[SRAM.scala 148:25:@42243.4]
  wire  _T_861; // @[SRAM.scala 148:15:@42244.4]
  wire  _T_862; // @[SRAM.scala 149:15:@42246.6]
  wire  _GEN_19; // @[SRAM.scala 148:48:@42245.4]
  reg  regs_20; // @[SRAM.scala 145:20:@42252.4]
  reg [31:0] _RAND_20;
  wire  _T_868; // @[SRAM.scala 148:37:@42253.4]
  wire  _T_869; // @[SRAM.scala 148:25:@42254.4]
  wire  _T_870; // @[SRAM.scala 148:15:@42255.4]
  wire  _T_871; // @[SRAM.scala 149:15:@42257.6]
  wire  _GEN_20; // @[SRAM.scala 148:48:@42256.4]
  reg  regs_21; // @[SRAM.scala 145:20:@42263.4]
  reg [31:0] _RAND_21;
  wire  _T_877; // @[SRAM.scala 148:37:@42264.4]
  wire  _T_878; // @[SRAM.scala 148:25:@42265.4]
  wire  _T_879; // @[SRAM.scala 148:15:@42266.4]
  wire  _T_880; // @[SRAM.scala 149:15:@42268.6]
  wire  _GEN_21; // @[SRAM.scala 148:48:@42267.4]
  reg  regs_22; // @[SRAM.scala 145:20:@42274.4]
  reg [31:0] _RAND_22;
  wire  _T_886; // @[SRAM.scala 148:37:@42275.4]
  wire  _T_887; // @[SRAM.scala 148:25:@42276.4]
  wire  _T_888; // @[SRAM.scala 148:15:@42277.4]
  wire  _T_889; // @[SRAM.scala 149:15:@42279.6]
  wire  _GEN_22; // @[SRAM.scala 148:48:@42278.4]
  reg  regs_23; // @[SRAM.scala 145:20:@42285.4]
  reg [31:0] _RAND_23;
  wire  _T_895; // @[SRAM.scala 148:37:@42286.4]
  wire  _T_896; // @[SRAM.scala 148:25:@42287.4]
  wire  _T_897; // @[SRAM.scala 148:15:@42288.4]
  wire  _T_898; // @[SRAM.scala 149:15:@42290.6]
  wire  _GEN_23; // @[SRAM.scala 148:48:@42289.4]
  reg  regs_24; // @[SRAM.scala 145:20:@42296.4]
  reg [31:0] _RAND_24;
  wire  _T_904; // @[SRAM.scala 148:37:@42297.4]
  wire  _T_905; // @[SRAM.scala 148:25:@42298.4]
  wire  _T_906; // @[SRAM.scala 148:15:@42299.4]
  wire  _T_907; // @[SRAM.scala 149:15:@42301.6]
  wire  _GEN_24; // @[SRAM.scala 148:48:@42300.4]
  reg  regs_25; // @[SRAM.scala 145:20:@42307.4]
  reg [31:0] _RAND_25;
  wire  _T_913; // @[SRAM.scala 148:37:@42308.4]
  wire  _T_914; // @[SRAM.scala 148:25:@42309.4]
  wire  _T_915; // @[SRAM.scala 148:15:@42310.4]
  wire  _T_916; // @[SRAM.scala 149:15:@42312.6]
  wire  _GEN_25; // @[SRAM.scala 148:48:@42311.4]
  reg  regs_26; // @[SRAM.scala 145:20:@42318.4]
  reg [31:0] _RAND_26;
  wire  _T_922; // @[SRAM.scala 148:37:@42319.4]
  wire  _T_923; // @[SRAM.scala 148:25:@42320.4]
  wire  _T_924; // @[SRAM.scala 148:15:@42321.4]
  wire  _T_925; // @[SRAM.scala 149:15:@42323.6]
  wire  _GEN_26; // @[SRAM.scala 148:48:@42322.4]
  reg  regs_27; // @[SRAM.scala 145:20:@42329.4]
  reg [31:0] _RAND_27;
  wire  _T_931; // @[SRAM.scala 148:37:@42330.4]
  wire  _T_932; // @[SRAM.scala 148:25:@42331.4]
  wire  _T_933; // @[SRAM.scala 148:15:@42332.4]
  wire  _T_934; // @[SRAM.scala 149:15:@42334.6]
  wire  _GEN_27; // @[SRAM.scala 148:48:@42333.4]
  reg  regs_28; // @[SRAM.scala 145:20:@42340.4]
  reg [31:0] _RAND_28;
  wire  _T_940; // @[SRAM.scala 148:37:@42341.4]
  wire  _T_941; // @[SRAM.scala 148:25:@42342.4]
  wire  _T_942; // @[SRAM.scala 148:15:@42343.4]
  wire  _T_943; // @[SRAM.scala 149:15:@42345.6]
  wire  _GEN_28; // @[SRAM.scala 148:48:@42344.4]
  reg  regs_29; // @[SRAM.scala 145:20:@42351.4]
  reg [31:0] _RAND_29;
  wire  _T_949; // @[SRAM.scala 148:37:@42352.4]
  wire  _T_950; // @[SRAM.scala 148:25:@42353.4]
  wire  _T_951; // @[SRAM.scala 148:15:@42354.4]
  wire  _T_952; // @[SRAM.scala 149:15:@42356.6]
  wire  _GEN_29; // @[SRAM.scala 148:48:@42355.4]
  reg  regs_30; // @[SRAM.scala 145:20:@42362.4]
  reg [31:0] _RAND_30;
  wire  _T_958; // @[SRAM.scala 148:37:@42363.4]
  wire  _T_959; // @[SRAM.scala 148:25:@42364.4]
  wire  _T_960; // @[SRAM.scala 148:15:@42365.4]
  wire  _T_961; // @[SRAM.scala 149:15:@42367.6]
  wire  _GEN_30; // @[SRAM.scala 148:48:@42366.4]
  reg  regs_31; // @[SRAM.scala 145:20:@42373.4]
  reg [31:0] _RAND_31;
  wire  _T_967; // @[SRAM.scala 148:37:@42374.4]
  wire  _T_968; // @[SRAM.scala 148:25:@42375.4]
  wire  _T_969; // @[SRAM.scala 148:15:@42376.4]
  wire  _T_970; // @[SRAM.scala 149:15:@42378.6]
  wire  _GEN_31; // @[SRAM.scala 148:48:@42377.4]
  reg  regs_32; // @[SRAM.scala 145:20:@42384.4]
  reg [31:0] _RAND_32;
  wire  _T_976; // @[SRAM.scala 148:37:@42385.4]
  wire  _T_977; // @[SRAM.scala 148:25:@42386.4]
  wire  _T_978; // @[SRAM.scala 148:15:@42387.4]
  wire  _T_979; // @[SRAM.scala 149:15:@42389.6]
  wire  _GEN_32; // @[SRAM.scala 148:48:@42388.4]
  reg  regs_33; // @[SRAM.scala 145:20:@42395.4]
  reg [31:0] _RAND_33;
  wire  _T_985; // @[SRAM.scala 148:37:@42396.4]
  wire  _T_986; // @[SRAM.scala 148:25:@42397.4]
  wire  _T_987; // @[SRAM.scala 148:15:@42398.4]
  wire  _T_988; // @[SRAM.scala 149:15:@42400.6]
  wire  _GEN_33; // @[SRAM.scala 148:48:@42399.4]
  reg  regs_34; // @[SRAM.scala 145:20:@42406.4]
  reg [31:0] _RAND_34;
  wire  _T_994; // @[SRAM.scala 148:37:@42407.4]
  wire  _T_995; // @[SRAM.scala 148:25:@42408.4]
  wire  _T_996; // @[SRAM.scala 148:15:@42409.4]
  wire  _T_997; // @[SRAM.scala 149:15:@42411.6]
  wire  _GEN_34; // @[SRAM.scala 148:48:@42410.4]
  reg  regs_35; // @[SRAM.scala 145:20:@42417.4]
  reg [31:0] _RAND_35;
  wire  _T_1003; // @[SRAM.scala 148:37:@42418.4]
  wire  _T_1004; // @[SRAM.scala 148:25:@42419.4]
  wire  _T_1005; // @[SRAM.scala 148:15:@42420.4]
  wire  _T_1006; // @[SRAM.scala 149:15:@42422.6]
  wire  _GEN_35; // @[SRAM.scala 148:48:@42421.4]
  reg  regs_36; // @[SRAM.scala 145:20:@42428.4]
  reg [31:0] _RAND_36;
  wire  _T_1012; // @[SRAM.scala 148:37:@42429.4]
  wire  _T_1013; // @[SRAM.scala 148:25:@42430.4]
  wire  _T_1014; // @[SRAM.scala 148:15:@42431.4]
  wire  _T_1015; // @[SRAM.scala 149:15:@42433.6]
  wire  _GEN_36; // @[SRAM.scala 148:48:@42432.4]
  reg  regs_37; // @[SRAM.scala 145:20:@42439.4]
  reg [31:0] _RAND_37;
  wire  _T_1021; // @[SRAM.scala 148:37:@42440.4]
  wire  _T_1022; // @[SRAM.scala 148:25:@42441.4]
  wire  _T_1023; // @[SRAM.scala 148:15:@42442.4]
  wire  _T_1024; // @[SRAM.scala 149:15:@42444.6]
  wire  _GEN_37; // @[SRAM.scala 148:48:@42443.4]
  reg  regs_38; // @[SRAM.scala 145:20:@42450.4]
  reg [31:0] _RAND_38;
  wire  _T_1030; // @[SRAM.scala 148:37:@42451.4]
  wire  _T_1031; // @[SRAM.scala 148:25:@42452.4]
  wire  _T_1032; // @[SRAM.scala 148:15:@42453.4]
  wire  _T_1033; // @[SRAM.scala 149:15:@42455.6]
  wire  _GEN_38; // @[SRAM.scala 148:48:@42454.4]
  reg  regs_39; // @[SRAM.scala 145:20:@42461.4]
  reg [31:0] _RAND_39;
  wire  _T_1039; // @[SRAM.scala 148:37:@42462.4]
  wire  _T_1040; // @[SRAM.scala 148:25:@42463.4]
  wire  _T_1041; // @[SRAM.scala 148:15:@42464.4]
  wire  _T_1042; // @[SRAM.scala 149:15:@42466.6]
  wire  _GEN_39; // @[SRAM.scala 148:48:@42465.4]
  reg  regs_40; // @[SRAM.scala 145:20:@42472.4]
  reg [31:0] _RAND_40;
  wire  _T_1048; // @[SRAM.scala 148:37:@42473.4]
  wire  _T_1049; // @[SRAM.scala 148:25:@42474.4]
  wire  _T_1050; // @[SRAM.scala 148:15:@42475.4]
  wire  _T_1051; // @[SRAM.scala 149:15:@42477.6]
  wire  _GEN_40; // @[SRAM.scala 148:48:@42476.4]
  reg  regs_41; // @[SRAM.scala 145:20:@42483.4]
  reg [31:0] _RAND_41;
  wire  _T_1057; // @[SRAM.scala 148:37:@42484.4]
  wire  _T_1058; // @[SRAM.scala 148:25:@42485.4]
  wire  _T_1059; // @[SRAM.scala 148:15:@42486.4]
  wire  _T_1060; // @[SRAM.scala 149:15:@42488.6]
  wire  _GEN_41; // @[SRAM.scala 148:48:@42487.4]
  reg  regs_42; // @[SRAM.scala 145:20:@42494.4]
  reg [31:0] _RAND_42;
  wire  _T_1066; // @[SRAM.scala 148:37:@42495.4]
  wire  _T_1067; // @[SRAM.scala 148:25:@42496.4]
  wire  _T_1068; // @[SRAM.scala 148:15:@42497.4]
  wire  _T_1069; // @[SRAM.scala 149:15:@42499.6]
  wire  _GEN_42; // @[SRAM.scala 148:48:@42498.4]
  reg  regs_43; // @[SRAM.scala 145:20:@42505.4]
  reg [31:0] _RAND_43;
  wire  _T_1075; // @[SRAM.scala 148:37:@42506.4]
  wire  _T_1076; // @[SRAM.scala 148:25:@42507.4]
  wire  _T_1077; // @[SRAM.scala 148:15:@42508.4]
  wire  _T_1078; // @[SRAM.scala 149:15:@42510.6]
  wire  _GEN_43; // @[SRAM.scala 148:48:@42509.4]
  reg  regs_44; // @[SRAM.scala 145:20:@42516.4]
  reg [31:0] _RAND_44;
  wire  _T_1084; // @[SRAM.scala 148:37:@42517.4]
  wire  _T_1085; // @[SRAM.scala 148:25:@42518.4]
  wire  _T_1086; // @[SRAM.scala 148:15:@42519.4]
  wire  _T_1087; // @[SRAM.scala 149:15:@42521.6]
  wire  _GEN_44; // @[SRAM.scala 148:48:@42520.4]
  reg  regs_45; // @[SRAM.scala 145:20:@42527.4]
  reg [31:0] _RAND_45;
  wire  _T_1093; // @[SRAM.scala 148:37:@42528.4]
  wire  _T_1094; // @[SRAM.scala 148:25:@42529.4]
  wire  _T_1095; // @[SRAM.scala 148:15:@42530.4]
  wire  _T_1096; // @[SRAM.scala 149:15:@42532.6]
  wire  _GEN_45; // @[SRAM.scala 148:48:@42531.4]
  reg  regs_46; // @[SRAM.scala 145:20:@42538.4]
  reg [31:0] _RAND_46;
  wire  _T_1102; // @[SRAM.scala 148:37:@42539.4]
  wire  _T_1103; // @[SRAM.scala 148:25:@42540.4]
  wire  _T_1104; // @[SRAM.scala 148:15:@42541.4]
  wire  _T_1105; // @[SRAM.scala 149:15:@42543.6]
  wire  _GEN_46; // @[SRAM.scala 148:48:@42542.4]
  reg  regs_47; // @[SRAM.scala 145:20:@42549.4]
  reg [31:0] _RAND_47;
  wire  _T_1111; // @[SRAM.scala 148:37:@42550.4]
  wire  _T_1112; // @[SRAM.scala 148:25:@42551.4]
  wire  _T_1113; // @[SRAM.scala 148:15:@42552.4]
  wire  _T_1114; // @[SRAM.scala 149:15:@42554.6]
  wire  _GEN_47; // @[SRAM.scala 148:48:@42553.4]
  reg  regs_48; // @[SRAM.scala 145:20:@42560.4]
  reg [31:0] _RAND_48;
  wire  _T_1120; // @[SRAM.scala 148:37:@42561.4]
  wire  _T_1121; // @[SRAM.scala 148:25:@42562.4]
  wire  _T_1122; // @[SRAM.scala 148:15:@42563.4]
  wire  _T_1123; // @[SRAM.scala 149:15:@42565.6]
  wire  _GEN_48; // @[SRAM.scala 148:48:@42564.4]
  reg  regs_49; // @[SRAM.scala 145:20:@42571.4]
  reg [31:0] _RAND_49;
  wire  _T_1129; // @[SRAM.scala 148:37:@42572.4]
  wire  _T_1130; // @[SRAM.scala 148:25:@42573.4]
  wire  _T_1131; // @[SRAM.scala 148:15:@42574.4]
  wire  _T_1132; // @[SRAM.scala 149:15:@42576.6]
  wire  _GEN_49; // @[SRAM.scala 148:48:@42575.4]
  reg  regs_50; // @[SRAM.scala 145:20:@42582.4]
  reg [31:0] _RAND_50;
  wire  _T_1138; // @[SRAM.scala 148:37:@42583.4]
  wire  _T_1139; // @[SRAM.scala 148:25:@42584.4]
  wire  _T_1140; // @[SRAM.scala 148:15:@42585.4]
  wire  _T_1141; // @[SRAM.scala 149:15:@42587.6]
  wire  _GEN_50; // @[SRAM.scala 148:48:@42586.4]
  reg  regs_51; // @[SRAM.scala 145:20:@42593.4]
  reg [31:0] _RAND_51;
  wire  _T_1147; // @[SRAM.scala 148:37:@42594.4]
  wire  _T_1148; // @[SRAM.scala 148:25:@42595.4]
  wire  _T_1149; // @[SRAM.scala 148:15:@42596.4]
  wire  _T_1150; // @[SRAM.scala 149:15:@42598.6]
  wire  _GEN_51; // @[SRAM.scala 148:48:@42597.4]
  reg  regs_52; // @[SRAM.scala 145:20:@42604.4]
  reg [31:0] _RAND_52;
  wire  _T_1156; // @[SRAM.scala 148:37:@42605.4]
  wire  _T_1157; // @[SRAM.scala 148:25:@42606.4]
  wire  _T_1158; // @[SRAM.scala 148:15:@42607.4]
  wire  _T_1159; // @[SRAM.scala 149:15:@42609.6]
  wire  _GEN_52; // @[SRAM.scala 148:48:@42608.4]
  reg  regs_53; // @[SRAM.scala 145:20:@42615.4]
  reg [31:0] _RAND_53;
  wire  _T_1165; // @[SRAM.scala 148:37:@42616.4]
  wire  _T_1166; // @[SRAM.scala 148:25:@42617.4]
  wire  _T_1167; // @[SRAM.scala 148:15:@42618.4]
  wire  _T_1168; // @[SRAM.scala 149:15:@42620.6]
  wire  _GEN_53; // @[SRAM.scala 148:48:@42619.4]
  reg  regs_54; // @[SRAM.scala 145:20:@42626.4]
  reg [31:0] _RAND_54;
  wire  _T_1174; // @[SRAM.scala 148:37:@42627.4]
  wire  _T_1175; // @[SRAM.scala 148:25:@42628.4]
  wire  _T_1176; // @[SRAM.scala 148:15:@42629.4]
  wire  _T_1177; // @[SRAM.scala 149:15:@42631.6]
  wire  _GEN_54; // @[SRAM.scala 148:48:@42630.4]
  reg  regs_55; // @[SRAM.scala 145:20:@42637.4]
  reg [31:0] _RAND_55;
  wire  _T_1183; // @[SRAM.scala 148:37:@42638.4]
  wire  _T_1184; // @[SRAM.scala 148:25:@42639.4]
  wire  _T_1185; // @[SRAM.scala 148:15:@42640.4]
  wire  _T_1186; // @[SRAM.scala 149:15:@42642.6]
  wire  _GEN_55; // @[SRAM.scala 148:48:@42641.4]
  reg  regs_56; // @[SRAM.scala 145:20:@42648.4]
  reg [31:0] _RAND_56;
  wire  _T_1192; // @[SRAM.scala 148:37:@42649.4]
  wire  _T_1193; // @[SRAM.scala 148:25:@42650.4]
  wire  _T_1194; // @[SRAM.scala 148:15:@42651.4]
  wire  _T_1195; // @[SRAM.scala 149:15:@42653.6]
  wire  _GEN_56; // @[SRAM.scala 148:48:@42652.4]
  reg  regs_57; // @[SRAM.scala 145:20:@42659.4]
  reg [31:0] _RAND_57;
  wire  _T_1201; // @[SRAM.scala 148:37:@42660.4]
  wire  _T_1202; // @[SRAM.scala 148:25:@42661.4]
  wire  _T_1203; // @[SRAM.scala 148:15:@42662.4]
  wire  _T_1204; // @[SRAM.scala 149:15:@42664.6]
  wire  _GEN_57; // @[SRAM.scala 148:48:@42663.4]
  reg  regs_58; // @[SRAM.scala 145:20:@42670.4]
  reg [31:0] _RAND_58;
  wire  _T_1210; // @[SRAM.scala 148:37:@42671.4]
  wire  _T_1211; // @[SRAM.scala 148:25:@42672.4]
  wire  _T_1212; // @[SRAM.scala 148:15:@42673.4]
  wire  _T_1213; // @[SRAM.scala 149:15:@42675.6]
  wire  _GEN_58; // @[SRAM.scala 148:48:@42674.4]
  reg  regs_59; // @[SRAM.scala 145:20:@42681.4]
  reg [31:0] _RAND_59;
  wire  _T_1219; // @[SRAM.scala 148:37:@42682.4]
  wire  _T_1220; // @[SRAM.scala 148:25:@42683.4]
  wire  _T_1221; // @[SRAM.scala 148:15:@42684.4]
  wire  _T_1222; // @[SRAM.scala 149:15:@42686.6]
  wire  _GEN_59; // @[SRAM.scala 148:48:@42685.4]
  reg  regs_60; // @[SRAM.scala 145:20:@42692.4]
  reg [31:0] _RAND_60;
  wire  _T_1228; // @[SRAM.scala 148:37:@42693.4]
  wire  _T_1229; // @[SRAM.scala 148:25:@42694.4]
  wire  _T_1230; // @[SRAM.scala 148:15:@42695.4]
  wire  _T_1231; // @[SRAM.scala 149:15:@42697.6]
  wire  _GEN_60; // @[SRAM.scala 148:48:@42696.4]
  reg  regs_61; // @[SRAM.scala 145:20:@42703.4]
  reg [31:0] _RAND_61;
  wire  _T_1237; // @[SRAM.scala 148:37:@42704.4]
  wire  _T_1238; // @[SRAM.scala 148:25:@42705.4]
  wire  _T_1239; // @[SRAM.scala 148:15:@42706.4]
  wire  _T_1240; // @[SRAM.scala 149:15:@42708.6]
  wire  _GEN_61; // @[SRAM.scala 148:48:@42707.4]
  reg  regs_62; // @[SRAM.scala 145:20:@42714.4]
  reg [31:0] _RAND_62;
  wire  _T_1246; // @[SRAM.scala 148:37:@42715.4]
  wire  _T_1247; // @[SRAM.scala 148:25:@42716.4]
  wire  _T_1248; // @[SRAM.scala 148:15:@42717.4]
  wire  _T_1249; // @[SRAM.scala 149:15:@42719.6]
  wire  _GEN_62; // @[SRAM.scala 148:48:@42718.4]
  reg  regs_63; // @[SRAM.scala 145:20:@42725.4]
  reg [31:0] _RAND_63;
  wire  _T_1255; // @[SRAM.scala 148:37:@42726.4]
  wire  _T_1256; // @[SRAM.scala 148:25:@42727.4]
  wire  _T_1257; // @[SRAM.scala 148:15:@42728.4]
  wire  _T_1258; // @[SRAM.scala 149:15:@42730.6]
  wire  _GEN_63; // @[SRAM.scala 148:48:@42729.4]
  wire  _GEN_65; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_66; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_67; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_68; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_69; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_70; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_71; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_72; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_73; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_74; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_75; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_76; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_77; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_78; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_79; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_80; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_81; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_82; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_83; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_84; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_85; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_86; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_87; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_88; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_89; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_90; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_91; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_92; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_93; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_94; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_95; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_96; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_97; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_98; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_99; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_100; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_101; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_102; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_103; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_104; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_105; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_106; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_107; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_108; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_109; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_110; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_111; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_112; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_113; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_114; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_115; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_116; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_117; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_118; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_119; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_120; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_121; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_122; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_123; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_124; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_125; // @[SRAM.scala 155:12:@42799.4]
  wire  _GEN_126; // @[SRAM.scala 155:12:@42799.4]
  assign _T_688 = io_waddr == 6'h0; // @[SRAM.scala 148:37:@42033.4]
  assign _T_689 = io_wen & _T_688; // @[SRAM.scala 148:25:@42034.4]
  assign _T_690 = io_banks_0_wdata_valid | _T_689; // @[SRAM.scala 148:15:@42035.4]
  assign _T_691 = io_banks_0_wdata_valid ? io_banks_0_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42037.6]
  assign _GEN_0 = _T_690 ? _T_691 : regs_0; // @[SRAM.scala 148:48:@42036.4]
  assign _T_697 = io_waddr == 6'h1; // @[SRAM.scala 148:37:@42044.4]
  assign _T_698 = io_wen & _T_697; // @[SRAM.scala 148:25:@42045.4]
  assign _T_699 = io_banks_1_wdata_valid | _T_698; // @[SRAM.scala 148:15:@42046.4]
  assign _T_700 = io_banks_1_wdata_valid ? io_banks_1_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42048.6]
  assign _GEN_1 = _T_699 ? _T_700 : regs_1; // @[SRAM.scala 148:48:@42047.4]
  assign _T_706 = io_waddr == 6'h2; // @[SRAM.scala 148:37:@42055.4]
  assign _T_707 = io_wen & _T_706; // @[SRAM.scala 148:25:@42056.4]
  assign _T_708 = io_banks_2_wdata_valid | _T_707; // @[SRAM.scala 148:15:@42057.4]
  assign _T_709 = io_banks_2_wdata_valid ? io_banks_2_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42059.6]
  assign _GEN_2 = _T_708 ? _T_709 : regs_2; // @[SRAM.scala 148:48:@42058.4]
  assign _T_715 = io_waddr == 6'h3; // @[SRAM.scala 148:37:@42066.4]
  assign _T_716 = io_wen & _T_715; // @[SRAM.scala 148:25:@42067.4]
  assign _T_717 = io_banks_3_wdata_valid | _T_716; // @[SRAM.scala 148:15:@42068.4]
  assign _T_718 = io_banks_3_wdata_valid ? io_banks_3_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42070.6]
  assign _GEN_3 = _T_717 ? _T_718 : regs_3; // @[SRAM.scala 148:48:@42069.4]
  assign _T_724 = io_waddr == 6'h4; // @[SRAM.scala 148:37:@42077.4]
  assign _T_725 = io_wen & _T_724; // @[SRAM.scala 148:25:@42078.4]
  assign _T_726 = io_banks_4_wdata_valid | _T_725; // @[SRAM.scala 148:15:@42079.4]
  assign _T_727 = io_banks_4_wdata_valid ? io_banks_4_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42081.6]
  assign _GEN_4 = _T_726 ? _T_727 : regs_4; // @[SRAM.scala 148:48:@42080.4]
  assign _T_733 = io_waddr == 6'h5; // @[SRAM.scala 148:37:@42088.4]
  assign _T_734 = io_wen & _T_733; // @[SRAM.scala 148:25:@42089.4]
  assign _T_735 = io_banks_5_wdata_valid | _T_734; // @[SRAM.scala 148:15:@42090.4]
  assign _T_736 = io_banks_5_wdata_valid ? io_banks_5_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42092.6]
  assign _GEN_5 = _T_735 ? _T_736 : regs_5; // @[SRAM.scala 148:48:@42091.4]
  assign _T_742 = io_waddr == 6'h6; // @[SRAM.scala 148:37:@42099.4]
  assign _T_743 = io_wen & _T_742; // @[SRAM.scala 148:25:@42100.4]
  assign _T_744 = io_banks_6_wdata_valid | _T_743; // @[SRAM.scala 148:15:@42101.4]
  assign _T_745 = io_banks_6_wdata_valid ? io_banks_6_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42103.6]
  assign _GEN_6 = _T_744 ? _T_745 : regs_6; // @[SRAM.scala 148:48:@42102.4]
  assign _T_751 = io_waddr == 6'h7; // @[SRAM.scala 148:37:@42110.4]
  assign _T_752 = io_wen & _T_751; // @[SRAM.scala 148:25:@42111.4]
  assign _T_753 = io_banks_7_wdata_valid | _T_752; // @[SRAM.scala 148:15:@42112.4]
  assign _T_754 = io_banks_7_wdata_valid ? io_banks_7_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42114.6]
  assign _GEN_7 = _T_753 ? _T_754 : regs_7; // @[SRAM.scala 148:48:@42113.4]
  assign _T_760 = io_waddr == 6'h8; // @[SRAM.scala 148:37:@42121.4]
  assign _T_761 = io_wen & _T_760; // @[SRAM.scala 148:25:@42122.4]
  assign _T_762 = io_banks_8_wdata_valid | _T_761; // @[SRAM.scala 148:15:@42123.4]
  assign _T_763 = io_banks_8_wdata_valid ? io_banks_8_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42125.6]
  assign _GEN_8 = _T_762 ? _T_763 : regs_8; // @[SRAM.scala 148:48:@42124.4]
  assign _T_769 = io_waddr == 6'h9; // @[SRAM.scala 148:37:@42132.4]
  assign _T_770 = io_wen & _T_769; // @[SRAM.scala 148:25:@42133.4]
  assign _T_771 = io_banks_9_wdata_valid | _T_770; // @[SRAM.scala 148:15:@42134.4]
  assign _T_772 = io_banks_9_wdata_valid ? io_banks_9_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42136.6]
  assign _GEN_9 = _T_771 ? _T_772 : regs_9; // @[SRAM.scala 148:48:@42135.4]
  assign _T_778 = io_waddr == 6'ha; // @[SRAM.scala 148:37:@42143.4]
  assign _T_779 = io_wen & _T_778; // @[SRAM.scala 148:25:@42144.4]
  assign _T_780 = io_banks_10_wdata_valid | _T_779; // @[SRAM.scala 148:15:@42145.4]
  assign _T_781 = io_banks_10_wdata_valid ? io_banks_10_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42147.6]
  assign _GEN_10 = _T_780 ? _T_781 : regs_10; // @[SRAM.scala 148:48:@42146.4]
  assign _T_787 = io_waddr == 6'hb; // @[SRAM.scala 148:37:@42154.4]
  assign _T_788 = io_wen & _T_787; // @[SRAM.scala 148:25:@42155.4]
  assign _T_789 = io_banks_11_wdata_valid | _T_788; // @[SRAM.scala 148:15:@42156.4]
  assign _T_790 = io_banks_11_wdata_valid ? io_banks_11_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42158.6]
  assign _GEN_11 = _T_789 ? _T_790 : regs_11; // @[SRAM.scala 148:48:@42157.4]
  assign _T_796 = io_waddr == 6'hc; // @[SRAM.scala 148:37:@42165.4]
  assign _T_797 = io_wen & _T_796; // @[SRAM.scala 148:25:@42166.4]
  assign _T_798 = io_banks_12_wdata_valid | _T_797; // @[SRAM.scala 148:15:@42167.4]
  assign _T_799 = io_banks_12_wdata_valid ? io_banks_12_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42169.6]
  assign _GEN_12 = _T_798 ? _T_799 : regs_12; // @[SRAM.scala 148:48:@42168.4]
  assign _T_805 = io_waddr == 6'hd; // @[SRAM.scala 148:37:@42176.4]
  assign _T_806 = io_wen & _T_805; // @[SRAM.scala 148:25:@42177.4]
  assign _T_807 = io_banks_13_wdata_valid | _T_806; // @[SRAM.scala 148:15:@42178.4]
  assign _T_808 = io_banks_13_wdata_valid ? io_banks_13_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42180.6]
  assign _GEN_13 = _T_807 ? _T_808 : regs_13; // @[SRAM.scala 148:48:@42179.4]
  assign _T_814 = io_waddr == 6'he; // @[SRAM.scala 148:37:@42187.4]
  assign _T_815 = io_wen & _T_814; // @[SRAM.scala 148:25:@42188.4]
  assign _T_816 = io_banks_14_wdata_valid | _T_815; // @[SRAM.scala 148:15:@42189.4]
  assign _T_817 = io_banks_14_wdata_valid ? io_banks_14_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42191.6]
  assign _GEN_14 = _T_816 ? _T_817 : regs_14; // @[SRAM.scala 148:48:@42190.4]
  assign _T_823 = io_waddr == 6'hf; // @[SRAM.scala 148:37:@42198.4]
  assign _T_824 = io_wen & _T_823; // @[SRAM.scala 148:25:@42199.4]
  assign _T_825 = io_banks_15_wdata_valid | _T_824; // @[SRAM.scala 148:15:@42200.4]
  assign _T_826 = io_banks_15_wdata_valid ? io_banks_15_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42202.6]
  assign _GEN_15 = _T_825 ? _T_826 : regs_15; // @[SRAM.scala 148:48:@42201.4]
  assign _T_832 = io_waddr == 6'h10; // @[SRAM.scala 148:37:@42209.4]
  assign _T_833 = io_wen & _T_832; // @[SRAM.scala 148:25:@42210.4]
  assign _T_834 = io_banks_16_wdata_valid | _T_833; // @[SRAM.scala 148:15:@42211.4]
  assign _T_835 = io_banks_16_wdata_valid ? io_banks_16_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42213.6]
  assign _GEN_16 = _T_834 ? _T_835 : regs_16; // @[SRAM.scala 148:48:@42212.4]
  assign _T_841 = io_waddr == 6'h11; // @[SRAM.scala 148:37:@42220.4]
  assign _T_842 = io_wen & _T_841; // @[SRAM.scala 148:25:@42221.4]
  assign _T_843 = io_banks_17_wdata_valid | _T_842; // @[SRAM.scala 148:15:@42222.4]
  assign _T_844 = io_banks_17_wdata_valid ? io_banks_17_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42224.6]
  assign _GEN_17 = _T_843 ? _T_844 : regs_17; // @[SRAM.scala 148:48:@42223.4]
  assign _T_850 = io_waddr == 6'h12; // @[SRAM.scala 148:37:@42231.4]
  assign _T_851 = io_wen & _T_850; // @[SRAM.scala 148:25:@42232.4]
  assign _T_852 = io_banks_18_wdata_valid | _T_851; // @[SRAM.scala 148:15:@42233.4]
  assign _T_853 = io_banks_18_wdata_valid ? io_banks_18_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42235.6]
  assign _GEN_18 = _T_852 ? _T_853 : regs_18; // @[SRAM.scala 148:48:@42234.4]
  assign _T_859 = io_waddr == 6'h13; // @[SRAM.scala 148:37:@42242.4]
  assign _T_860 = io_wen & _T_859; // @[SRAM.scala 148:25:@42243.4]
  assign _T_861 = io_banks_19_wdata_valid | _T_860; // @[SRAM.scala 148:15:@42244.4]
  assign _T_862 = io_banks_19_wdata_valid ? io_banks_19_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42246.6]
  assign _GEN_19 = _T_861 ? _T_862 : regs_19; // @[SRAM.scala 148:48:@42245.4]
  assign _T_868 = io_waddr == 6'h14; // @[SRAM.scala 148:37:@42253.4]
  assign _T_869 = io_wen & _T_868; // @[SRAM.scala 148:25:@42254.4]
  assign _T_870 = io_banks_20_wdata_valid | _T_869; // @[SRAM.scala 148:15:@42255.4]
  assign _T_871 = io_banks_20_wdata_valid ? io_banks_20_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42257.6]
  assign _GEN_20 = _T_870 ? _T_871 : regs_20; // @[SRAM.scala 148:48:@42256.4]
  assign _T_877 = io_waddr == 6'h15; // @[SRAM.scala 148:37:@42264.4]
  assign _T_878 = io_wen & _T_877; // @[SRAM.scala 148:25:@42265.4]
  assign _T_879 = io_banks_21_wdata_valid | _T_878; // @[SRAM.scala 148:15:@42266.4]
  assign _T_880 = io_banks_21_wdata_valid ? io_banks_21_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42268.6]
  assign _GEN_21 = _T_879 ? _T_880 : regs_21; // @[SRAM.scala 148:48:@42267.4]
  assign _T_886 = io_waddr == 6'h16; // @[SRAM.scala 148:37:@42275.4]
  assign _T_887 = io_wen & _T_886; // @[SRAM.scala 148:25:@42276.4]
  assign _T_888 = io_banks_22_wdata_valid | _T_887; // @[SRAM.scala 148:15:@42277.4]
  assign _T_889 = io_banks_22_wdata_valid ? io_banks_22_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42279.6]
  assign _GEN_22 = _T_888 ? _T_889 : regs_22; // @[SRAM.scala 148:48:@42278.4]
  assign _T_895 = io_waddr == 6'h17; // @[SRAM.scala 148:37:@42286.4]
  assign _T_896 = io_wen & _T_895; // @[SRAM.scala 148:25:@42287.4]
  assign _T_897 = io_banks_23_wdata_valid | _T_896; // @[SRAM.scala 148:15:@42288.4]
  assign _T_898 = io_banks_23_wdata_valid ? io_banks_23_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42290.6]
  assign _GEN_23 = _T_897 ? _T_898 : regs_23; // @[SRAM.scala 148:48:@42289.4]
  assign _T_904 = io_waddr == 6'h18; // @[SRAM.scala 148:37:@42297.4]
  assign _T_905 = io_wen & _T_904; // @[SRAM.scala 148:25:@42298.4]
  assign _T_906 = io_banks_24_wdata_valid | _T_905; // @[SRAM.scala 148:15:@42299.4]
  assign _T_907 = io_banks_24_wdata_valid ? io_banks_24_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42301.6]
  assign _GEN_24 = _T_906 ? _T_907 : regs_24; // @[SRAM.scala 148:48:@42300.4]
  assign _T_913 = io_waddr == 6'h19; // @[SRAM.scala 148:37:@42308.4]
  assign _T_914 = io_wen & _T_913; // @[SRAM.scala 148:25:@42309.4]
  assign _T_915 = io_banks_25_wdata_valid | _T_914; // @[SRAM.scala 148:15:@42310.4]
  assign _T_916 = io_banks_25_wdata_valid ? io_banks_25_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42312.6]
  assign _GEN_25 = _T_915 ? _T_916 : regs_25; // @[SRAM.scala 148:48:@42311.4]
  assign _T_922 = io_waddr == 6'h1a; // @[SRAM.scala 148:37:@42319.4]
  assign _T_923 = io_wen & _T_922; // @[SRAM.scala 148:25:@42320.4]
  assign _T_924 = io_banks_26_wdata_valid | _T_923; // @[SRAM.scala 148:15:@42321.4]
  assign _T_925 = io_banks_26_wdata_valid ? io_banks_26_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42323.6]
  assign _GEN_26 = _T_924 ? _T_925 : regs_26; // @[SRAM.scala 148:48:@42322.4]
  assign _T_931 = io_waddr == 6'h1b; // @[SRAM.scala 148:37:@42330.4]
  assign _T_932 = io_wen & _T_931; // @[SRAM.scala 148:25:@42331.4]
  assign _T_933 = io_banks_27_wdata_valid | _T_932; // @[SRAM.scala 148:15:@42332.4]
  assign _T_934 = io_banks_27_wdata_valid ? io_banks_27_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42334.6]
  assign _GEN_27 = _T_933 ? _T_934 : regs_27; // @[SRAM.scala 148:48:@42333.4]
  assign _T_940 = io_waddr == 6'h1c; // @[SRAM.scala 148:37:@42341.4]
  assign _T_941 = io_wen & _T_940; // @[SRAM.scala 148:25:@42342.4]
  assign _T_942 = io_banks_28_wdata_valid | _T_941; // @[SRAM.scala 148:15:@42343.4]
  assign _T_943 = io_banks_28_wdata_valid ? io_banks_28_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42345.6]
  assign _GEN_28 = _T_942 ? _T_943 : regs_28; // @[SRAM.scala 148:48:@42344.4]
  assign _T_949 = io_waddr == 6'h1d; // @[SRAM.scala 148:37:@42352.4]
  assign _T_950 = io_wen & _T_949; // @[SRAM.scala 148:25:@42353.4]
  assign _T_951 = io_banks_29_wdata_valid | _T_950; // @[SRAM.scala 148:15:@42354.4]
  assign _T_952 = io_banks_29_wdata_valid ? io_banks_29_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42356.6]
  assign _GEN_29 = _T_951 ? _T_952 : regs_29; // @[SRAM.scala 148:48:@42355.4]
  assign _T_958 = io_waddr == 6'h1e; // @[SRAM.scala 148:37:@42363.4]
  assign _T_959 = io_wen & _T_958; // @[SRAM.scala 148:25:@42364.4]
  assign _T_960 = io_banks_30_wdata_valid | _T_959; // @[SRAM.scala 148:15:@42365.4]
  assign _T_961 = io_banks_30_wdata_valid ? io_banks_30_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42367.6]
  assign _GEN_30 = _T_960 ? _T_961 : regs_30; // @[SRAM.scala 148:48:@42366.4]
  assign _T_967 = io_waddr == 6'h1f; // @[SRAM.scala 148:37:@42374.4]
  assign _T_968 = io_wen & _T_967; // @[SRAM.scala 148:25:@42375.4]
  assign _T_969 = io_banks_31_wdata_valid | _T_968; // @[SRAM.scala 148:15:@42376.4]
  assign _T_970 = io_banks_31_wdata_valid ? io_banks_31_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42378.6]
  assign _GEN_31 = _T_969 ? _T_970 : regs_31; // @[SRAM.scala 148:48:@42377.4]
  assign _T_976 = io_waddr == 6'h20; // @[SRAM.scala 148:37:@42385.4]
  assign _T_977 = io_wen & _T_976; // @[SRAM.scala 148:25:@42386.4]
  assign _T_978 = io_banks_32_wdata_valid | _T_977; // @[SRAM.scala 148:15:@42387.4]
  assign _T_979 = io_banks_32_wdata_valid ? io_banks_32_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42389.6]
  assign _GEN_32 = _T_978 ? _T_979 : regs_32; // @[SRAM.scala 148:48:@42388.4]
  assign _T_985 = io_waddr == 6'h21; // @[SRAM.scala 148:37:@42396.4]
  assign _T_986 = io_wen & _T_985; // @[SRAM.scala 148:25:@42397.4]
  assign _T_987 = io_banks_33_wdata_valid | _T_986; // @[SRAM.scala 148:15:@42398.4]
  assign _T_988 = io_banks_33_wdata_valid ? io_banks_33_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42400.6]
  assign _GEN_33 = _T_987 ? _T_988 : regs_33; // @[SRAM.scala 148:48:@42399.4]
  assign _T_994 = io_waddr == 6'h22; // @[SRAM.scala 148:37:@42407.4]
  assign _T_995 = io_wen & _T_994; // @[SRAM.scala 148:25:@42408.4]
  assign _T_996 = io_banks_34_wdata_valid | _T_995; // @[SRAM.scala 148:15:@42409.4]
  assign _T_997 = io_banks_34_wdata_valid ? io_banks_34_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42411.6]
  assign _GEN_34 = _T_996 ? _T_997 : regs_34; // @[SRAM.scala 148:48:@42410.4]
  assign _T_1003 = io_waddr == 6'h23; // @[SRAM.scala 148:37:@42418.4]
  assign _T_1004 = io_wen & _T_1003; // @[SRAM.scala 148:25:@42419.4]
  assign _T_1005 = io_banks_35_wdata_valid | _T_1004; // @[SRAM.scala 148:15:@42420.4]
  assign _T_1006 = io_banks_35_wdata_valid ? io_banks_35_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42422.6]
  assign _GEN_35 = _T_1005 ? _T_1006 : regs_35; // @[SRAM.scala 148:48:@42421.4]
  assign _T_1012 = io_waddr == 6'h24; // @[SRAM.scala 148:37:@42429.4]
  assign _T_1013 = io_wen & _T_1012; // @[SRAM.scala 148:25:@42430.4]
  assign _T_1014 = io_banks_36_wdata_valid | _T_1013; // @[SRAM.scala 148:15:@42431.4]
  assign _T_1015 = io_banks_36_wdata_valid ? io_banks_36_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42433.6]
  assign _GEN_36 = _T_1014 ? _T_1015 : regs_36; // @[SRAM.scala 148:48:@42432.4]
  assign _T_1021 = io_waddr == 6'h25; // @[SRAM.scala 148:37:@42440.4]
  assign _T_1022 = io_wen & _T_1021; // @[SRAM.scala 148:25:@42441.4]
  assign _T_1023 = io_banks_37_wdata_valid | _T_1022; // @[SRAM.scala 148:15:@42442.4]
  assign _T_1024 = io_banks_37_wdata_valid ? io_banks_37_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42444.6]
  assign _GEN_37 = _T_1023 ? _T_1024 : regs_37; // @[SRAM.scala 148:48:@42443.4]
  assign _T_1030 = io_waddr == 6'h26; // @[SRAM.scala 148:37:@42451.4]
  assign _T_1031 = io_wen & _T_1030; // @[SRAM.scala 148:25:@42452.4]
  assign _T_1032 = io_banks_38_wdata_valid | _T_1031; // @[SRAM.scala 148:15:@42453.4]
  assign _T_1033 = io_banks_38_wdata_valid ? io_banks_38_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42455.6]
  assign _GEN_38 = _T_1032 ? _T_1033 : regs_38; // @[SRAM.scala 148:48:@42454.4]
  assign _T_1039 = io_waddr == 6'h27; // @[SRAM.scala 148:37:@42462.4]
  assign _T_1040 = io_wen & _T_1039; // @[SRAM.scala 148:25:@42463.4]
  assign _T_1041 = io_banks_39_wdata_valid | _T_1040; // @[SRAM.scala 148:15:@42464.4]
  assign _T_1042 = io_banks_39_wdata_valid ? io_banks_39_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42466.6]
  assign _GEN_39 = _T_1041 ? _T_1042 : regs_39; // @[SRAM.scala 148:48:@42465.4]
  assign _T_1048 = io_waddr == 6'h28; // @[SRAM.scala 148:37:@42473.4]
  assign _T_1049 = io_wen & _T_1048; // @[SRAM.scala 148:25:@42474.4]
  assign _T_1050 = io_banks_40_wdata_valid | _T_1049; // @[SRAM.scala 148:15:@42475.4]
  assign _T_1051 = io_banks_40_wdata_valid ? io_banks_40_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42477.6]
  assign _GEN_40 = _T_1050 ? _T_1051 : regs_40; // @[SRAM.scala 148:48:@42476.4]
  assign _T_1057 = io_waddr == 6'h29; // @[SRAM.scala 148:37:@42484.4]
  assign _T_1058 = io_wen & _T_1057; // @[SRAM.scala 148:25:@42485.4]
  assign _T_1059 = io_banks_41_wdata_valid | _T_1058; // @[SRAM.scala 148:15:@42486.4]
  assign _T_1060 = io_banks_41_wdata_valid ? io_banks_41_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42488.6]
  assign _GEN_41 = _T_1059 ? _T_1060 : regs_41; // @[SRAM.scala 148:48:@42487.4]
  assign _T_1066 = io_waddr == 6'h2a; // @[SRAM.scala 148:37:@42495.4]
  assign _T_1067 = io_wen & _T_1066; // @[SRAM.scala 148:25:@42496.4]
  assign _T_1068 = io_banks_42_wdata_valid | _T_1067; // @[SRAM.scala 148:15:@42497.4]
  assign _T_1069 = io_banks_42_wdata_valid ? io_banks_42_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42499.6]
  assign _GEN_42 = _T_1068 ? _T_1069 : regs_42; // @[SRAM.scala 148:48:@42498.4]
  assign _T_1075 = io_waddr == 6'h2b; // @[SRAM.scala 148:37:@42506.4]
  assign _T_1076 = io_wen & _T_1075; // @[SRAM.scala 148:25:@42507.4]
  assign _T_1077 = io_banks_43_wdata_valid | _T_1076; // @[SRAM.scala 148:15:@42508.4]
  assign _T_1078 = io_banks_43_wdata_valid ? io_banks_43_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42510.6]
  assign _GEN_43 = _T_1077 ? _T_1078 : regs_43; // @[SRAM.scala 148:48:@42509.4]
  assign _T_1084 = io_waddr == 6'h2c; // @[SRAM.scala 148:37:@42517.4]
  assign _T_1085 = io_wen & _T_1084; // @[SRAM.scala 148:25:@42518.4]
  assign _T_1086 = io_banks_44_wdata_valid | _T_1085; // @[SRAM.scala 148:15:@42519.4]
  assign _T_1087 = io_banks_44_wdata_valid ? io_banks_44_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42521.6]
  assign _GEN_44 = _T_1086 ? _T_1087 : regs_44; // @[SRAM.scala 148:48:@42520.4]
  assign _T_1093 = io_waddr == 6'h2d; // @[SRAM.scala 148:37:@42528.4]
  assign _T_1094 = io_wen & _T_1093; // @[SRAM.scala 148:25:@42529.4]
  assign _T_1095 = io_banks_45_wdata_valid | _T_1094; // @[SRAM.scala 148:15:@42530.4]
  assign _T_1096 = io_banks_45_wdata_valid ? io_banks_45_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42532.6]
  assign _GEN_45 = _T_1095 ? _T_1096 : regs_45; // @[SRAM.scala 148:48:@42531.4]
  assign _T_1102 = io_waddr == 6'h2e; // @[SRAM.scala 148:37:@42539.4]
  assign _T_1103 = io_wen & _T_1102; // @[SRAM.scala 148:25:@42540.4]
  assign _T_1104 = io_banks_46_wdata_valid | _T_1103; // @[SRAM.scala 148:15:@42541.4]
  assign _T_1105 = io_banks_46_wdata_valid ? io_banks_46_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42543.6]
  assign _GEN_46 = _T_1104 ? _T_1105 : regs_46; // @[SRAM.scala 148:48:@42542.4]
  assign _T_1111 = io_waddr == 6'h2f; // @[SRAM.scala 148:37:@42550.4]
  assign _T_1112 = io_wen & _T_1111; // @[SRAM.scala 148:25:@42551.4]
  assign _T_1113 = io_banks_47_wdata_valid | _T_1112; // @[SRAM.scala 148:15:@42552.4]
  assign _T_1114 = io_banks_47_wdata_valid ? io_banks_47_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42554.6]
  assign _GEN_47 = _T_1113 ? _T_1114 : regs_47; // @[SRAM.scala 148:48:@42553.4]
  assign _T_1120 = io_waddr == 6'h30; // @[SRAM.scala 148:37:@42561.4]
  assign _T_1121 = io_wen & _T_1120; // @[SRAM.scala 148:25:@42562.4]
  assign _T_1122 = io_banks_48_wdata_valid | _T_1121; // @[SRAM.scala 148:15:@42563.4]
  assign _T_1123 = io_banks_48_wdata_valid ? io_banks_48_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42565.6]
  assign _GEN_48 = _T_1122 ? _T_1123 : regs_48; // @[SRAM.scala 148:48:@42564.4]
  assign _T_1129 = io_waddr == 6'h31; // @[SRAM.scala 148:37:@42572.4]
  assign _T_1130 = io_wen & _T_1129; // @[SRAM.scala 148:25:@42573.4]
  assign _T_1131 = io_banks_49_wdata_valid | _T_1130; // @[SRAM.scala 148:15:@42574.4]
  assign _T_1132 = io_banks_49_wdata_valid ? io_banks_49_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42576.6]
  assign _GEN_49 = _T_1131 ? _T_1132 : regs_49; // @[SRAM.scala 148:48:@42575.4]
  assign _T_1138 = io_waddr == 6'h32; // @[SRAM.scala 148:37:@42583.4]
  assign _T_1139 = io_wen & _T_1138; // @[SRAM.scala 148:25:@42584.4]
  assign _T_1140 = io_banks_50_wdata_valid | _T_1139; // @[SRAM.scala 148:15:@42585.4]
  assign _T_1141 = io_banks_50_wdata_valid ? io_banks_50_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42587.6]
  assign _GEN_50 = _T_1140 ? _T_1141 : regs_50; // @[SRAM.scala 148:48:@42586.4]
  assign _T_1147 = io_waddr == 6'h33; // @[SRAM.scala 148:37:@42594.4]
  assign _T_1148 = io_wen & _T_1147; // @[SRAM.scala 148:25:@42595.4]
  assign _T_1149 = io_banks_51_wdata_valid | _T_1148; // @[SRAM.scala 148:15:@42596.4]
  assign _T_1150 = io_banks_51_wdata_valid ? io_banks_51_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42598.6]
  assign _GEN_51 = _T_1149 ? _T_1150 : regs_51; // @[SRAM.scala 148:48:@42597.4]
  assign _T_1156 = io_waddr == 6'h34; // @[SRAM.scala 148:37:@42605.4]
  assign _T_1157 = io_wen & _T_1156; // @[SRAM.scala 148:25:@42606.4]
  assign _T_1158 = io_banks_52_wdata_valid | _T_1157; // @[SRAM.scala 148:15:@42607.4]
  assign _T_1159 = io_banks_52_wdata_valid ? io_banks_52_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42609.6]
  assign _GEN_52 = _T_1158 ? _T_1159 : regs_52; // @[SRAM.scala 148:48:@42608.4]
  assign _T_1165 = io_waddr == 6'h35; // @[SRAM.scala 148:37:@42616.4]
  assign _T_1166 = io_wen & _T_1165; // @[SRAM.scala 148:25:@42617.4]
  assign _T_1167 = io_banks_53_wdata_valid | _T_1166; // @[SRAM.scala 148:15:@42618.4]
  assign _T_1168 = io_banks_53_wdata_valid ? io_banks_53_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42620.6]
  assign _GEN_53 = _T_1167 ? _T_1168 : regs_53; // @[SRAM.scala 148:48:@42619.4]
  assign _T_1174 = io_waddr == 6'h36; // @[SRAM.scala 148:37:@42627.4]
  assign _T_1175 = io_wen & _T_1174; // @[SRAM.scala 148:25:@42628.4]
  assign _T_1176 = io_banks_54_wdata_valid | _T_1175; // @[SRAM.scala 148:15:@42629.4]
  assign _T_1177 = io_banks_54_wdata_valid ? io_banks_54_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42631.6]
  assign _GEN_54 = _T_1176 ? _T_1177 : regs_54; // @[SRAM.scala 148:48:@42630.4]
  assign _T_1183 = io_waddr == 6'h37; // @[SRAM.scala 148:37:@42638.4]
  assign _T_1184 = io_wen & _T_1183; // @[SRAM.scala 148:25:@42639.4]
  assign _T_1185 = io_banks_55_wdata_valid | _T_1184; // @[SRAM.scala 148:15:@42640.4]
  assign _T_1186 = io_banks_55_wdata_valid ? io_banks_55_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42642.6]
  assign _GEN_55 = _T_1185 ? _T_1186 : regs_55; // @[SRAM.scala 148:48:@42641.4]
  assign _T_1192 = io_waddr == 6'h38; // @[SRAM.scala 148:37:@42649.4]
  assign _T_1193 = io_wen & _T_1192; // @[SRAM.scala 148:25:@42650.4]
  assign _T_1194 = io_banks_56_wdata_valid | _T_1193; // @[SRAM.scala 148:15:@42651.4]
  assign _T_1195 = io_banks_56_wdata_valid ? io_banks_56_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42653.6]
  assign _GEN_56 = _T_1194 ? _T_1195 : regs_56; // @[SRAM.scala 148:48:@42652.4]
  assign _T_1201 = io_waddr == 6'h39; // @[SRAM.scala 148:37:@42660.4]
  assign _T_1202 = io_wen & _T_1201; // @[SRAM.scala 148:25:@42661.4]
  assign _T_1203 = io_banks_57_wdata_valid | _T_1202; // @[SRAM.scala 148:15:@42662.4]
  assign _T_1204 = io_banks_57_wdata_valid ? io_banks_57_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42664.6]
  assign _GEN_57 = _T_1203 ? _T_1204 : regs_57; // @[SRAM.scala 148:48:@42663.4]
  assign _T_1210 = io_waddr == 6'h3a; // @[SRAM.scala 148:37:@42671.4]
  assign _T_1211 = io_wen & _T_1210; // @[SRAM.scala 148:25:@42672.4]
  assign _T_1212 = io_banks_58_wdata_valid | _T_1211; // @[SRAM.scala 148:15:@42673.4]
  assign _T_1213 = io_banks_58_wdata_valid ? io_banks_58_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42675.6]
  assign _GEN_58 = _T_1212 ? _T_1213 : regs_58; // @[SRAM.scala 148:48:@42674.4]
  assign _T_1219 = io_waddr == 6'h3b; // @[SRAM.scala 148:37:@42682.4]
  assign _T_1220 = io_wen & _T_1219; // @[SRAM.scala 148:25:@42683.4]
  assign _T_1221 = io_banks_59_wdata_valid | _T_1220; // @[SRAM.scala 148:15:@42684.4]
  assign _T_1222 = io_banks_59_wdata_valid ? io_banks_59_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42686.6]
  assign _GEN_59 = _T_1221 ? _T_1222 : regs_59; // @[SRAM.scala 148:48:@42685.4]
  assign _T_1228 = io_waddr == 6'h3c; // @[SRAM.scala 148:37:@42693.4]
  assign _T_1229 = io_wen & _T_1228; // @[SRAM.scala 148:25:@42694.4]
  assign _T_1230 = io_banks_60_wdata_valid | _T_1229; // @[SRAM.scala 148:15:@42695.4]
  assign _T_1231 = io_banks_60_wdata_valid ? io_banks_60_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42697.6]
  assign _GEN_60 = _T_1230 ? _T_1231 : regs_60; // @[SRAM.scala 148:48:@42696.4]
  assign _T_1237 = io_waddr == 6'h3d; // @[SRAM.scala 148:37:@42704.4]
  assign _T_1238 = io_wen & _T_1237; // @[SRAM.scala 148:25:@42705.4]
  assign _T_1239 = io_banks_61_wdata_valid | _T_1238; // @[SRAM.scala 148:15:@42706.4]
  assign _T_1240 = io_banks_61_wdata_valid ? io_banks_61_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42708.6]
  assign _GEN_61 = _T_1239 ? _T_1240 : regs_61; // @[SRAM.scala 148:48:@42707.4]
  assign _T_1246 = io_waddr == 6'h3e; // @[SRAM.scala 148:37:@42715.4]
  assign _T_1247 = io_wen & _T_1246; // @[SRAM.scala 148:25:@42716.4]
  assign _T_1248 = io_banks_62_wdata_valid | _T_1247; // @[SRAM.scala 148:15:@42717.4]
  assign _T_1249 = io_banks_62_wdata_valid ? io_banks_62_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42719.6]
  assign _GEN_62 = _T_1248 ? _T_1249 : regs_62; // @[SRAM.scala 148:48:@42718.4]
  assign _T_1255 = io_waddr == 6'h3f; // @[SRAM.scala 148:37:@42726.4]
  assign _T_1256 = io_wen & _T_1255; // @[SRAM.scala 148:25:@42727.4]
  assign _T_1257 = io_banks_63_wdata_valid | _T_1256; // @[SRAM.scala 148:15:@42728.4]
  assign _T_1258 = io_banks_63_wdata_valid ? io_banks_63_wdata_bits : io_wdata; // @[SRAM.scala 149:15:@42730.6]
  assign _GEN_63 = _T_1257 ? _T_1258 : regs_63; // @[SRAM.scala 148:48:@42729.4]
  assign _GEN_65 = 6'h1 == io_raddr ? regs_1 : regs_0; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_66 = 6'h2 == io_raddr ? regs_2 : _GEN_65; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_67 = 6'h3 == io_raddr ? regs_3 : _GEN_66; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_68 = 6'h4 == io_raddr ? regs_4 : _GEN_67; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_69 = 6'h5 == io_raddr ? regs_5 : _GEN_68; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_70 = 6'h6 == io_raddr ? regs_6 : _GEN_69; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_71 = 6'h7 == io_raddr ? regs_7 : _GEN_70; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_72 = 6'h8 == io_raddr ? regs_8 : _GEN_71; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_73 = 6'h9 == io_raddr ? regs_9 : _GEN_72; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_74 = 6'ha == io_raddr ? regs_10 : _GEN_73; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_75 = 6'hb == io_raddr ? regs_11 : _GEN_74; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_76 = 6'hc == io_raddr ? regs_12 : _GEN_75; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_77 = 6'hd == io_raddr ? regs_13 : _GEN_76; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_78 = 6'he == io_raddr ? regs_14 : _GEN_77; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_79 = 6'hf == io_raddr ? regs_15 : _GEN_78; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_80 = 6'h10 == io_raddr ? regs_16 : _GEN_79; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_81 = 6'h11 == io_raddr ? regs_17 : _GEN_80; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_82 = 6'h12 == io_raddr ? regs_18 : _GEN_81; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_83 = 6'h13 == io_raddr ? regs_19 : _GEN_82; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_84 = 6'h14 == io_raddr ? regs_20 : _GEN_83; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_85 = 6'h15 == io_raddr ? regs_21 : _GEN_84; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_86 = 6'h16 == io_raddr ? regs_22 : _GEN_85; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_87 = 6'h17 == io_raddr ? regs_23 : _GEN_86; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_88 = 6'h18 == io_raddr ? regs_24 : _GEN_87; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_89 = 6'h19 == io_raddr ? regs_25 : _GEN_88; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_90 = 6'h1a == io_raddr ? regs_26 : _GEN_89; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_91 = 6'h1b == io_raddr ? regs_27 : _GEN_90; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_92 = 6'h1c == io_raddr ? regs_28 : _GEN_91; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_93 = 6'h1d == io_raddr ? regs_29 : _GEN_92; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_94 = 6'h1e == io_raddr ? regs_30 : _GEN_93; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_95 = 6'h1f == io_raddr ? regs_31 : _GEN_94; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_96 = 6'h20 == io_raddr ? regs_32 : _GEN_95; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_97 = 6'h21 == io_raddr ? regs_33 : _GEN_96; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_98 = 6'h22 == io_raddr ? regs_34 : _GEN_97; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_99 = 6'h23 == io_raddr ? regs_35 : _GEN_98; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_100 = 6'h24 == io_raddr ? regs_36 : _GEN_99; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_101 = 6'h25 == io_raddr ? regs_37 : _GEN_100; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_102 = 6'h26 == io_raddr ? regs_38 : _GEN_101; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_103 = 6'h27 == io_raddr ? regs_39 : _GEN_102; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_104 = 6'h28 == io_raddr ? regs_40 : _GEN_103; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_105 = 6'h29 == io_raddr ? regs_41 : _GEN_104; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_106 = 6'h2a == io_raddr ? regs_42 : _GEN_105; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_107 = 6'h2b == io_raddr ? regs_43 : _GEN_106; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_108 = 6'h2c == io_raddr ? regs_44 : _GEN_107; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_109 = 6'h2d == io_raddr ? regs_45 : _GEN_108; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_110 = 6'h2e == io_raddr ? regs_46 : _GEN_109; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_111 = 6'h2f == io_raddr ? regs_47 : _GEN_110; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_112 = 6'h30 == io_raddr ? regs_48 : _GEN_111; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_113 = 6'h31 == io_raddr ? regs_49 : _GEN_112; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_114 = 6'h32 == io_raddr ? regs_50 : _GEN_113; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_115 = 6'h33 == io_raddr ? regs_51 : _GEN_114; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_116 = 6'h34 == io_raddr ? regs_52 : _GEN_115; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_117 = 6'h35 == io_raddr ? regs_53 : _GEN_116; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_118 = 6'h36 == io_raddr ? regs_54 : _GEN_117; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_119 = 6'h37 == io_raddr ? regs_55 : _GEN_118; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_120 = 6'h38 == io_raddr ? regs_56 : _GEN_119; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_121 = 6'h39 == io_raddr ? regs_57 : _GEN_120; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_122 = 6'h3a == io_raddr ? regs_58 : _GEN_121; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_123 = 6'h3b == io_raddr ? regs_59 : _GEN_122; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_124 = 6'h3c == io_raddr ? regs_60 : _GEN_123; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_125 = 6'h3d == io_raddr ? regs_61 : _GEN_124; // @[SRAM.scala 155:12:@42799.4]
  assign _GEN_126 = 6'h3e == io_raddr ? regs_62 : _GEN_125; // @[SRAM.scala 155:12:@42799.4]
  assign io_rdata = 6'h3f == io_raddr ? regs_63 : _GEN_126; // @[SRAM.scala 155:12:@42799.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regs_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regs_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regs_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regs_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regs_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regs_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regs_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regs_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regs_8 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regs_9 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regs_10 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regs_11 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regs_12 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regs_13 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regs_14 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regs_15 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regs_16 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regs_17 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regs_18 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regs_19 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regs_20 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regs_21 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regs_22 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regs_23 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regs_24 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regs_25 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regs_26 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regs_27 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regs_28 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regs_29 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regs_30 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regs_31 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  regs_32 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  regs_33 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  regs_34 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  regs_35 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  regs_36 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  regs_37 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  regs_38 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  regs_39 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  regs_40 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  regs_41 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  regs_42 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  regs_43 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  regs_44 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  regs_45 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  regs_46 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  regs_47 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  regs_48 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  regs_49 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  regs_50 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  regs_51 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  regs_52 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  regs_53 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  regs_54 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  regs_55 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  regs_56 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  regs_57 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  regs_58 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  regs_59 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  regs_60 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  regs_61 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  regs_62 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  regs_63 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      regs_0 <= 1'h0;
    end else begin
      if (_T_690) begin
        if (io_banks_0_wdata_valid) begin
          regs_0 <= io_banks_0_wdata_bits;
        end else begin
          regs_0 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_1 <= 1'h0;
    end else begin
      if (_T_699) begin
        if (io_banks_1_wdata_valid) begin
          regs_1 <= io_banks_1_wdata_bits;
        end else begin
          regs_1 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_2 <= 1'h0;
    end else begin
      if (_T_708) begin
        if (io_banks_2_wdata_valid) begin
          regs_2 <= io_banks_2_wdata_bits;
        end else begin
          regs_2 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_3 <= 1'h0;
    end else begin
      if (_T_717) begin
        if (io_banks_3_wdata_valid) begin
          regs_3 <= io_banks_3_wdata_bits;
        end else begin
          regs_3 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_4 <= 1'h0;
    end else begin
      if (_T_726) begin
        if (io_banks_4_wdata_valid) begin
          regs_4 <= io_banks_4_wdata_bits;
        end else begin
          regs_4 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_5 <= 1'h0;
    end else begin
      if (_T_735) begin
        if (io_banks_5_wdata_valid) begin
          regs_5 <= io_banks_5_wdata_bits;
        end else begin
          regs_5 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_6 <= 1'h0;
    end else begin
      if (_T_744) begin
        if (io_banks_6_wdata_valid) begin
          regs_6 <= io_banks_6_wdata_bits;
        end else begin
          regs_6 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_7 <= 1'h0;
    end else begin
      if (_T_753) begin
        if (io_banks_7_wdata_valid) begin
          regs_7 <= io_banks_7_wdata_bits;
        end else begin
          regs_7 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_8 <= 1'h0;
    end else begin
      if (_T_762) begin
        if (io_banks_8_wdata_valid) begin
          regs_8 <= io_banks_8_wdata_bits;
        end else begin
          regs_8 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_9 <= 1'h0;
    end else begin
      if (_T_771) begin
        if (io_banks_9_wdata_valid) begin
          regs_9 <= io_banks_9_wdata_bits;
        end else begin
          regs_9 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_10 <= 1'h0;
    end else begin
      if (_T_780) begin
        if (io_banks_10_wdata_valid) begin
          regs_10 <= io_banks_10_wdata_bits;
        end else begin
          regs_10 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_11 <= 1'h0;
    end else begin
      if (_T_789) begin
        if (io_banks_11_wdata_valid) begin
          regs_11 <= io_banks_11_wdata_bits;
        end else begin
          regs_11 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_12 <= 1'h0;
    end else begin
      if (_T_798) begin
        if (io_banks_12_wdata_valid) begin
          regs_12 <= io_banks_12_wdata_bits;
        end else begin
          regs_12 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_13 <= 1'h0;
    end else begin
      if (_T_807) begin
        if (io_banks_13_wdata_valid) begin
          regs_13 <= io_banks_13_wdata_bits;
        end else begin
          regs_13 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_14 <= 1'h0;
    end else begin
      if (_T_816) begin
        if (io_banks_14_wdata_valid) begin
          regs_14 <= io_banks_14_wdata_bits;
        end else begin
          regs_14 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_15 <= 1'h0;
    end else begin
      if (_T_825) begin
        if (io_banks_15_wdata_valid) begin
          regs_15 <= io_banks_15_wdata_bits;
        end else begin
          regs_15 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_16 <= 1'h0;
    end else begin
      if (_T_834) begin
        if (io_banks_16_wdata_valid) begin
          regs_16 <= io_banks_16_wdata_bits;
        end else begin
          regs_16 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_17 <= 1'h0;
    end else begin
      if (_T_843) begin
        if (io_banks_17_wdata_valid) begin
          regs_17 <= io_banks_17_wdata_bits;
        end else begin
          regs_17 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_18 <= 1'h0;
    end else begin
      if (_T_852) begin
        if (io_banks_18_wdata_valid) begin
          regs_18 <= io_banks_18_wdata_bits;
        end else begin
          regs_18 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_19 <= 1'h0;
    end else begin
      if (_T_861) begin
        if (io_banks_19_wdata_valid) begin
          regs_19 <= io_banks_19_wdata_bits;
        end else begin
          regs_19 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_20 <= 1'h0;
    end else begin
      if (_T_870) begin
        if (io_banks_20_wdata_valid) begin
          regs_20 <= io_banks_20_wdata_bits;
        end else begin
          regs_20 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_21 <= 1'h0;
    end else begin
      if (_T_879) begin
        if (io_banks_21_wdata_valid) begin
          regs_21 <= io_banks_21_wdata_bits;
        end else begin
          regs_21 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_22 <= 1'h0;
    end else begin
      if (_T_888) begin
        if (io_banks_22_wdata_valid) begin
          regs_22 <= io_banks_22_wdata_bits;
        end else begin
          regs_22 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_23 <= 1'h0;
    end else begin
      if (_T_897) begin
        if (io_banks_23_wdata_valid) begin
          regs_23 <= io_banks_23_wdata_bits;
        end else begin
          regs_23 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_24 <= 1'h0;
    end else begin
      if (_T_906) begin
        if (io_banks_24_wdata_valid) begin
          regs_24 <= io_banks_24_wdata_bits;
        end else begin
          regs_24 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_25 <= 1'h0;
    end else begin
      if (_T_915) begin
        if (io_banks_25_wdata_valid) begin
          regs_25 <= io_banks_25_wdata_bits;
        end else begin
          regs_25 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_26 <= 1'h0;
    end else begin
      if (_T_924) begin
        if (io_banks_26_wdata_valid) begin
          regs_26 <= io_banks_26_wdata_bits;
        end else begin
          regs_26 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_27 <= 1'h0;
    end else begin
      if (_T_933) begin
        if (io_banks_27_wdata_valid) begin
          regs_27 <= io_banks_27_wdata_bits;
        end else begin
          regs_27 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_28 <= 1'h0;
    end else begin
      if (_T_942) begin
        if (io_banks_28_wdata_valid) begin
          regs_28 <= io_banks_28_wdata_bits;
        end else begin
          regs_28 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_29 <= 1'h0;
    end else begin
      if (_T_951) begin
        if (io_banks_29_wdata_valid) begin
          regs_29 <= io_banks_29_wdata_bits;
        end else begin
          regs_29 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_30 <= 1'h0;
    end else begin
      if (_T_960) begin
        if (io_banks_30_wdata_valid) begin
          regs_30 <= io_banks_30_wdata_bits;
        end else begin
          regs_30 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_31 <= 1'h0;
    end else begin
      if (_T_969) begin
        if (io_banks_31_wdata_valid) begin
          regs_31 <= io_banks_31_wdata_bits;
        end else begin
          regs_31 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_32 <= 1'h0;
    end else begin
      if (_T_978) begin
        if (io_banks_32_wdata_valid) begin
          regs_32 <= io_banks_32_wdata_bits;
        end else begin
          regs_32 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_33 <= 1'h0;
    end else begin
      if (_T_987) begin
        if (io_banks_33_wdata_valid) begin
          regs_33 <= io_banks_33_wdata_bits;
        end else begin
          regs_33 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_34 <= 1'h0;
    end else begin
      if (_T_996) begin
        if (io_banks_34_wdata_valid) begin
          regs_34 <= io_banks_34_wdata_bits;
        end else begin
          regs_34 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_35 <= 1'h0;
    end else begin
      if (_T_1005) begin
        if (io_banks_35_wdata_valid) begin
          regs_35 <= io_banks_35_wdata_bits;
        end else begin
          regs_35 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_36 <= 1'h0;
    end else begin
      if (_T_1014) begin
        if (io_banks_36_wdata_valid) begin
          regs_36 <= io_banks_36_wdata_bits;
        end else begin
          regs_36 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_37 <= 1'h0;
    end else begin
      if (_T_1023) begin
        if (io_banks_37_wdata_valid) begin
          regs_37 <= io_banks_37_wdata_bits;
        end else begin
          regs_37 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_38 <= 1'h0;
    end else begin
      if (_T_1032) begin
        if (io_banks_38_wdata_valid) begin
          regs_38 <= io_banks_38_wdata_bits;
        end else begin
          regs_38 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_39 <= 1'h0;
    end else begin
      if (_T_1041) begin
        if (io_banks_39_wdata_valid) begin
          regs_39 <= io_banks_39_wdata_bits;
        end else begin
          regs_39 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_40 <= 1'h0;
    end else begin
      if (_T_1050) begin
        if (io_banks_40_wdata_valid) begin
          regs_40 <= io_banks_40_wdata_bits;
        end else begin
          regs_40 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_41 <= 1'h0;
    end else begin
      if (_T_1059) begin
        if (io_banks_41_wdata_valid) begin
          regs_41 <= io_banks_41_wdata_bits;
        end else begin
          regs_41 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_42 <= 1'h0;
    end else begin
      if (_T_1068) begin
        if (io_banks_42_wdata_valid) begin
          regs_42 <= io_banks_42_wdata_bits;
        end else begin
          regs_42 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_43 <= 1'h0;
    end else begin
      if (_T_1077) begin
        if (io_banks_43_wdata_valid) begin
          regs_43 <= io_banks_43_wdata_bits;
        end else begin
          regs_43 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_44 <= 1'h0;
    end else begin
      if (_T_1086) begin
        if (io_banks_44_wdata_valid) begin
          regs_44 <= io_banks_44_wdata_bits;
        end else begin
          regs_44 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_45 <= 1'h0;
    end else begin
      if (_T_1095) begin
        if (io_banks_45_wdata_valid) begin
          regs_45 <= io_banks_45_wdata_bits;
        end else begin
          regs_45 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_46 <= 1'h0;
    end else begin
      if (_T_1104) begin
        if (io_banks_46_wdata_valid) begin
          regs_46 <= io_banks_46_wdata_bits;
        end else begin
          regs_46 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_47 <= 1'h0;
    end else begin
      if (_T_1113) begin
        if (io_banks_47_wdata_valid) begin
          regs_47 <= io_banks_47_wdata_bits;
        end else begin
          regs_47 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_48 <= 1'h0;
    end else begin
      if (_T_1122) begin
        if (io_banks_48_wdata_valid) begin
          regs_48 <= io_banks_48_wdata_bits;
        end else begin
          regs_48 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_49 <= 1'h0;
    end else begin
      if (_T_1131) begin
        if (io_banks_49_wdata_valid) begin
          regs_49 <= io_banks_49_wdata_bits;
        end else begin
          regs_49 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_50 <= 1'h0;
    end else begin
      if (_T_1140) begin
        if (io_banks_50_wdata_valid) begin
          regs_50 <= io_banks_50_wdata_bits;
        end else begin
          regs_50 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_51 <= 1'h0;
    end else begin
      if (_T_1149) begin
        if (io_banks_51_wdata_valid) begin
          regs_51 <= io_banks_51_wdata_bits;
        end else begin
          regs_51 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_52 <= 1'h0;
    end else begin
      if (_T_1158) begin
        if (io_banks_52_wdata_valid) begin
          regs_52 <= io_banks_52_wdata_bits;
        end else begin
          regs_52 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_53 <= 1'h0;
    end else begin
      if (_T_1167) begin
        if (io_banks_53_wdata_valid) begin
          regs_53 <= io_banks_53_wdata_bits;
        end else begin
          regs_53 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_54 <= 1'h0;
    end else begin
      if (_T_1176) begin
        if (io_banks_54_wdata_valid) begin
          regs_54 <= io_banks_54_wdata_bits;
        end else begin
          regs_54 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_55 <= 1'h0;
    end else begin
      if (_T_1185) begin
        if (io_banks_55_wdata_valid) begin
          regs_55 <= io_banks_55_wdata_bits;
        end else begin
          regs_55 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_56 <= 1'h0;
    end else begin
      if (_T_1194) begin
        if (io_banks_56_wdata_valid) begin
          regs_56 <= io_banks_56_wdata_bits;
        end else begin
          regs_56 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_57 <= 1'h0;
    end else begin
      if (_T_1203) begin
        if (io_banks_57_wdata_valid) begin
          regs_57 <= io_banks_57_wdata_bits;
        end else begin
          regs_57 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_58 <= 1'h0;
    end else begin
      if (_T_1212) begin
        if (io_banks_58_wdata_valid) begin
          regs_58 <= io_banks_58_wdata_bits;
        end else begin
          regs_58 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_59 <= 1'h0;
    end else begin
      if (_T_1221) begin
        if (io_banks_59_wdata_valid) begin
          regs_59 <= io_banks_59_wdata_bits;
        end else begin
          regs_59 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_60 <= 1'h0;
    end else begin
      if (_T_1230) begin
        if (io_banks_60_wdata_valid) begin
          regs_60 <= io_banks_60_wdata_bits;
        end else begin
          regs_60 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_61 <= 1'h0;
    end else begin
      if (_T_1239) begin
        if (io_banks_61_wdata_valid) begin
          regs_61 <= io_banks_61_wdata_bits;
        end else begin
          regs_61 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_62 <= 1'h0;
    end else begin
      if (_T_1248) begin
        if (io_banks_62_wdata_valid) begin
          regs_62 <= io_banks_62_wdata_bits;
        end else begin
          regs_62 <= io_wdata;
        end
      end
    end
    if (reset) begin
      regs_63 <= 1'h0;
    end else begin
      if (_T_1257) begin
        if (io_banks_63_wdata_valid) begin
          regs_63 <= io_banks_63_wdata_bits;
        end else begin
          regs_63 <= io_wdata;
        end
      end
    end
  end
endmodule
module FIFO_33( // @[:@42801.2]
  input   clock, // @[:@42802.4]
  input   reset, // @[:@42803.4]
  output  io_in_ready, // @[:@42804.4]
  input   io_in_valid, // @[:@42804.4]
  input   io_in_bits, // @[:@42804.4]
  input   io_out_ready, // @[:@42804.4]
  output  io_out_valid, // @[:@42804.4]
  output  io_out_bits, // @[:@42804.4]
  input   io_banks_0_wdata_valid, // @[:@42804.4]
  input   io_banks_0_wdata_bits, // @[:@42804.4]
  input   io_banks_1_wdata_valid, // @[:@42804.4]
  input   io_banks_1_wdata_bits, // @[:@42804.4]
  input   io_banks_2_wdata_valid, // @[:@42804.4]
  input   io_banks_2_wdata_bits, // @[:@42804.4]
  input   io_banks_3_wdata_valid, // @[:@42804.4]
  input   io_banks_3_wdata_bits, // @[:@42804.4]
  input   io_banks_4_wdata_valid, // @[:@42804.4]
  input   io_banks_4_wdata_bits, // @[:@42804.4]
  input   io_banks_5_wdata_valid, // @[:@42804.4]
  input   io_banks_5_wdata_bits, // @[:@42804.4]
  input   io_banks_6_wdata_valid, // @[:@42804.4]
  input   io_banks_6_wdata_bits, // @[:@42804.4]
  input   io_banks_7_wdata_valid, // @[:@42804.4]
  input   io_banks_7_wdata_bits, // @[:@42804.4]
  input   io_banks_8_wdata_valid, // @[:@42804.4]
  input   io_banks_8_wdata_bits, // @[:@42804.4]
  input   io_banks_9_wdata_valid, // @[:@42804.4]
  input   io_banks_9_wdata_bits, // @[:@42804.4]
  input   io_banks_10_wdata_valid, // @[:@42804.4]
  input   io_banks_10_wdata_bits, // @[:@42804.4]
  input   io_banks_11_wdata_valid, // @[:@42804.4]
  input   io_banks_11_wdata_bits, // @[:@42804.4]
  input   io_banks_12_wdata_valid, // @[:@42804.4]
  input   io_banks_12_wdata_bits, // @[:@42804.4]
  input   io_banks_13_wdata_valid, // @[:@42804.4]
  input   io_banks_13_wdata_bits, // @[:@42804.4]
  input   io_banks_14_wdata_valid, // @[:@42804.4]
  input   io_banks_14_wdata_bits, // @[:@42804.4]
  input   io_banks_15_wdata_valid, // @[:@42804.4]
  input   io_banks_15_wdata_bits, // @[:@42804.4]
  input   io_banks_16_wdata_valid, // @[:@42804.4]
  input   io_banks_16_wdata_bits, // @[:@42804.4]
  input   io_banks_17_wdata_valid, // @[:@42804.4]
  input   io_banks_17_wdata_bits, // @[:@42804.4]
  input   io_banks_18_wdata_valid, // @[:@42804.4]
  input   io_banks_18_wdata_bits, // @[:@42804.4]
  input   io_banks_19_wdata_valid, // @[:@42804.4]
  input   io_banks_19_wdata_bits, // @[:@42804.4]
  input   io_banks_20_wdata_valid, // @[:@42804.4]
  input   io_banks_20_wdata_bits, // @[:@42804.4]
  input   io_banks_21_wdata_valid, // @[:@42804.4]
  input   io_banks_21_wdata_bits, // @[:@42804.4]
  input   io_banks_22_wdata_valid, // @[:@42804.4]
  input   io_banks_22_wdata_bits, // @[:@42804.4]
  input   io_banks_23_wdata_valid, // @[:@42804.4]
  input   io_banks_23_wdata_bits, // @[:@42804.4]
  input   io_banks_24_wdata_valid, // @[:@42804.4]
  input   io_banks_24_wdata_bits, // @[:@42804.4]
  input   io_banks_25_wdata_valid, // @[:@42804.4]
  input   io_banks_25_wdata_bits, // @[:@42804.4]
  input   io_banks_26_wdata_valid, // @[:@42804.4]
  input   io_banks_26_wdata_bits, // @[:@42804.4]
  input   io_banks_27_wdata_valid, // @[:@42804.4]
  input   io_banks_27_wdata_bits, // @[:@42804.4]
  input   io_banks_28_wdata_valid, // @[:@42804.4]
  input   io_banks_28_wdata_bits, // @[:@42804.4]
  input   io_banks_29_wdata_valid, // @[:@42804.4]
  input   io_banks_29_wdata_bits, // @[:@42804.4]
  input   io_banks_30_wdata_valid, // @[:@42804.4]
  input   io_banks_30_wdata_bits, // @[:@42804.4]
  input   io_banks_31_wdata_valid, // @[:@42804.4]
  input   io_banks_31_wdata_bits, // @[:@42804.4]
  input   io_banks_32_wdata_valid, // @[:@42804.4]
  input   io_banks_32_wdata_bits, // @[:@42804.4]
  input   io_banks_33_wdata_valid, // @[:@42804.4]
  input   io_banks_33_wdata_bits, // @[:@42804.4]
  input   io_banks_34_wdata_valid, // @[:@42804.4]
  input   io_banks_34_wdata_bits, // @[:@42804.4]
  input   io_banks_35_wdata_valid, // @[:@42804.4]
  input   io_banks_35_wdata_bits, // @[:@42804.4]
  input   io_banks_36_wdata_valid, // @[:@42804.4]
  input   io_banks_36_wdata_bits, // @[:@42804.4]
  input   io_banks_37_wdata_valid, // @[:@42804.4]
  input   io_banks_37_wdata_bits, // @[:@42804.4]
  input   io_banks_38_wdata_valid, // @[:@42804.4]
  input   io_banks_38_wdata_bits, // @[:@42804.4]
  input   io_banks_39_wdata_valid, // @[:@42804.4]
  input   io_banks_39_wdata_bits, // @[:@42804.4]
  input   io_banks_40_wdata_valid, // @[:@42804.4]
  input   io_banks_40_wdata_bits, // @[:@42804.4]
  input   io_banks_41_wdata_valid, // @[:@42804.4]
  input   io_banks_41_wdata_bits, // @[:@42804.4]
  input   io_banks_42_wdata_valid, // @[:@42804.4]
  input   io_banks_42_wdata_bits, // @[:@42804.4]
  input   io_banks_43_wdata_valid, // @[:@42804.4]
  input   io_banks_43_wdata_bits, // @[:@42804.4]
  input   io_banks_44_wdata_valid, // @[:@42804.4]
  input   io_banks_44_wdata_bits, // @[:@42804.4]
  input   io_banks_45_wdata_valid, // @[:@42804.4]
  input   io_banks_45_wdata_bits, // @[:@42804.4]
  input   io_banks_46_wdata_valid, // @[:@42804.4]
  input   io_banks_46_wdata_bits, // @[:@42804.4]
  input   io_banks_47_wdata_valid, // @[:@42804.4]
  input   io_banks_47_wdata_bits, // @[:@42804.4]
  input   io_banks_48_wdata_valid, // @[:@42804.4]
  input   io_banks_48_wdata_bits, // @[:@42804.4]
  input   io_banks_49_wdata_valid, // @[:@42804.4]
  input   io_banks_49_wdata_bits, // @[:@42804.4]
  input   io_banks_50_wdata_valid, // @[:@42804.4]
  input   io_banks_50_wdata_bits, // @[:@42804.4]
  input   io_banks_51_wdata_valid, // @[:@42804.4]
  input   io_banks_51_wdata_bits, // @[:@42804.4]
  input   io_banks_52_wdata_valid, // @[:@42804.4]
  input   io_banks_52_wdata_bits, // @[:@42804.4]
  input   io_banks_53_wdata_valid, // @[:@42804.4]
  input   io_banks_53_wdata_bits, // @[:@42804.4]
  input   io_banks_54_wdata_valid, // @[:@42804.4]
  input   io_banks_54_wdata_bits, // @[:@42804.4]
  input   io_banks_55_wdata_valid, // @[:@42804.4]
  input   io_banks_55_wdata_bits, // @[:@42804.4]
  input   io_banks_56_wdata_valid, // @[:@42804.4]
  input   io_banks_56_wdata_bits, // @[:@42804.4]
  input   io_banks_57_wdata_valid, // @[:@42804.4]
  input   io_banks_57_wdata_bits, // @[:@42804.4]
  input   io_banks_58_wdata_valid, // @[:@42804.4]
  input   io_banks_58_wdata_bits, // @[:@42804.4]
  input   io_banks_59_wdata_valid, // @[:@42804.4]
  input   io_banks_59_wdata_bits, // @[:@42804.4]
  input   io_banks_60_wdata_valid, // @[:@42804.4]
  input   io_banks_60_wdata_bits, // @[:@42804.4]
  input   io_banks_61_wdata_valid, // @[:@42804.4]
  input   io_banks_61_wdata_bits, // @[:@42804.4]
  input   io_banks_62_wdata_valid, // @[:@42804.4]
  input   io_banks_62_wdata_bits, // @[:@42804.4]
  input   io_banks_63_wdata_valid, // @[:@42804.4]
  input   io_banks_63_wdata_bits // @[:@42804.4]
);
  wire  enqCounter_clock; // @[FIFO.scala 34:26:@43070.4]
  wire  enqCounter_reset; // @[FIFO.scala 34:26:@43070.4]
  wire  enqCounter_io_enable; // @[FIFO.scala 34:26:@43070.4]
  wire [5:0] enqCounter_io_out; // @[FIFO.scala 34:26:@43070.4]
  wire [5:0] enqCounter_io_next; // @[FIFO.scala 34:26:@43070.4]
  wire  deqCounter_clock; // @[FIFO.scala 38:26:@43080.4]
  wire  deqCounter_reset; // @[FIFO.scala 38:26:@43080.4]
  wire  deqCounter_io_enable; // @[FIFO.scala 38:26:@43080.4]
  wire [5:0] deqCounter_io_out; // @[FIFO.scala 38:26:@43080.4]
  wire [5:0] deqCounter_io_next; // @[FIFO.scala 38:26:@43080.4]
  wire  FFRAM_clock; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_reset; // @[FIFO.scala 49:19:@43095.4]
  wire [5:0] FFRAM_io_raddr; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_wen; // @[FIFO.scala 49:19:@43095.4]
  wire [5:0] FFRAM_io_waddr; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_wdata; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_rdata; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_0_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_0_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_1_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_1_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_2_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_2_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_3_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_3_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_4_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_4_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_5_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_5_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_6_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_6_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_7_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_7_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_8_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_8_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_9_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_9_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_10_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_10_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_11_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_11_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_12_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_12_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_13_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_13_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_14_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_14_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_15_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_15_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_16_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_16_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_17_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_17_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_18_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_18_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_19_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_19_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_20_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_20_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_21_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_21_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_22_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_22_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_23_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_23_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_24_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_24_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_25_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_25_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_26_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_26_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_27_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_27_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_28_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_28_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_29_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_29_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_30_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_30_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_31_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_31_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_32_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_32_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_33_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_33_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_34_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_34_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_35_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_35_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_36_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_36_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_37_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_37_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_38_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_38_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_39_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_39_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_40_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_40_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_41_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_41_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_42_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_42_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_43_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_43_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_44_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_44_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_45_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_45_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_46_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_46_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_47_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_47_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_48_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_48_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_49_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_49_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_50_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_50_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_51_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_51_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_52_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_52_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_53_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_53_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_54_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_54_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_55_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_55_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_56_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_56_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_57_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_57_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_58_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_58_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_59_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_59_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_60_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_60_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_61_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_61_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_62_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_62_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_63_wdata_valid; // @[FIFO.scala 49:19:@43095.4]
  wire  FFRAM_io_banks_63_wdata_bits; // @[FIFO.scala 49:19:@43095.4]
  wire  writeEn; // @[FIFO.scala 30:29:@43068.4]
  wire  readEn; // @[FIFO.scala 31:29:@43069.4]
  reg  maybeFull; // @[FIFO.scala 42:26:@43090.4]
  reg [31:0] _RAND_0;
  wire  ptrMatch; // @[FIFO.scala 44:36:@43091.4]
  wire  _T_824; // @[FIFO.scala 45:27:@43092.4]
  wire  empty; // @[FIFO.scala 45:24:@43093.4]
  wire  full; // @[FIFO.scala 46:23:@43094.4]
  wire  _T_1657; // @[FIFO.scala 83:17:@44261.4]
  wire  _GEN_64; // @[FIFO.scala 83:29:@44262.4]
  Counter enqCounter ( // @[FIFO.scala 34:26:@43070.4]
    .clock(enqCounter_clock),
    .reset(enqCounter_reset),
    .io_enable(enqCounter_io_enable),
    .io_out(enqCounter_io_out),
    .io_next(enqCounter_io_next)
  );
  Counter deqCounter ( // @[FIFO.scala 38:26:@43080.4]
    .clock(deqCounter_clock),
    .reset(deqCounter_reset),
    .io_enable(deqCounter_io_enable),
    .io_out(deqCounter_io_out),
    .io_next(deqCounter_io_next)
  );
  FFRAM_16 FFRAM ( // @[FIFO.scala 49:19:@43095.4]
    .clock(FFRAM_clock),
    .reset(FFRAM_reset),
    .io_raddr(FFRAM_io_raddr),
    .io_wen(FFRAM_io_wen),
    .io_waddr(FFRAM_io_waddr),
    .io_wdata(FFRAM_io_wdata),
    .io_rdata(FFRAM_io_rdata),
    .io_banks_0_wdata_valid(FFRAM_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(FFRAM_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(FFRAM_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(FFRAM_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(FFRAM_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(FFRAM_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(FFRAM_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(FFRAM_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(FFRAM_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(FFRAM_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(FFRAM_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(FFRAM_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(FFRAM_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(FFRAM_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(FFRAM_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(FFRAM_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(FFRAM_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(FFRAM_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(FFRAM_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(FFRAM_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(FFRAM_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(FFRAM_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(FFRAM_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(FFRAM_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(FFRAM_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(FFRAM_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(FFRAM_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(FFRAM_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(FFRAM_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(FFRAM_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(FFRAM_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(FFRAM_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(FFRAM_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(FFRAM_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(FFRAM_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(FFRAM_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(FFRAM_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(FFRAM_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(FFRAM_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(FFRAM_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(FFRAM_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(FFRAM_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(FFRAM_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(FFRAM_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(FFRAM_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(FFRAM_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(FFRAM_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(FFRAM_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(FFRAM_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(FFRAM_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(FFRAM_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(FFRAM_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(FFRAM_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(FFRAM_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(FFRAM_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(FFRAM_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(FFRAM_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(FFRAM_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(FFRAM_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(FFRAM_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(FFRAM_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(FFRAM_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(FFRAM_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(FFRAM_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(FFRAM_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(FFRAM_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(FFRAM_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(FFRAM_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(FFRAM_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(FFRAM_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(FFRAM_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(FFRAM_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(FFRAM_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(FFRAM_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(FFRAM_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(FFRAM_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(FFRAM_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(FFRAM_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(FFRAM_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(FFRAM_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(FFRAM_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(FFRAM_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(FFRAM_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(FFRAM_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(FFRAM_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(FFRAM_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(FFRAM_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(FFRAM_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(FFRAM_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(FFRAM_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(FFRAM_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(FFRAM_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(FFRAM_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(FFRAM_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(FFRAM_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(FFRAM_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(FFRAM_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(FFRAM_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(FFRAM_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(FFRAM_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(FFRAM_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(FFRAM_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(FFRAM_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(FFRAM_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(FFRAM_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(FFRAM_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(FFRAM_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(FFRAM_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(FFRAM_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(FFRAM_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(FFRAM_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(FFRAM_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(FFRAM_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(FFRAM_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(FFRAM_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(FFRAM_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(FFRAM_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(FFRAM_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(FFRAM_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(FFRAM_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(FFRAM_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(FFRAM_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(FFRAM_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(FFRAM_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(FFRAM_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(FFRAM_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(FFRAM_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(FFRAM_io_banks_63_wdata_bits)
  );
  assign writeEn = io_in_valid & io_in_ready; // @[FIFO.scala 30:29:@43068.4]
  assign readEn = io_out_valid & io_out_ready; // @[FIFO.scala 31:29:@43069.4]
  assign ptrMatch = enqCounter_io_out == deqCounter_io_out; // @[FIFO.scala 44:36:@43091.4]
  assign _T_824 = maybeFull == 1'h0; // @[FIFO.scala 45:27:@43092.4]
  assign empty = ptrMatch & _T_824; // @[FIFO.scala 45:24:@43093.4]
  assign full = ptrMatch & maybeFull; // @[FIFO.scala 46:23:@43094.4]
  assign _T_1657 = writeEn != readEn; // @[FIFO.scala 83:17:@44261.4]
  assign _GEN_64 = _T_1657 ? writeEn : maybeFull; // @[FIFO.scala 83:29:@44262.4]
  assign io_in_ready = full == 1'h0; // @[FIFO.scala 88:15:@44268.4]
  assign io_out_valid = empty == 1'h0; // @[FIFO.scala 87:16:@44266.4]
  assign io_out_bits = FFRAM_io_rdata; // @[FIFO.scala 56:17:@43300.4]
  assign enqCounter_clock = clock; // @[:@43071.4]
  assign enqCounter_reset = reset; // @[:@43072.4]
  assign enqCounter_io_enable = io_in_valid & io_in_ready; // @[FIFO.scala 36:24:@43078.4]
  assign deqCounter_clock = clock; // @[:@43081.4]
  assign deqCounter_reset = reset; // @[:@43082.4]
  assign deqCounter_io_enable = io_out_valid & io_out_ready; // @[FIFO.scala 40:24:@43088.4]
  assign FFRAM_clock = clock; // @[:@43096.4]
  assign FFRAM_reset = reset; // @[:@43097.4]
  assign FFRAM_io_raddr = deqCounter_io_out; // @[FIFO.scala 52:16:@43296.4]
  assign FFRAM_io_wen = io_in_valid & io_in_ready; // @[FIFO.scala 53:14:@43297.4]
  assign FFRAM_io_waddr = enqCounter_io_out; // @[FIFO.scala 54:16:@43298.4]
  assign FFRAM_io_wdata = io_in_bits; // @[FIFO.scala 55:16:@43299.4]
  assign FFRAM_io_banks_0_wdata_valid = io_banks_0_wdata_valid; // @[FIFO.scala 59:15:@43302.4]
  assign FFRAM_io_banks_0_wdata_bits = io_banks_0_wdata_bits; // @[FIFO.scala 59:15:@43301.4]
  assign FFRAM_io_banks_1_wdata_valid = io_banks_1_wdata_valid; // @[FIFO.scala 59:15:@43305.4]
  assign FFRAM_io_banks_1_wdata_bits = io_banks_1_wdata_bits; // @[FIFO.scala 59:15:@43304.4]
  assign FFRAM_io_banks_2_wdata_valid = io_banks_2_wdata_valid; // @[FIFO.scala 59:15:@43308.4]
  assign FFRAM_io_banks_2_wdata_bits = io_banks_2_wdata_bits; // @[FIFO.scala 59:15:@43307.4]
  assign FFRAM_io_banks_3_wdata_valid = io_banks_3_wdata_valid; // @[FIFO.scala 59:15:@43311.4]
  assign FFRAM_io_banks_3_wdata_bits = io_banks_3_wdata_bits; // @[FIFO.scala 59:15:@43310.4]
  assign FFRAM_io_banks_4_wdata_valid = io_banks_4_wdata_valid; // @[FIFO.scala 59:15:@43314.4]
  assign FFRAM_io_banks_4_wdata_bits = io_banks_4_wdata_bits; // @[FIFO.scala 59:15:@43313.4]
  assign FFRAM_io_banks_5_wdata_valid = io_banks_5_wdata_valid; // @[FIFO.scala 59:15:@43317.4]
  assign FFRAM_io_banks_5_wdata_bits = io_banks_5_wdata_bits; // @[FIFO.scala 59:15:@43316.4]
  assign FFRAM_io_banks_6_wdata_valid = io_banks_6_wdata_valid; // @[FIFO.scala 59:15:@43320.4]
  assign FFRAM_io_banks_6_wdata_bits = io_banks_6_wdata_bits; // @[FIFO.scala 59:15:@43319.4]
  assign FFRAM_io_banks_7_wdata_valid = io_banks_7_wdata_valid; // @[FIFO.scala 59:15:@43323.4]
  assign FFRAM_io_banks_7_wdata_bits = io_banks_7_wdata_bits; // @[FIFO.scala 59:15:@43322.4]
  assign FFRAM_io_banks_8_wdata_valid = io_banks_8_wdata_valid; // @[FIFO.scala 59:15:@43326.4]
  assign FFRAM_io_banks_8_wdata_bits = io_banks_8_wdata_bits; // @[FIFO.scala 59:15:@43325.4]
  assign FFRAM_io_banks_9_wdata_valid = io_banks_9_wdata_valid; // @[FIFO.scala 59:15:@43329.4]
  assign FFRAM_io_banks_9_wdata_bits = io_banks_9_wdata_bits; // @[FIFO.scala 59:15:@43328.4]
  assign FFRAM_io_banks_10_wdata_valid = io_banks_10_wdata_valid; // @[FIFO.scala 59:15:@43332.4]
  assign FFRAM_io_banks_10_wdata_bits = io_banks_10_wdata_bits; // @[FIFO.scala 59:15:@43331.4]
  assign FFRAM_io_banks_11_wdata_valid = io_banks_11_wdata_valid; // @[FIFO.scala 59:15:@43335.4]
  assign FFRAM_io_banks_11_wdata_bits = io_banks_11_wdata_bits; // @[FIFO.scala 59:15:@43334.4]
  assign FFRAM_io_banks_12_wdata_valid = io_banks_12_wdata_valid; // @[FIFO.scala 59:15:@43338.4]
  assign FFRAM_io_banks_12_wdata_bits = io_banks_12_wdata_bits; // @[FIFO.scala 59:15:@43337.4]
  assign FFRAM_io_banks_13_wdata_valid = io_banks_13_wdata_valid; // @[FIFO.scala 59:15:@43341.4]
  assign FFRAM_io_banks_13_wdata_bits = io_banks_13_wdata_bits; // @[FIFO.scala 59:15:@43340.4]
  assign FFRAM_io_banks_14_wdata_valid = io_banks_14_wdata_valid; // @[FIFO.scala 59:15:@43344.4]
  assign FFRAM_io_banks_14_wdata_bits = io_banks_14_wdata_bits; // @[FIFO.scala 59:15:@43343.4]
  assign FFRAM_io_banks_15_wdata_valid = io_banks_15_wdata_valid; // @[FIFO.scala 59:15:@43347.4]
  assign FFRAM_io_banks_15_wdata_bits = io_banks_15_wdata_bits; // @[FIFO.scala 59:15:@43346.4]
  assign FFRAM_io_banks_16_wdata_valid = io_banks_16_wdata_valid; // @[FIFO.scala 59:15:@43350.4]
  assign FFRAM_io_banks_16_wdata_bits = io_banks_16_wdata_bits; // @[FIFO.scala 59:15:@43349.4]
  assign FFRAM_io_banks_17_wdata_valid = io_banks_17_wdata_valid; // @[FIFO.scala 59:15:@43353.4]
  assign FFRAM_io_banks_17_wdata_bits = io_banks_17_wdata_bits; // @[FIFO.scala 59:15:@43352.4]
  assign FFRAM_io_banks_18_wdata_valid = io_banks_18_wdata_valid; // @[FIFO.scala 59:15:@43356.4]
  assign FFRAM_io_banks_18_wdata_bits = io_banks_18_wdata_bits; // @[FIFO.scala 59:15:@43355.4]
  assign FFRAM_io_banks_19_wdata_valid = io_banks_19_wdata_valid; // @[FIFO.scala 59:15:@43359.4]
  assign FFRAM_io_banks_19_wdata_bits = io_banks_19_wdata_bits; // @[FIFO.scala 59:15:@43358.4]
  assign FFRAM_io_banks_20_wdata_valid = io_banks_20_wdata_valid; // @[FIFO.scala 59:15:@43362.4]
  assign FFRAM_io_banks_20_wdata_bits = io_banks_20_wdata_bits; // @[FIFO.scala 59:15:@43361.4]
  assign FFRAM_io_banks_21_wdata_valid = io_banks_21_wdata_valid; // @[FIFO.scala 59:15:@43365.4]
  assign FFRAM_io_banks_21_wdata_bits = io_banks_21_wdata_bits; // @[FIFO.scala 59:15:@43364.4]
  assign FFRAM_io_banks_22_wdata_valid = io_banks_22_wdata_valid; // @[FIFO.scala 59:15:@43368.4]
  assign FFRAM_io_banks_22_wdata_bits = io_banks_22_wdata_bits; // @[FIFO.scala 59:15:@43367.4]
  assign FFRAM_io_banks_23_wdata_valid = io_banks_23_wdata_valid; // @[FIFO.scala 59:15:@43371.4]
  assign FFRAM_io_banks_23_wdata_bits = io_banks_23_wdata_bits; // @[FIFO.scala 59:15:@43370.4]
  assign FFRAM_io_banks_24_wdata_valid = io_banks_24_wdata_valid; // @[FIFO.scala 59:15:@43374.4]
  assign FFRAM_io_banks_24_wdata_bits = io_banks_24_wdata_bits; // @[FIFO.scala 59:15:@43373.4]
  assign FFRAM_io_banks_25_wdata_valid = io_banks_25_wdata_valid; // @[FIFO.scala 59:15:@43377.4]
  assign FFRAM_io_banks_25_wdata_bits = io_banks_25_wdata_bits; // @[FIFO.scala 59:15:@43376.4]
  assign FFRAM_io_banks_26_wdata_valid = io_banks_26_wdata_valid; // @[FIFO.scala 59:15:@43380.4]
  assign FFRAM_io_banks_26_wdata_bits = io_banks_26_wdata_bits; // @[FIFO.scala 59:15:@43379.4]
  assign FFRAM_io_banks_27_wdata_valid = io_banks_27_wdata_valid; // @[FIFO.scala 59:15:@43383.4]
  assign FFRAM_io_banks_27_wdata_bits = io_banks_27_wdata_bits; // @[FIFO.scala 59:15:@43382.4]
  assign FFRAM_io_banks_28_wdata_valid = io_banks_28_wdata_valid; // @[FIFO.scala 59:15:@43386.4]
  assign FFRAM_io_banks_28_wdata_bits = io_banks_28_wdata_bits; // @[FIFO.scala 59:15:@43385.4]
  assign FFRAM_io_banks_29_wdata_valid = io_banks_29_wdata_valid; // @[FIFO.scala 59:15:@43389.4]
  assign FFRAM_io_banks_29_wdata_bits = io_banks_29_wdata_bits; // @[FIFO.scala 59:15:@43388.4]
  assign FFRAM_io_banks_30_wdata_valid = io_banks_30_wdata_valid; // @[FIFO.scala 59:15:@43392.4]
  assign FFRAM_io_banks_30_wdata_bits = io_banks_30_wdata_bits; // @[FIFO.scala 59:15:@43391.4]
  assign FFRAM_io_banks_31_wdata_valid = io_banks_31_wdata_valid; // @[FIFO.scala 59:15:@43395.4]
  assign FFRAM_io_banks_31_wdata_bits = io_banks_31_wdata_bits; // @[FIFO.scala 59:15:@43394.4]
  assign FFRAM_io_banks_32_wdata_valid = io_banks_32_wdata_valid; // @[FIFO.scala 59:15:@43398.4]
  assign FFRAM_io_banks_32_wdata_bits = io_banks_32_wdata_bits; // @[FIFO.scala 59:15:@43397.4]
  assign FFRAM_io_banks_33_wdata_valid = io_banks_33_wdata_valid; // @[FIFO.scala 59:15:@43401.4]
  assign FFRAM_io_banks_33_wdata_bits = io_banks_33_wdata_bits; // @[FIFO.scala 59:15:@43400.4]
  assign FFRAM_io_banks_34_wdata_valid = io_banks_34_wdata_valid; // @[FIFO.scala 59:15:@43404.4]
  assign FFRAM_io_banks_34_wdata_bits = io_banks_34_wdata_bits; // @[FIFO.scala 59:15:@43403.4]
  assign FFRAM_io_banks_35_wdata_valid = io_banks_35_wdata_valid; // @[FIFO.scala 59:15:@43407.4]
  assign FFRAM_io_banks_35_wdata_bits = io_banks_35_wdata_bits; // @[FIFO.scala 59:15:@43406.4]
  assign FFRAM_io_banks_36_wdata_valid = io_banks_36_wdata_valid; // @[FIFO.scala 59:15:@43410.4]
  assign FFRAM_io_banks_36_wdata_bits = io_banks_36_wdata_bits; // @[FIFO.scala 59:15:@43409.4]
  assign FFRAM_io_banks_37_wdata_valid = io_banks_37_wdata_valid; // @[FIFO.scala 59:15:@43413.4]
  assign FFRAM_io_banks_37_wdata_bits = io_banks_37_wdata_bits; // @[FIFO.scala 59:15:@43412.4]
  assign FFRAM_io_banks_38_wdata_valid = io_banks_38_wdata_valid; // @[FIFO.scala 59:15:@43416.4]
  assign FFRAM_io_banks_38_wdata_bits = io_banks_38_wdata_bits; // @[FIFO.scala 59:15:@43415.4]
  assign FFRAM_io_banks_39_wdata_valid = io_banks_39_wdata_valid; // @[FIFO.scala 59:15:@43419.4]
  assign FFRAM_io_banks_39_wdata_bits = io_banks_39_wdata_bits; // @[FIFO.scala 59:15:@43418.4]
  assign FFRAM_io_banks_40_wdata_valid = io_banks_40_wdata_valid; // @[FIFO.scala 59:15:@43422.4]
  assign FFRAM_io_banks_40_wdata_bits = io_banks_40_wdata_bits; // @[FIFO.scala 59:15:@43421.4]
  assign FFRAM_io_banks_41_wdata_valid = io_banks_41_wdata_valid; // @[FIFO.scala 59:15:@43425.4]
  assign FFRAM_io_banks_41_wdata_bits = io_banks_41_wdata_bits; // @[FIFO.scala 59:15:@43424.4]
  assign FFRAM_io_banks_42_wdata_valid = io_banks_42_wdata_valid; // @[FIFO.scala 59:15:@43428.4]
  assign FFRAM_io_banks_42_wdata_bits = io_banks_42_wdata_bits; // @[FIFO.scala 59:15:@43427.4]
  assign FFRAM_io_banks_43_wdata_valid = io_banks_43_wdata_valid; // @[FIFO.scala 59:15:@43431.4]
  assign FFRAM_io_banks_43_wdata_bits = io_banks_43_wdata_bits; // @[FIFO.scala 59:15:@43430.4]
  assign FFRAM_io_banks_44_wdata_valid = io_banks_44_wdata_valid; // @[FIFO.scala 59:15:@43434.4]
  assign FFRAM_io_banks_44_wdata_bits = io_banks_44_wdata_bits; // @[FIFO.scala 59:15:@43433.4]
  assign FFRAM_io_banks_45_wdata_valid = io_banks_45_wdata_valid; // @[FIFO.scala 59:15:@43437.4]
  assign FFRAM_io_banks_45_wdata_bits = io_banks_45_wdata_bits; // @[FIFO.scala 59:15:@43436.4]
  assign FFRAM_io_banks_46_wdata_valid = io_banks_46_wdata_valid; // @[FIFO.scala 59:15:@43440.4]
  assign FFRAM_io_banks_46_wdata_bits = io_banks_46_wdata_bits; // @[FIFO.scala 59:15:@43439.4]
  assign FFRAM_io_banks_47_wdata_valid = io_banks_47_wdata_valid; // @[FIFO.scala 59:15:@43443.4]
  assign FFRAM_io_banks_47_wdata_bits = io_banks_47_wdata_bits; // @[FIFO.scala 59:15:@43442.4]
  assign FFRAM_io_banks_48_wdata_valid = io_banks_48_wdata_valid; // @[FIFO.scala 59:15:@43446.4]
  assign FFRAM_io_banks_48_wdata_bits = io_banks_48_wdata_bits; // @[FIFO.scala 59:15:@43445.4]
  assign FFRAM_io_banks_49_wdata_valid = io_banks_49_wdata_valid; // @[FIFO.scala 59:15:@43449.4]
  assign FFRAM_io_banks_49_wdata_bits = io_banks_49_wdata_bits; // @[FIFO.scala 59:15:@43448.4]
  assign FFRAM_io_banks_50_wdata_valid = io_banks_50_wdata_valid; // @[FIFO.scala 59:15:@43452.4]
  assign FFRAM_io_banks_50_wdata_bits = io_banks_50_wdata_bits; // @[FIFO.scala 59:15:@43451.4]
  assign FFRAM_io_banks_51_wdata_valid = io_banks_51_wdata_valid; // @[FIFO.scala 59:15:@43455.4]
  assign FFRAM_io_banks_51_wdata_bits = io_banks_51_wdata_bits; // @[FIFO.scala 59:15:@43454.4]
  assign FFRAM_io_banks_52_wdata_valid = io_banks_52_wdata_valid; // @[FIFO.scala 59:15:@43458.4]
  assign FFRAM_io_banks_52_wdata_bits = io_banks_52_wdata_bits; // @[FIFO.scala 59:15:@43457.4]
  assign FFRAM_io_banks_53_wdata_valid = io_banks_53_wdata_valid; // @[FIFO.scala 59:15:@43461.4]
  assign FFRAM_io_banks_53_wdata_bits = io_banks_53_wdata_bits; // @[FIFO.scala 59:15:@43460.4]
  assign FFRAM_io_banks_54_wdata_valid = io_banks_54_wdata_valid; // @[FIFO.scala 59:15:@43464.4]
  assign FFRAM_io_banks_54_wdata_bits = io_banks_54_wdata_bits; // @[FIFO.scala 59:15:@43463.4]
  assign FFRAM_io_banks_55_wdata_valid = io_banks_55_wdata_valid; // @[FIFO.scala 59:15:@43467.4]
  assign FFRAM_io_banks_55_wdata_bits = io_banks_55_wdata_bits; // @[FIFO.scala 59:15:@43466.4]
  assign FFRAM_io_banks_56_wdata_valid = io_banks_56_wdata_valid; // @[FIFO.scala 59:15:@43470.4]
  assign FFRAM_io_banks_56_wdata_bits = io_banks_56_wdata_bits; // @[FIFO.scala 59:15:@43469.4]
  assign FFRAM_io_banks_57_wdata_valid = io_banks_57_wdata_valid; // @[FIFO.scala 59:15:@43473.4]
  assign FFRAM_io_banks_57_wdata_bits = io_banks_57_wdata_bits; // @[FIFO.scala 59:15:@43472.4]
  assign FFRAM_io_banks_58_wdata_valid = io_banks_58_wdata_valid; // @[FIFO.scala 59:15:@43476.4]
  assign FFRAM_io_banks_58_wdata_bits = io_banks_58_wdata_bits; // @[FIFO.scala 59:15:@43475.4]
  assign FFRAM_io_banks_59_wdata_valid = io_banks_59_wdata_valid; // @[FIFO.scala 59:15:@43479.4]
  assign FFRAM_io_banks_59_wdata_bits = io_banks_59_wdata_bits; // @[FIFO.scala 59:15:@43478.4]
  assign FFRAM_io_banks_60_wdata_valid = io_banks_60_wdata_valid; // @[FIFO.scala 59:15:@43482.4]
  assign FFRAM_io_banks_60_wdata_bits = io_banks_60_wdata_bits; // @[FIFO.scala 59:15:@43481.4]
  assign FFRAM_io_banks_61_wdata_valid = io_banks_61_wdata_valid; // @[FIFO.scala 59:15:@43485.4]
  assign FFRAM_io_banks_61_wdata_bits = io_banks_61_wdata_bits; // @[FIFO.scala 59:15:@43484.4]
  assign FFRAM_io_banks_62_wdata_valid = io_banks_62_wdata_valid; // @[FIFO.scala 59:15:@43488.4]
  assign FFRAM_io_banks_62_wdata_bits = io_banks_62_wdata_bits; // @[FIFO.scala 59:15:@43487.4]
  assign FFRAM_io_banks_63_wdata_valid = io_banks_63_wdata_valid; // @[FIFO.scala 59:15:@43491.4]
  assign FFRAM_io_banks_63_wdata_bits = io_banks_63_wdata_bits; // @[FIFO.scala 59:15:@43490.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  maybeFull = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      maybeFull <= 1'h0;
    end else begin
      if (_T_1657) begin
        maybeFull <= writeEn;
      end
    end
  end
endmodule
module StreamControllerStore( // @[:@44270.2]
  input         clock, // @[:@44271.4]
  input         reset, // @[:@44272.4]
  input         io_dram_cmd_ready, // @[:@44273.4]
  output        io_dram_cmd_valid, // @[:@44273.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@44273.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@44273.4]
  input         io_dram_wdata_ready, // @[:@44273.4]
  output        io_dram_wdata_valid, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@44273.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@44273.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@44273.4]
  output        io_dram_wresp_ready, // @[:@44273.4]
  input         io_dram_wresp_valid, // @[:@44273.4]
  output        io_store_cmd_ready, // @[:@44273.4]
  input         io_store_cmd_valid, // @[:@44273.4]
  input  [63:0] io_store_cmd_bits_addr, // @[:@44273.4]
  input  [31:0] io_store_cmd_bits_size, // @[:@44273.4]
  output        io_store_data_ready, // @[:@44273.4]
  input         io_store_data_valid, // @[:@44273.4]
  input  [31:0] io_store_data_bits_wdata_0, // @[:@44273.4]
  input         io_store_data_bits_wstrb, // @[:@44273.4]
  input         io_store_wresp_ready, // @[:@44273.4]
  output        io_store_wresp_valid, // @[:@44273.4]
  output        io_store_wresp_bits // @[:@44273.4]
);
  wire  cmd_clock; // @[StreamController.scala 75:19:@44398.4]
  wire  cmd_reset; // @[StreamController.scala 75:19:@44398.4]
  wire  cmd_io_in_ready; // @[StreamController.scala 75:19:@44398.4]
  wire  cmd_io_in_valid; // @[StreamController.scala 75:19:@44398.4]
  wire [63:0] cmd_io_in_bits_addr; // @[StreamController.scala 75:19:@44398.4]
  wire [31:0] cmd_io_in_bits_size; // @[StreamController.scala 75:19:@44398.4]
  wire  cmd_io_out_ready; // @[StreamController.scala 75:19:@44398.4]
  wire  cmd_io_out_valid; // @[StreamController.scala 75:19:@44398.4]
  wire [63:0] cmd_io_out_bits_addr; // @[StreamController.scala 75:19:@44398.4]
  wire [31:0] cmd_io_out_bits_size; // @[StreamController.scala 75:19:@44398.4]
  wire  wdata_clock; // @[StreamController.scala 88:21:@44804.4]
  wire  wdata_reset; // @[StreamController.scala 88:21:@44804.4]
  wire  wdata_io_in_ready; // @[StreamController.scala 88:21:@44804.4]
  wire  wdata_io_in_valid; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_in_bits_data_0; // @[StreamController.scala 88:21:@44804.4]
  wire  wdata_io_in_bits_strobe; // @[StreamController.scala 88:21:@44804.4]
  wire  wdata_io_out_ready; // @[StreamController.scala 88:21:@44804.4]
  wire  wdata_io_out_valid; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_0; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_1; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_2; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_3; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_4; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_5; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_6; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_7; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_8; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_9; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_10; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_11; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_12; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_13; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_14; // @[StreamController.scala 88:21:@44804.4]
  wire [31:0] wdata_io_out_bits_data_15; // @[StreamController.scala 88:21:@44804.4]
  wire [63:0] wdata_io_out_bits_strobe; // @[StreamController.scala 88:21:@44804.4]
  wire  wresp_clock; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_reset; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_in_ready; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_in_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_in_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_out_ready; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_out_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_out_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_0_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_0_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_1_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_1_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_2_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_2_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_3_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_3_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_4_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_4_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_5_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_5_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_6_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_6_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_7_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_7_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_8_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_8_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_9_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_9_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_10_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_10_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_11_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_11_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_12_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_12_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_13_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_13_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_14_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_14_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_15_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_15_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_16_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_16_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_17_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_17_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_18_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_18_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_19_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_19_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_20_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_20_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_21_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_21_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_22_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_22_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_23_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_23_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_24_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_24_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_25_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_25_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_26_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_26_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_27_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_27_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_28_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_28_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_29_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_29_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_30_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_30_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_31_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_31_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_32_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_32_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_33_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_33_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_34_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_34_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_35_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_35_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_36_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_36_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_37_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_37_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_38_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_38_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_39_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_39_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_40_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_40_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_41_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_41_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_42_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_42_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_43_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_43_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_44_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_44_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_45_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_45_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_46_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_46_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_47_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_47_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_48_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_48_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_49_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_49_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_50_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_50_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_51_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_51_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_52_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_52_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_53_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_53_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_54_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_54_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_55_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_55_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_56_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_56_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_57_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_57_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_58_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_58_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_59_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_59_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_60_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_60_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_61_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_61_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_62_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_62_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_63_wdata_valid; // @[StreamController.scala 100:21:@45045.4]
  wire  wresp_io_banks_63_wdata_bits; // @[StreamController.scala 100:21:@45045.4]
  wire [25:0] _T_111; // @[StreamController.scala 21:10:@44801.4]
  FIFO cmd ( // @[StreamController.scala 75:19:@44398.4]
    .clock(cmd_clock),
    .reset(cmd_reset),
    .io_in_ready(cmd_io_in_ready),
    .io_in_valid(cmd_io_in_valid),
    .io_in_bits_addr(cmd_io_in_bits_addr),
    .io_in_bits_size(cmd_io_in_bits_size),
    .io_out_ready(cmd_io_out_ready),
    .io_out_valid(cmd_io_out_valid),
    .io_out_bits_addr(cmd_io_out_bits_addr),
    .io_out_bits_size(cmd_io_out_bits_size)
  );
  FIFOWidthConvert wdata ( // @[StreamController.scala 88:21:@44804.4]
    .clock(wdata_clock),
    .reset(wdata_reset),
    .io_in_ready(wdata_io_in_ready),
    .io_in_valid(wdata_io_in_valid),
    .io_in_bits_data_0(wdata_io_in_bits_data_0),
    .io_in_bits_strobe(wdata_io_in_bits_strobe),
    .io_out_ready(wdata_io_out_ready),
    .io_out_valid(wdata_io_out_valid),
    .io_out_bits_data_0(wdata_io_out_bits_data_0),
    .io_out_bits_data_1(wdata_io_out_bits_data_1),
    .io_out_bits_data_2(wdata_io_out_bits_data_2),
    .io_out_bits_data_3(wdata_io_out_bits_data_3),
    .io_out_bits_data_4(wdata_io_out_bits_data_4),
    .io_out_bits_data_5(wdata_io_out_bits_data_5),
    .io_out_bits_data_6(wdata_io_out_bits_data_6),
    .io_out_bits_data_7(wdata_io_out_bits_data_7),
    .io_out_bits_data_8(wdata_io_out_bits_data_8),
    .io_out_bits_data_9(wdata_io_out_bits_data_9),
    .io_out_bits_data_10(wdata_io_out_bits_data_10),
    .io_out_bits_data_11(wdata_io_out_bits_data_11),
    .io_out_bits_data_12(wdata_io_out_bits_data_12),
    .io_out_bits_data_13(wdata_io_out_bits_data_13),
    .io_out_bits_data_14(wdata_io_out_bits_data_14),
    .io_out_bits_data_15(wdata_io_out_bits_data_15),
    .io_out_bits_strobe(wdata_io_out_bits_strobe)
  );
  FIFO_33 wresp ( // @[StreamController.scala 100:21:@45045.4]
    .clock(wresp_clock),
    .reset(wresp_reset),
    .io_in_ready(wresp_io_in_ready),
    .io_in_valid(wresp_io_in_valid),
    .io_in_bits(wresp_io_in_bits),
    .io_out_ready(wresp_io_out_ready),
    .io_out_valid(wresp_io_out_valid),
    .io_out_bits(wresp_io_out_bits),
    .io_banks_0_wdata_valid(wresp_io_banks_0_wdata_valid),
    .io_banks_0_wdata_bits(wresp_io_banks_0_wdata_bits),
    .io_banks_1_wdata_valid(wresp_io_banks_1_wdata_valid),
    .io_banks_1_wdata_bits(wresp_io_banks_1_wdata_bits),
    .io_banks_2_wdata_valid(wresp_io_banks_2_wdata_valid),
    .io_banks_2_wdata_bits(wresp_io_banks_2_wdata_bits),
    .io_banks_3_wdata_valid(wresp_io_banks_3_wdata_valid),
    .io_banks_3_wdata_bits(wresp_io_banks_3_wdata_bits),
    .io_banks_4_wdata_valid(wresp_io_banks_4_wdata_valid),
    .io_banks_4_wdata_bits(wresp_io_banks_4_wdata_bits),
    .io_banks_5_wdata_valid(wresp_io_banks_5_wdata_valid),
    .io_banks_5_wdata_bits(wresp_io_banks_5_wdata_bits),
    .io_banks_6_wdata_valid(wresp_io_banks_6_wdata_valid),
    .io_banks_6_wdata_bits(wresp_io_banks_6_wdata_bits),
    .io_banks_7_wdata_valid(wresp_io_banks_7_wdata_valid),
    .io_banks_7_wdata_bits(wresp_io_banks_7_wdata_bits),
    .io_banks_8_wdata_valid(wresp_io_banks_8_wdata_valid),
    .io_banks_8_wdata_bits(wresp_io_banks_8_wdata_bits),
    .io_banks_9_wdata_valid(wresp_io_banks_9_wdata_valid),
    .io_banks_9_wdata_bits(wresp_io_banks_9_wdata_bits),
    .io_banks_10_wdata_valid(wresp_io_banks_10_wdata_valid),
    .io_banks_10_wdata_bits(wresp_io_banks_10_wdata_bits),
    .io_banks_11_wdata_valid(wresp_io_banks_11_wdata_valid),
    .io_banks_11_wdata_bits(wresp_io_banks_11_wdata_bits),
    .io_banks_12_wdata_valid(wresp_io_banks_12_wdata_valid),
    .io_banks_12_wdata_bits(wresp_io_banks_12_wdata_bits),
    .io_banks_13_wdata_valid(wresp_io_banks_13_wdata_valid),
    .io_banks_13_wdata_bits(wresp_io_banks_13_wdata_bits),
    .io_banks_14_wdata_valid(wresp_io_banks_14_wdata_valid),
    .io_banks_14_wdata_bits(wresp_io_banks_14_wdata_bits),
    .io_banks_15_wdata_valid(wresp_io_banks_15_wdata_valid),
    .io_banks_15_wdata_bits(wresp_io_banks_15_wdata_bits),
    .io_banks_16_wdata_valid(wresp_io_banks_16_wdata_valid),
    .io_banks_16_wdata_bits(wresp_io_banks_16_wdata_bits),
    .io_banks_17_wdata_valid(wresp_io_banks_17_wdata_valid),
    .io_banks_17_wdata_bits(wresp_io_banks_17_wdata_bits),
    .io_banks_18_wdata_valid(wresp_io_banks_18_wdata_valid),
    .io_banks_18_wdata_bits(wresp_io_banks_18_wdata_bits),
    .io_banks_19_wdata_valid(wresp_io_banks_19_wdata_valid),
    .io_banks_19_wdata_bits(wresp_io_banks_19_wdata_bits),
    .io_banks_20_wdata_valid(wresp_io_banks_20_wdata_valid),
    .io_banks_20_wdata_bits(wresp_io_banks_20_wdata_bits),
    .io_banks_21_wdata_valid(wresp_io_banks_21_wdata_valid),
    .io_banks_21_wdata_bits(wresp_io_banks_21_wdata_bits),
    .io_banks_22_wdata_valid(wresp_io_banks_22_wdata_valid),
    .io_banks_22_wdata_bits(wresp_io_banks_22_wdata_bits),
    .io_banks_23_wdata_valid(wresp_io_banks_23_wdata_valid),
    .io_banks_23_wdata_bits(wresp_io_banks_23_wdata_bits),
    .io_banks_24_wdata_valid(wresp_io_banks_24_wdata_valid),
    .io_banks_24_wdata_bits(wresp_io_banks_24_wdata_bits),
    .io_banks_25_wdata_valid(wresp_io_banks_25_wdata_valid),
    .io_banks_25_wdata_bits(wresp_io_banks_25_wdata_bits),
    .io_banks_26_wdata_valid(wresp_io_banks_26_wdata_valid),
    .io_banks_26_wdata_bits(wresp_io_banks_26_wdata_bits),
    .io_banks_27_wdata_valid(wresp_io_banks_27_wdata_valid),
    .io_banks_27_wdata_bits(wresp_io_banks_27_wdata_bits),
    .io_banks_28_wdata_valid(wresp_io_banks_28_wdata_valid),
    .io_banks_28_wdata_bits(wresp_io_banks_28_wdata_bits),
    .io_banks_29_wdata_valid(wresp_io_banks_29_wdata_valid),
    .io_banks_29_wdata_bits(wresp_io_banks_29_wdata_bits),
    .io_banks_30_wdata_valid(wresp_io_banks_30_wdata_valid),
    .io_banks_30_wdata_bits(wresp_io_banks_30_wdata_bits),
    .io_banks_31_wdata_valid(wresp_io_banks_31_wdata_valid),
    .io_banks_31_wdata_bits(wresp_io_banks_31_wdata_bits),
    .io_banks_32_wdata_valid(wresp_io_banks_32_wdata_valid),
    .io_banks_32_wdata_bits(wresp_io_banks_32_wdata_bits),
    .io_banks_33_wdata_valid(wresp_io_banks_33_wdata_valid),
    .io_banks_33_wdata_bits(wresp_io_banks_33_wdata_bits),
    .io_banks_34_wdata_valid(wresp_io_banks_34_wdata_valid),
    .io_banks_34_wdata_bits(wresp_io_banks_34_wdata_bits),
    .io_banks_35_wdata_valid(wresp_io_banks_35_wdata_valid),
    .io_banks_35_wdata_bits(wresp_io_banks_35_wdata_bits),
    .io_banks_36_wdata_valid(wresp_io_banks_36_wdata_valid),
    .io_banks_36_wdata_bits(wresp_io_banks_36_wdata_bits),
    .io_banks_37_wdata_valid(wresp_io_banks_37_wdata_valid),
    .io_banks_37_wdata_bits(wresp_io_banks_37_wdata_bits),
    .io_banks_38_wdata_valid(wresp_io_banks_38_wdata_valid),
    .io_banks_38_wdata_bits(wresp_io_banks_38_wdata_bits),
    .io_banks_39_wdata_valid(wresp_io_banks_39_wdata_valid),
    .io_banks_39_wdata_bits(wresp_io_banks_39_wdata_bits),
    .io_banks_40_wdata_valid(wresp_io_banks_40_wdata_valid),
    .io_banks_40_wdata_bits(wresp_io_banks_40_wdata_bits),
    .io_banks_41_wdata_valid(wresp_io_banks_41_wdata_valid),
    .io_banks_41_wdata_bits(wresp_io_banks_41_wdata_bits),
    .io_banks_42_wdata_valid(wresp_io_banks_42_wdata_valid),
    .io_banks_42_wdata_bits(wresp_io_banks_42_wdata_bits),
    .io_banks_43_wdata_valid(wresp_io_banks_43_wdata_valid),
    .io_banks_43_wdata_bits(wresp_io_banks_43_wdata_bits),
    .io_banks_44_wdata_valid(wresp_io_banks_44_wdata_valid),
    .io_banks_44_wdata_bits(wresp_io_banks_44_wdata_bits),
    .io_banks_45_wdata_valid(wresp_io_banks_45_wdata_valid),
    .io_banks_45_wdata_bits(wresp_io_banks_45_wdata_bits),
    .io_banks_46_wdata_valid(wresp_io_banks_46_wdata_valid),
    .io_banks_46_wdata_bits(wresp_io_banks_46_wdata_bits),
    .io_banks_47_wdata_valid(wresp_io_banks_47_wdata_valid),
    .io_banks_47_wdata_bits(wresp_io_banks_47_wdata_bits),
    .io_banks_48_wdata_valid(wresp_io_banks_48_wdata_valid),
    .io_banks_48_wdata_bits(wresp_io_banks_48_wdata_bits),
    .io_banks_49_wdata_valid(wresp_io_banks_49_wdata_valid),
    .io_banks_49_wdata_bits(wresp_io_banks_49_wdata_bits),
    .io_banks_50_wdata_valid(wresp_io_banks_50_wdata_valid),
    .io_banks_50_wdata_bits(wresp_io_banks_50_wdata_bits),
    .io_banks_51_wdata_valid(wresp_io_banks_51_wdata_valid),
    .io_banks_51_wdata_bits(wresp_io_banks_51_wdata_bits),
    .io_banks_52_wdata_valid(wresp_io_banks_52_wdata_valid),
    .io_banks_52_wdata_bits(wresp_io_banks_52_wdata_bits),
    .io_banks_53_wdata_valid(wresp_io_banks_53_wdata_valid),
    .io_banks_53_wdata_bits(wresp_io_banks_53_wdata_bits),
    .io_banks_54_wdata_valid(wresp_io_banks_54_wdata_valid),
    .io_banks_54_wdata_bits(wresp_io_banks_54_wdata_bits),
    .io_banks_55_wdata_valid(wresp_io_banks_55_wdata_valid),
    .io_banks_55_wdata_bits(wresp_io_banks_55_wdata_bits),
    .io_banks_56_wdata_valid(wresp_io_banks_56_wdata_valid),
    .io_banks_56_wdata_bits(wresp_io_banks_56_wdata_bits),
    .io_banks_57_wdata_valid(wresp_io_banks_57_wdata_valid),
    .io_banks_57_wdata_bits(wresp_io_banks_57_wdata_bits),
    .io_banks_58_wdata_valid(wresp_io_banks_58_wdata_valid),
    .io_banks_58_wdata_bits(wresp_io_banks_58_wdata_bits),
    .io_banks_59_wdata_valid(wresp_io_banks_59_wdata_valid),
    .io_banks_59_wdata_bits(wresp_io_banks_59_wdata_bits),
    .io_banks_60_wdata_valid(wresp_io_banks_60_wdata_valid),
    .io_banks_60_wdata_bits(wresp_io_banks_60_wdata_bits),
    .io_banks_61_wdata_valid(wresp_io_banks_61_wdata_valid),
    .io_banks_61_wdata_bits(wresp_io_banks_61_wdata_bits),
    .io_banks_62_wdata_valid(wresp_io_banks_62_wdata_valid),
    .io_banks_62_wdata_bits(wresp_io_banks_62_wdata_bits),
    .io_banks_63_wdata_valid(wresp_io_banks_63_wdata_valid),
    .io_banks_63_wdata_bits(wresp_io_banks_63_wdata_bits)
  );
  assign _T_111 = cmd_io_out_bits_size[31:6]; // @[StreamController.scala 21:10:@44801.4]
  assign io_dram_cmd_valid = cmd_io_out_valid; // @[StreamController.scala 81:21:@44798.4]
  assign io_dram_cmd_bits_addr = cmd_io_out_bits_addr; // @[StreamController.scala 83:25:@44799.4]
  assign io_dram_cmd_bits_size = {{6'd0}, _T_111}; // @[StreamController.scala 85:25:@44802.4]
  assign io_dram_wdata_valid = wdata_io_out_valid; // @[StreamController.scala 95:23:@44834.4]
  assign io_dram_wdata_bits_wdata_0 = wdata_io_out_bits_data_0; // @[StreamController.scala 96:28:@44835.4]
  assign io_dram_wdata_bits_wdata_1 = wdata_io_out_bits_data_1; // @[StreamController.scala 96:28:@44836.4]
  assign io_dram_wdata_bits_wdata_2 = wdata_io_out_bits_data_2; // @[StreamController.scala 96:28:@44837.4]
  assign io_dram_wdata_bits_wdata_3 = wdata_io_out_bits_data_3; // @[StreamController.scala 96:28:@44838.4]
  assign io_dram_wdata_bits_wdata_4 = wdata_io_out_bits_data_4; // @[StreamController.scala 96:28:@44839.4]
  assign io_dram_wdata_bits_wdata_5 = wdata_io_out_bits_data_5; // @[StreamController.scala 96:28:@44840.4]
  assign io_dram_wdata_bits_wdata_6 = wdata_io_out_bits_data_6; // @[StreamController.scala 96:28:@44841.4]
  assign io_dram_wdata_bits_wdata_7 = wdata_io_out_bits_data_7; // @[StreamController.scala 96:28:@44842.4]
  assign io_dram_wdata_bits_wdata_8 = wdata_io_out_bits_data_8; // @[StreamController.scala 96:28:@44843.4]
  assign io_dram_wdata_bits_wdata_9 = wdata_io_out_bits_data_9; // @[StreamController.scala 96:28:@44844.4]
  assign io_dram_wdata_bits_wdata_10 = wdata_io_out_bits_data_10; // @[StreamController.scala 96:28:@44845.4]
  assign io_dram_wdata_bits_wdata_11 = wdata_io_out_bits_data_11; // @[StreamController.scala 96:28:@44846.4]
  assign io_dram_wdata_bits_wdata_12 = wdata_io_out_bits_data_12; // @[StreamController.scala 96:28:@44847.4]
  assign io_dram_wdata_bits_wdata_13 = wdata_io_out_bits_data_13; // @[StreamController.scala 96:28:@44848.4]
  assign io_dram_wdata_bits_wdata_14 = wdata_io_out_bits_data_14; // @[StreamController.scala 96:28:@44849.4]
  assign io_dram_wdata_bits_wdata_15 = wdata_io_out_bits_data_15; // @[StreamController.scala 96:28:@44850.4]
  assign io_dram_wdata_bits_wstrb_0 = wdata_io_out_bits_strobe[63]; // @[StreamController.scala 97:28:@44980.4]
  assign io_dram_wdata_bits_wstrb_1 = wdata_io_out_bits_strobe[62]; // @[StreamController.scala 97:28:@44981.4]
  assign io_dram_wdata_bits_wstrb_2 = wdata_io_out_bits_strobe[61]; // @[StreamController.scala 97:28:@44982.4]
  assign io_dram_wdata_bits_wstrb_3 = wdata_io_out_bits_strobe[60]; // @[StreamController.scala 97:28:@44983.4]
  assign io_dram_wdata_bits_wstrb_4 = wdata_io_out_bits_strobe[59]; // @[StreamController.scala 97:28:@44984.4]
  assign io_dram_wdata_bits_wstrb_5 = wdata_io_out_bits_strobe[58]; // @[StreamController.scala 97:28:@44985.4]
  assign io_dram_wdata_bits_wstrb_6 = wdata_io_out_bits_strobe[57]; // @[StreamController.scala 97:28:@44986.4]
  assign io_dram_wdata_bits_wstrb_7 = wdata_io_out_bits_strobe[56]; // @[StreamController.scala 97:28:@44987.4]
  assign io_dram_wdata_bits_wstrb_8 = wdata_io_out_bits_strobe[55]; // @[StreamController.scala 97:28:@44988.4]
  assign io_dram_wdata_bits_wstrb_9 = wdata_io_out_bits_strobe[54]; // @[StreamController.scala 97:28:@44989.4]
  assign io_dram_wdata_bits_wstrb_10 = wdata_io_out_bits_strobe[53]; // @[StreamController.scala 97:28:@44990.4]
  assign io_dram_wdata_bits_wstrb_11 = wdata_io_out_bits_strobe[52]; // @[StreamController.scala 97:28:@44991.4]
  assign io_dram_wdata_bits_wstrb_12 = wdata_io_out_bits_strobe[51]; // @[StreamController.scala 97:28:@44992.4]
  assign io_dram_wdata_bits_wstrb_13 = wdata_io_out_bits_strobe[50]; // @[StreamController.scala 97:28:@44993.4]
  assign io_dram_wdata_bits_wstrb_14 = wdata_io_out_bits_strobe[49]; // @[StreamController.scala 97:28:@44994.4]
  assign io_dram_wdata_bits_wstrb_15 = wdata_io_out_bits_strobe[48]; // @[StreamController.scala 97:28:@44995.4]
  assign io_dram_wdata_bits_wstrb_16 = wdata_io_out_bits_strobe[47]; // @[StreamController.scala 97:28:@44996.4]
  assign io_dram_wdata_bits_wstrb_17 = wdata_io_out_bits_strobe[46]; // @[StreamController.scala 97:28:@44997.4]
  assign io_dram_wdata_bits_wstrb_18 = wdata_io_out_bits_strobe[45]; // @[StreamController.scala 97:28:@44998.4]
  assign io_dram_wdata_bits_wstrb_19 = wdata_io_out_bits_strobe[44]; // @[StreamController.scala 97:28:@44999.4]
  assign io_dram_wdata_bits_wstrb_20 = wdata_io_out_bits_strobe[43]; // @[StreamController.scala 97:28:@45000.4]
  assign io_dram_wdata_bits_wstrb_21 = wdata_io_out_bits_strobe[42]; // @[StreamController.scala 97:28:@45001.4]
  assign io_dram_wdata_bits_wstrb_22 = wdata_io_out_bits_strobe[41]; // @[StreamController.scala 97:28:@45002.4]
  assign io_dram_wdata_bits_wstrb_23 = wdata_io_out_bits_strobe[40]; // @[StreamController.scala 97:28:@45003.4]
  assign io_dram_wdata_bits_wstrb_24 = wdata_io_out_bits_strobe[39]; // @[StreamController.scala 97:28:@45004.4]
  assign io_dram_wdata_bits_wstrb_25 = wdata_io_out_bits_strobe[38]; // @[StreamController.scala 97:28:@45005.4]
  assign io_dram_wdata_bits_wstrb_26 = wdata_io_out_bits_strobe[37]; // @[StreamController.scala 97:28:@45006.4]
  assign io_dram_wdata_bits_wstrb_27 = wdata_io_out_bits_strobe[36]; // @[StreamController.scala 97:28:@45007.4]
  assign io_dram_wdata_bits_wstrb_28 = wdata_io_out_bits_strobe[35]; // @[StreamController.scala 97:28:@45008.4]
  assign io_dram_wdata_bits_wstrb_29 = wdata_io_out_bits_strobe[34]; // @[StreamController.scala 97:28:@45009.4]
  assign io_dram_wdata_bits_wstrb_30 = wdata_io_out_bits_strobe[33]; // @[StreamController.scala 97:28:@45010.4]
  assign io_dram_wdata_bits_wstrb_31 = wdata_io_out_bits_strobe[32]; // @[StreamController.scala 97:28:@45011.4]
  assign io_dram_wdata_bits_wstrb_32 = wdata_io_out_bits_strobe[31]; // @[StreamController.scala 97:28:@45012.4]
  assign io_dram_wdata_bits_wstrb_33 = wdata_io_out_bits_strobe[30]; // @[StreamController.scala 97:28:@45013.4]
  assign io_dram_wdata_bits_wstrb_34 = wdata_io_out_bits_strobe[29]; // @[StreamController.scala 97:28:@45014.4]
  assign io_dram_wdata_bits_wstrb_35 = wdata_io_out_bits_strobe[28]; // @[StreamController.scala 97:28:@45015.4]
  assign io_dram_wdata_bits_wstrb_36 = wdata_io_out_bits_strobe[27]; // @[StreamController.scala 97:28:@45016.4]
  assign io_dram_wdata_bits_wstrb_37 = wdata_io_out_bits_strobe[26]; // @[StreamController.scala 97:28:@45017.4]
  assign io_dram_wdata_bits_wstrb_38 = wdata_io_out_bits_strobe[25]; // @[StreamController.scala 97:28:@45018.4]
  assign io_dram_wdata_bits_wstrb_39 = wdata_io_out_bits_strobe[24]; // @[StreamController.scala 97:28:@45019.4]
  assign io_dram_wdata_bits_wstrb_40 = wdata_io_out_bits_strobe[23]; // @[StreamController.scala 97:28:@45020.4]
  assign io_dram_wdata_bits_wstrb_41 = wdata_io_out_bits_strobe[22]; // @[StreamController.scala 97:28:@45021.4]
  assign io_dram_wdata_bits_wstrb_42 = wdata_io_out_bits_strobe[21]; // @[StreamController.scala 97:28:@45022.4]
  assign io_dram_wdata_bits_wstrb_43 = wdata_io_out_bits_strobe[20]; // @[StreamController.scala 97:28:@45023.4]
  assign io_dram_wdata_bits_wstrb_44 = wdata_io_out_bits_strobe[19]; // @[StreamController.scala 97:28:@45024.4]
  assign io_dram_wdata_bits_wstrb_45 = wdata_io_out_bits_strobe[18]; // @[StreamController.scala 97:28:@45025.4]
  assign io_dram_wdata_bits_wstrb_46 = wdata_io_out_bits_strobe[17]; // @[StreamController.scala 97:28:@45026.4]
  assign io_dram_wdata_bits_wstrb_47 = wdata_io_out_bits_strobe[16]; // @[StreamController.scala 97:28:@45027.4]
  assign io_dram_wdata_bits_wstrb_48 = wdata_io_out_bits_strobe[15]; // @[StreamController.scala 97:28:@45028.4]
  assign io_dram_wdata_bits_wstrb_49 = wdata_io_out_bits_strobe[14]; // @[StreamController.scala 97:28:@45029.4]
  assign io_dram_wdata_bits_wstrb_50 = wdata_io_out_bits_strobe[13]; // @[StreamController.scala 97:28:@45030.4]
  assign io_dram_wdata_bits_wstrb_51 = wdata_io_out_bits_strobe[12]; // @[StreamController.scala 97:28:@45031.4]
  assign io_dram_wdata_bits_wstrb_52 = wdata_io_out_bits_strobe[11]; // @[StreamController.scala 97:28:@45032.4]
  assign io_dram_wdata_bits_wstrb_53 = wdata_io_out_bits_strobe[10]; // @[StreamController.scala 97:28:@45033.4]
  assign io_dram_wdata_bits_wstrb_54 = wdata_io_out_bits_strobe[9]; // @[StreamController.scala 97:28:@45034.4]
  assign io_dram_wdata_bits_wstrb_55 = wdata_io_out_bits_strobe[8]; // @[StreamController.scala 97:28:@45035.4]
  assign io_dram_wdata_bits_wstrb_56 = wdata_io_out_bits_strobe[7]; // @[StreamController.scala 97:28:@45036.4]
  assign io_dram_wdata_bits_wstrb_57 = wdata_io_out_bits_strobe[6]; // @[StreamController.scala 97:28:@45037.4]
  assign io_dram_wdata_bits_wstrb_58 = wdata_io_out_bits_strobe[5]; // @[StreamController.scala 97:28:@45038.4]
  assign io_dram_wdata_bits_wstrb_59 = wdata_io_out_bits_strobe[4]; // @[StreamController.scala 97:28:@45039.4]
  assign io_dram_wdata_bits_wstrb_60 = wdata_io_out_bits_strobe[3]; // @[StreamController.scala 97:28:@45040.4]
  assign io_dram_wdata_bits_wstrb_61 = wdata_io_out_bits_strobe[2]; // @[StreamController.scala 97:28:@45041.4]
  assign io_dram_wdata_bits_wstrb_62 = wdata_io_out_bits_strobe[1]; // @[StreamController.scala 97:28:@45042.4]
  assign io_dram_wdata_bits_wstrb_63 = wdata_io_out_bits_strobe[0]; // @[StreamController.scala 97:28:@45043.4]
  assign io_dram_wresp_ready = wresp_io_in_ready; // @[StreamController.scala 104:23:@45312.4]
  assign io_store_cmd_ready = cmd_io_in_ready; // @[StreamController.scala 79:22:@44796.4]
  assign io_store_data_ready = wdata_io_in_ready; // @[StreamController.scala 93:23:@44833.4]
  assign io_store_wresp_valid = wresp_io_out_valid; // @[StreamController.scala 106:24:@45313.4]
  assign io_store_wresp_bits = wresp_io_out_bits; // @[StreamController.scala 107:23:@45314.4]
  assign cmd_clock = clock; // @[:@44399.4]
  assign cmd_reset = reset; // @[:@44400.4]
  assign cmd_io_in_valid = io_store_cmd_valid; // @[StreamController.scala 77:19:@44793.4]
  assign cmd_io_in_bits_addr = io_store_cmd_bits_addr; // @[StreamController.scala 78:18:@44795.4]
  assign cmd_io_in_bits_size = io_store_cmd_bits_size; // @[StreamController.scala 78:18:@44794.4]
  assign cmd_io_out_ready = io_dram_cmd_ready; // @[StreamController.scala 80:20:@44797.4]
  assign wdata_clock = clock; // @[:@44805.4]
  assign wdata_reset = reset; // @[:@44806.4]
  assign wdata_io_in_valid = io_store_data_valid; // @[StreamController.scala 90:21:@44830.4]
  assign wdata_io_in_bits_data_0 = io_store_data_bits_wdata_0; // @[StreamController.scala 91:25:@44831.4]
  assign wdata_io_in_bits_strobe = io_store_data_bits_wstrb; // @[StreamController.scala 92:27:@44832.4]
  assign wdata_io_out_ready = io_dram_wdata_ready; // @[StreamController.scala 98:22:@45044.4]
  assign wresp_clock = clock; // @[:@45046.4]
  assign wresp_reset = reset; // @[:@45047.4]
  assign wresp_io_in_valid = io_dram_wresp_valid; // @[StreamController.scala 102:21:@45310.4]
  assign wresp_io_in_bits = 1'h1; // @[StreamController.scala 103:20:@45311.4]
  assign wresp_io_out_ready = io_store_wresp_ready; // @[StreamController.scala 108:22:@45315.4]
  assign wresp_io_banks_0_wdata_valid = 1'h0;
  assign wresp_io_banks_0_wdata_bits = 1'h0;
  assign wresp_io_banks_1_wdata_valid = 1'h0;
  assign wresp_io_banks_1_wdata_bits = 1'h0;
  assign wresp_io_banks_2_wdata_valid = 1'h0;
  assign wresp_io_banks_2_wdata_bits = 1'h0;
  assign wresp_io_banks_3_wdata_valid = 1'h0;
  assign wresp_io_banks_3_wdata_bits = 1'h0;
  assign wresp_io_banks_4_wdata_valid = 1'h0;
  assign wresp_io_banks_4_wdata_bits = 1'h0;
  assign wresp_io_banks_5_wdata_valid = 1'h0;
  assign wresp_io_banks_5_wdata_bits = 1'h0;
  assign wresp_io_banks_6_wdata_valid = 1'h0;
  assign wresp_io_banks_6_wdata_bits = 1'h0;
  assign wresp_io_banks_7_wdata_valid = 1'h0;
  assign wresp_io_banks_7_wdata_bits = 1'h0;
  assign wresp_io_banks_8_wdata_valid = 1'h0;
  assign wresp_io_banks_8_wdata_bits = 1'h0;
  assign wresp_io_banks_9_wdata_valid = 1'h0;
  assign wresp_io_banks_9_wdata_bits = 1'h0;
  assign wresp_io_banks_10_wdata_valid = 1'h0;
  assign wresp_io_banks_10_wdata_bits = 1'h0;
  assign wresp_io_banks_11_wdata_valid = 1'h0;
  assign wresp_io_banks_11_wdata_bits = 1'h0;
  assign wresp_io_banks_12_wdata_valid = 1'h0;
  assign wresp_io_banks_12_wdata_bits = 1'h0;
  assign wresp_io_banks_13_wdata_valid = 1'h0;
  assign wresp_io_banks_13_wdata_bits = 1'h0;
  assign wresp_io_banks_14_wdata_valid = 1'h0;
  assign wresp_io_banks_14_wdata_bits = 1'h0;
  assign wresp_io_banks_15_wdata_valid = 1'h0;
  assign wresp_io_banks_15_wdata_bits = 1'h0;
  assign wresp_io_banks_16_wdata_valid = 1'h0;
  assign wresp_io_banks_16_wdata_bits = 1'h0;
  assign wresp_io_banks_17_wdata_valid = 1'h0;
  assign wresp_io_banks_17_wdata_bits = 1'h0;
  assign wresp_io_banks_18_wdata_valid = 1'h0;
  assign wresp_io_banks_18_wdata_bits = 1'h0;
  assign wresp_io_banks_19_wdata_valid = 1'h0;
  assign wresp_io_banks_19_wdata_bits = 1'h0;
  assign wresp_io_banks_20_wdata_valid = 1'h0;
  assign wresp_io_banks_20_wdata_bits = 1'h0;
  assign wresp_io_banks_21_wdata_valid = 1'h0;
  assign wresp_io_banks_21_wdata_bits = 1'h0;
  assign wresp_io_banks_22_wdata_valid = 1'h0;
  assign wresp_io_banks_22_wdata_bits = 1'h0;
  assign wresp_io_banks_23_wdata_valid = 1'h0;
  assign wresp_io_banks_23_wdata_bits = 1'h0;
  assign wresp_io_banks_24_wdata_valid = 1'h0;
  assign wresp_io_banks_24_wdata_bits = 1'h0;
  assign wresp_io_banks_25_wdata_valid = 1'h0;
  assign wresp_io_banks_25_wdata_bits = 1'h0;
  assign wresp_io_banks_26_wdata_valid = 1'h0;
  assign wresp_io_banks_26_wdata_bits = 1'h0;
  assign wresp_io_banks_27_wdata_valid = 1'h0;
  assign wresp_io_banks_27_wdata_bits = 1'h0;
  assign wresp_io_banks_28_wdata_valid = 1'h0;
  assign wresp_io_banks_28_wdata_bits = 1'h0;
  assign wresp_io_banks_29_wdata_valid = 1'h0;
  assign wresp_io_banks_29_wdata_bits = 1'h0;
  assign wresp_io_banks_30_wdata_valid = 1'h0;
  assign wresp_io_banks_30_wdata_bits = 1'h0;
  assign wresp_io_banks_31_wdata_valid = 1'h0;
  assign wresp_io_banks_31_wdata_bits = 1'h0;
  assign wresp_io_banks_32_wdata_valid = 1'h0;
  assign wresp_io_banks_32_wdata_bits = 1'h0;
  assign wresp_io_banks_33_wdata_valid = 1'h0;
  assign wresp_io_banks_33_wdata_bits = 1'h0;
  assign wresp_io_banks_34_wdata_valid = 1'h0;
  assign wresp_io_banks_34_wdata_bits = 1'h0;
  assign wresp_io_banks_35_wdata_valid = 1'h0;
  assign wresp_io_banks_35_wdata_bits = 1'h0;
  assign wresp_io_banks_36_wdata_valid = 1'h0;
  assign wresp_io_banks_36_wdata_bits = 1'h0;
  assign wresp_io_banks_37_wdata_valid = 1'h0;
  assign wresp_io_banks_37_wdata_bits = 1'h0;
  assign wresp_io_banks_38_wdata_valid = 1'h0;
  assign wresp_io_banks_38_wdata_bits = 1'h0;
  assign wresp_io_banks_39_wdata_valid = 1'h0;
  assign wresp_io_banks_39_wdata_bits = 1'h0;
  assign wresp_io_banks_40_wdata_valid = 1'h0;
  assign wresp_io_banks_40_wdata_bits = 1'h0;
  assign wresp_io_banks_41_wdata_valid = 1'h0;
  assign wresp_io_banks_41_wdata_bits = 1'h0;
  assign wresp_io_banks_42_wdata_valid = 1'h0;
  assign wresp_io_banks_42_wdata_bits = 1'h0;
  assign wresp_io_banks_43_wdata_valid = 1'h0;
  assign wresp_io_banks_43_wdata_bits = 1'h0;
  assign wresp_io_banks_44_wdata_valid = 1'h0;
  assign wresp_io_banks_44_wdata_bits = 1'h0;
  assign wresp_io_banks_45_wdata_valid = 1'h0;
  assign wresp_io_banks_45_wdata_bits = 1'h0;
  assign wresp_io_banks_46_wdata_valid = 1'h0;
  assign wresp_io_banks_46_wdata_bits = 1'h0;
  assign wresp_io_banks_47_wdata_valid = 1'h0;
  assign wresp_io_banks_47_wdata_bits = 1'h0;
  assign wresp_io_banks_48_wdata_valid = 1'h0;
  assign wresp_io_banks_48_wdata_bits = 1'h0;
  assign wresp_io_banks_49_wdata_valid = 1'h0;
  assign wresp_io_banks_49_wdata_bits = 1'h0;
  assign wresp_io_banks_50_wdata_valid = 1'h0;
  assign wresp_io_banks_50_wdata_bits = 1'h0;
  assign wresp_io_banks_51_wdata_valid = 1'h0;
  assign wresp_io_banks_51_wdata_bits = 1'h0;
  assign wresp_io_banks_52_wdata_valid = 1'h0;
  assign wresp_io_banks_52_wdata_bits = 1'h0;
  assign wresp_io_banks_53_wdata_valid = 1'h0;
  assign wresp_io_banks_53_wdata_bits = 1'h0;
  assign wresp_io_banks_54_wdata_valid = 1'h0;
  assign wresp_io_banks_54_wdata_bits = 1'h0;
  assign wresp_io_banks_55_wdata_valid = 1'h0;
  assign wresp_io_banks_55_wdata_bits = 1'h0;
  assign wresp_io_banks_56_wdata_valid = 1'h0;
  assign wresp_io_banks_56_wdata_bits = 1'h0;
  assign wresp_io_banks_57_wdata_valid = 1'h0;
  assign wresp_io_banks_57_wdata_bits = 1'h0;
  assign wresp_io_banks_58_wdata_valid = 1'h0;
  assign wresp_io_banks_58_wdata_bits = 1'h0;
  assign wresp_io_banks_59_wdata_valid = 1'h0;
  assign wresp_io_banks_59_wdata_bits = 1'h0;
  assign wresp_io_banks_60_wdata_valid = 1'h0;
  assign wresp_io_banks_60_wdata_bits = 1'h0;
  assign wresp_io_banks_61_wdata_valid = 1'h0;
  assign wresp_io_banks_61_wdata_bits = 1'h0;
  assign wresp_io_banks_62_wdata_valid = 1'h0;
  assign wresp_io_banks_62_wdata_bits = 1'h0;
  assign wresp_io_banks_63_wdata_valid = 1'h0;
  assign wresp_io_banks_63_wdata_bits = 1'h0;
endmodule
module MuxPipe( // @[:@45381.2]
  output        io_in_ready, // @[:@45384.4]
  input         io_in_valid, // @[:@45384.4]
  input  [63:0] io_in_bits_0_addr, // @[:@45384.4]
  input  [31:0] io_in_bits_0_size, // @[:@45384.4]
  input         io_in_bits_0_isWr, // @[:@45384.4]
  input  [31:0] io_in_bits_0_tag, // @[:@45384.4]
  input         io_out_ready, // @[:@45384.4]
  output        io_out_valid, // @[:@45384.4]
  output [63:0] io_out_bits_addr, // @[:@45384.4]
  output [31:0] io_out_bits_size, // @[:@45384.4]
  output        io_out_bits_isWr, // @[:@45384.4]
  output [31:0] io_out_bits_tag // @[:@45384.4]
);
  wire  _T_42; // @[MuxN.scala 28:31:@45386.4]
  assign _T_42 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@45386.4]
  assign io_in_ready = io_out_ready | _T_42; // @[MuxN.scala 71:15:@45395.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@45394.4]
  assign io_out_bits_addr = io_in_bits_0_addr; // @[MuxN.scala 72:15:@45400.4]
  assign io_out_bits_size = io_in_bits_0_size; // @[MuxN.scala 72:15:@45399.4]
  assign io_out_bits_isWr = io_in_bits_0_isWr; // @[MuxN.scala 72:15:@45397.4]
  assign io_out_bits_tag = io_in_bits_0_tag; // @[MuxN.scala 72:15:@45396.4]
endmodule
module MuxPipe_1( // @[:@45402.2]
  output        io_in_ready, // @[:@45405.4]
  input         io_in_valid, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_0, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_1, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_2, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_3, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_4, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_5, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_6, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_7, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_8, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_9, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_10, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_11, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_12, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_13, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_14, // @[:@45405.4]
  input  [31:0] io_in_bits_0_wdata_15, // @[:@45405.4]
  input         io_in_bits_0_wstrb_0, // @[:@45405.4]
  input         io_in_bits_0_wstrb_1, // @[:@45405.4]
  input         io_in_bits_0_wstrb_2, // @[:@45405.4]
  input         io_in_bits_0_wstrb_3, // @[:@45405.4]
  input         io_in_bits_0_wstrb_4, // @[:@45405.4]
  input         io_in_bits_0_wstrb_5, // @[:@45405.4]
  input         io_in_bits_0_wstrb_6, // @[:@45405.4]
  input         io_in_bits_0_wstrb_7, // @[:@45405.4]
  input         io_in_bits_0_wstrb_8, // @[:@45405.4]
  input         io_in_bits_0_wstrb_9, // @[:@45405.4]
  input         io_in_bits_0_wstrb_10, // @[:@45405.4]
  input         io_in_bits_0_wstrb_11, // @[:@45405.4]
  input         io_in_bits_0_wstrb_12, // @[:@45405.4]
  input         io_in_bits_0_wstrb_13, // @[:@45405.4]
  input         io_in_bits_0_wstrb_14, // @[:@45405.4]
  input         io_in_bits_0_wstrb_15, // @[:@45405.4]
  input         io_in_bits_0_wstrb_16, // @[:@45405.4]
  input         io_in_bits_0_wstrb_17, // @[:@45405.4]
  input         io_in_bits_0_wstrb_18, // @[:@45405.4]
  input         io_in_bits_0_wstrb_19, // @[:@45405.4]
  input         io_in_bits_0_wstrb_20, // @[:@45405.4]
  input         io_in_bits_0_wstrb_21, // @[:@45405.4]
  input         io_in_bits_0_wstrb_22, // @[:@45405.4]
  input         io_in_bits_0_wstrb_23, // @[:@45405.4]
  input         io_in_bits_0_wstrb_24, // @[:@45405.4]
  input         io_in_bits_0_wstrb_25, // @[:@45405.4]
  input         io_in_bits_0_wstrb_26, // @[:@45405.4]
  input         io_in_bits_0_wstrb_27, // @[:@45405.4]
  input         io_in_bits_0_wstrb_28, // @[:@45405.4]
  input         io_in_bits_0_wstrb_29, // @[:@45405.4]
  input         io_in_bits_0_wstrb_30, // @[:@45405.4]
  input         io_in_bits_0_wstrb_31, // @[:@45405.4]
  input         io_in_bits_0_wstrb_32, // @[:@45405.4]
  input         io_in_bits_0_wstrb_33, // @[:@45405.4]
  input         io_in_bits_0_wstrb_34, // @[:@45405.4]
  input         io_in_bits_0_wstrb_35, // @[:@45405.4]
  input         io_in_bits_0_wstrb_36, // @[:@45405.4]
  input         io_in_bits_0_wstrb_37, // @[:@45405.4]
  input         io_in_bits_0_wstrb_38, // @[:@45405.4]
  input         io_in_bits_0_wstrb_39, // @[:@45405.4]
  input         io_in_bits_0_wstrb_40, // @[:@45405.4]
  input         io_in_bits_0_wstrb_41, // @[:@45405.4]
  input         io_in_bits_0_wstrb_42, // @[:@45405.4]
  input         io_in_bits_0_wstrb_43, // @[:@45405.4]
  input         io_in_bits_0_wstrb_44, // @[:@45405.4]
  input         io_in_bits_0_wstrb_45, // @[:@45405.4]
  input         io_in_bits_0_wstrb_46, // @[:@45405.4]
  input         io_in_bits_0_wstrb_47, // @[:@45405.4]
  input         io_in_bits_0_wstrb_48, // @[:@45405.4]
  input         io_in_bits_0_wstrb_49, // @[:@45405.4]
  input         io_in_bits_0_wstrb_50, // @[:@45405.4]
  input         io_in_bits_0_wstrb_51, // @[:@45405.4]
  input         io_in_bits_0_wstrb_52, // @[:@45405.4]
  input         io_in_bits_0_wstrb_53, // @[:@45405.4]
  input         io_in_bits_0_wstrb_54, // @[:@45405.4]
  input         io_in_bits_0_wstrb_55, // @[:@45405.4]
  input         io_in_bits_0_wstrb_56, // @[:@45405.4]
  input         io_in_bits_0_wstrb_57, // @[:@45405.4]
  input         io_in_bits_0_wstrb_58, // @[:@45405.4]
  input         io_in_bits_0_wstrb_59, // @[:@45405.4]
  input         io_in_bits_0_wstrb_60, // @[:@45405.4]
  input         io_in_bits_0_wstrb_61, // @[:@45405.4]
  input         io_in_bits_0_wstrb_62, // @[:@45405.4]
  input         io_in_bits_0_wstrb_63, // @[:@45405.4]
  input         io_out_ready, // @[:@45405.4]
  output        io_out_valid, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_0, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_1, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_2, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_3, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_4, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_5, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_6, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_7, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_8, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_9, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_10, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_11, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_12, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_13, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_14, // @[:@45405.4]
  output [31:0] io_out_bits_wdata_15, // @[:@45405.4]
  output        io_out_bits_wstrb_0, // @[:@45405.4]
  output        io_out_bits_wstrb_1, // @[:@45405.4]
  output        io_out_bits_wstrb_2, // @[:@45405.4]
  output        io_out_bits_wstrb_3, // @[:@45405.4]
  output        io_out_bits_wstrb_4, // @[:@45405.4]
  output        io_out_bits_wstrb_5, // @[:@45405.4]
  output        io_out_bits_wstrb_6, // @[:@45405.4]
  output        io_out_bits_wstrb_7, // @[:@45405.4]
  output        io_out_bits_wstrb_8, // @[:@45405.4]
  output        io_out_bits_wstrb_9, // @[:@45405.4]
  output        io_out_bits_wstrb_10, // @[:@45405.4]
  output        io_out_bits_wstrb_11, // @[:@45405.4]
  output        io_out_bits_wstrb_12, // @[:@45405.4]
  output        io_out_bits_wstrb_13, // @[:@45405.4]
  output        io_out_bits_wstrb_14, // @[:@45405.4]
  output        io_out_bits_wstrb_15, // @[:@45405.4]
  output        io_out_bits_wstrb_16, // @[:@45405.4]
  output        io_out_bits_wstrb_17, // @[:@45405.4]
  output        io_out_bits_wstrb_18, // @[:@45405.4]
  output        io_out_bits_wstrb_19, // @[:@45405.4]
  output        io_out_bits_wstrb_20, // @[:@45405.4]
  output        io_out_bits_wstrb_21, // @[:@45405.4]
  output        io_out_bits_wstrb_22, // @[:@45405.4]
  output        io_out_bits_wstrb_23, // @[:@45405.4]
  output        io_out_bits_wstrb_24, // @[:@45405.4]
  output        io_out_bits_wstrb_25, // @[:@45405.4]
  output        io_out_bits_wstrb_26, // @[:@45405.4]
  output        io_out_bits_wstrb_27, // @[:@45405.4]
  output        io_out_bits_wstrb_28, // @[:@45405.4]
  output        io_out_bits_wstrb_29, // @[:@45405.4]
  output        io_out_bits_wstrb_30, // @[:@45405.4]
  output        io_out_bits_wstrb_31, // @[:@45405.4]
  output        io_out_bits_wstrb_32, // @[:@45405.4]
  output        io_out_bits_wstrb_33, // @[:@45405.4]
  output        io_out_bits_wstrb_34, // @[:@45405.4]
  output        io_out_bits_wstrb_35, // @[:@45405.4]
  output        io_out_bits_wstrb_36, // @[:@45405.4]
  output        io_out_bits_wstrb_37, // @[:@45405.4]
  output        io_out_bits_wstrb_38, // @[:@45405.4]
  output        io_out_bits_wstrb_39, // @[:@45405.4]
  output        io_out_bits_wstrb_40, // @[:@45405.4]
  output        io_out_bits_wstrb_41, // @[:@45405.4]
  output        io_out_bits_wstrb_42, // @[:@45405.4]
  output        io_out_bits_wstrb_43, // @[:@45405.4]
  output        io_out_bits_wstrb_44, // @[:@45405.4]
  output        io_out_bits_wstrb_45, // @[:@45405.4]
  output        io_out_bits_wstrb_46, // @[:@45405.4]
  output        io_out_bits_wstrb_47, // @[:@45405.4]
  output        io_out_bits_wstrb_48, // @[:@45405.4]
  output        io_out_bits_wstrb_49, // @[:@45405.4]
  output        io_out_bits_wstrb_50, // @[:@45405.4]
  output        io_out_bits_wstrb_51, // @[:@45405.4]
  output        io_out_bits_wstrb_52, // @[:@45405.4]
  output        io_out_bits_wstrb_53, // @[:@45405.4]
  output        io_out_bits_wstrb_54, // @[:@45405.4]
  output        io_out_bits_wstrb_55, // @[:@45405.4]
  output        io_out_bits_wstrb_56, // @[:@45405.4]
  output        io_out_bits_wstrb_57, // @[:@45405.4]
  output        io_out_bits_wstrb_58, // @[:@45405.4]
  output        io_out_bits_wstrb_59, // @[:@45405.4]
  output        io_out_bits_wstrb_60, // @[:@45405.4]
  output        io_out_bits_wstrb_61, // @[:@45405.4]
  output        io_out_bits_wstrb_62, // @[:@45405.4]
  output        io_out_bits_wstrb_63 // @[:@45405.4]
);
  wire  _T_146; // @[MuxN.scala 28:31:@45407.4]
  assign _T_146 = io_out_valid == 1'h0; // @[MuxN.scala 28:31:@45407.4]
  assign io_in_ready = io_out_ready | _T_146; // @[MuxN.scala 71:15:@45492.4]
  assign io_out_valid = io_in_valid; // @[MuxN.scala 70:16:@45491.4]
  assign io_out_bits_wdata_0 = io_in_bits_0_wdata_0; // @[MuxN.scala 72:15:@45558.4]
  assign io_out_bits_wdata_1 = io_in_bits_0_wdata_1; // @[MuxN.scala 72:15:@45559.4]
  assign io_out_bits_wdata_2 = io_in_bits_0_wdata_2; // @[MuxN.scala 72:15:@45560.4]
  assign io_out_bits_wdata_3 = io_in_bits_0_wdata_3; // @[MuxN.scala 72:15:@45561.4]
  assign io_out_bits_wdata_4 = io_in_bits_0_wdata_4; // @[MuxN.scala 72:15:@45562.4]
  assign io_out_bits_wdata_5 = io_in_bits_0_wdata_5; // @[MuxN.scala 72:15:@45563.4]
  assign io_out_bits_wdata_6 = io_in_bits_0_wdata_6; // @[MuxN.scala 72:15:@45564.4]
  assign io_out_bits_wdata_7 = io_in_bits_0_wdata_7; // @[MuxN.scala 72:15:@45565.4]
  assign io_out_bits_wdata_8 = io_in_bits_0_wdata_8; // @[MuxN.scala 72:15:@45566.4]
  assign io_out_bits_wdata_9 = io_in_bits_0_wdata_9; // @[MuxN.scala 72:15:@45567.4]
  assign io_out_bits_wdata_10 = io_in_bits_0_wdata_10; // @[MuxN.scala 72:15:@45568.4]
  assign io_out_bits_wdata_11 = io_in_bits_0_wdata_11; // @[MuxN.scala 72:15:@45569.4]
  assign io_out_bits_wdata_12 = io_in_bits_0_wdata_12; // @[MuxN.scala 72:15:@45570.4]
  assign io_out_bits_wdata_13 = io_in_bits_0_wdata_13; // @[MuxN.scala 72:15:@45571.4]
  assign io_out_bits_wdata_14 = io_in_bits_0_wdata_14; // @[MuxN.scala 72:15:@45572.4]
  assign io_out_bits_wdata_15 = io_in_bits_0_wdata_15; // @[MuxN.scala 72:15:@45573.4]
  assign io_out_bits_wstrb_0 = io_in_bits_0_wstrb_0; // @[MuxN.scala 72:15:@45494.4]
  assign io_out_bits_wstrb_1 = io_in_bits_0_wstrb_1; // @[MuxN.scala 72:15:@45495.4]
  assign io_out_bits_wstrb_2 = io_in_bits_0_wstrb_2; // @[MuxN.scala 72:15:@45496.4]
  assign io_out_bits_wstrb_3 = io_in_bits_0_wstrb_3; // @[MuxN.scala 72:15:@45497.4]
  assign io_out_bits_wstrb_4 = io_in_bits_0_wstrb_4; // @[MuxN.scala 72:15:@45498.4]
  assign io_out_bits_wstrb_5 = io_in_bits_0_wstrb_5; // @[MuxN.scala 72:15:@45499.4]
  assign io_out_bits_wstrb_6 = io_in_bits_0_wstrb_6; // @[MuxN.scala 72:15:@45500.4]
  assign io_out_bits_wstrb_7 = io_in_bits_0_wstrb_7; // @[MuxN.scala 72:15:@45501.4]
  assign io_out_bits_wstrb_8 = io_in_bits_0_wstrb_8; // @[MuxN.scala 72:15:@45502.4]
  assign io_out_bits_wstrb_9 = io_in_bits_0_wstrb_9; // @[MuxN.scala 72:15:@45503.4]
  assign io_out_bits_wstrb_10 = io_in_bits_0_wstrb_10; // @[MuxN.scala 72:15:@45504.4]
  assign io_out_bits_wstrb_11 = io_in_bits_0_wstrb_11; // @[MuxN.scala 72:15:@45505.4]
  assign io_out_bits_wstrb_12 = io_in_bits_0_wstrb_12; // @[MuxN.scala 72:15:@45506.4]
  assign io_out_bits_wstrb_13 = io_in_bits_0_wstrb_13; // @[MuxN.scala 72:15:@45507.4]
  assign io_out_bits_wstrb_14 = io_in_bits_0_wstrb_14; // @[MuxN.scala 72:15:@45508.4]
  assign io_out_bits_wstrb_15 = io_in_bits_0_wstrb_15; // @[MuxN.scala 72:15:@45509.4]
  assign io_out_bits_wstrb_16 = io_in_bits_0_wstrb_16; // @[MuxN.scala 72:15:@45510.4]
  assign io_out_bits_wstrb_17 = io_in_bits_0_wstrb_17; // @[MuxN.scala 72:15:@45511.4]
  assign io_out_bits_wstrb_18 = io_in_bits_0_wstrb_18; // @[MuxN.scala 72:15:@45512.4]
  assign io_out_bits_wstrb_19 = io_in_bits_0_wstrb_19; // @[MuxN.scala 72:15:@45513.4]
  assign io_out_bits_wstrb_20 = io_in_bits_0_wstrb_20; // @[MuxN.scala 72:15:@45514.4]
  assign io_out_bits_wstrb_21 = io_in_bits_0_wstrb_21; // @[MuxN.scala 72:15:@45515.4]
  assign io_out_bits_wstrb_22 = io_in_bits_0_wstrb_22; // @[MuxN.scala 72:15:@45516.4]
  assign io_out_bits_wstrb_23 = io_in_bits_0_wstrb_23; // @[MuxN.scala 72:15:@45517.4]
  assign io_out_bits_wstrb_24 = io_in_bits_0_wstrb_24; // @[MuxN.scala 72:15:@45518.4]
  assign io_out_bits_wstrb_25 = io_in_bits_0_wstrb_25; // @[MuxN.scala 72:15:@45519.4]
  assign io_out_bits_wstrb_26 = io_in_bits_0_wstrb_26; // @[MuxN.scala 72:15:@45520.4]
  assign io_out_bits_wstrb_27 = io_in_bits_0_wstrb_27; // @[MuxN.scala 72:15:@45521.4]
  assign io_out_bits_wstrb_28 = io_in_bits_0_wstrb_28; // @[MuxN.scala 72:15:@45522.4]
  assign io_out_bits_wstrb_29 = io_in_bits_0_wstrb_29; // @[MuxN.scala 72:15:@45523.4]
  assign io_out_bits_wstrb_30 = io_in_bits_0_wstrb_30; // @[MuxN.scala 72:15:@45524.4]
  assign io_out_bits_wstrb_31 = io_in_bits_0_wstrb_31; // @[MuxN.scala 72:15:@45525.4]
  assign io_out_bits_wstrb_32 = io_in_bits_0_wstrb_32; // @[MuxN.scala 72:15:@45526.4]
  assign io_out_bits_wstrb_33 = io_in_bits_0_wstrb_33; // @[MuxN.scala 72:15:@45527.4]
  assign io_out_bits_wstrb_34 = io_in_bits_0_wstrb_34; // @[MuxN.scala 72:15:@45528.4]
  assign io_out_bits_wstrb_35 = io_in_bits_0_wstrb_35; // @[MuxN.scala 72:15:@45529.4]
  assign io_out_bits_wstrb_36 = io_in_bits_0_wstrb_36; // @[MuxN.scala 72:15:@45530.4]
  assign io_out_bits_wstrb_37 = io_in_bits_0_wstrb_37; // @[MuxN.scala 72:15:@45531.4]
  assign io_out_bits_wstrb_38 = io_in_bits_0_wstrb_38; // @[MuxN.scala 72:15:@45532.4]
  assign io_out_bits_wstrb_39 = io_in_bits_0_wstrb_39; // @[MuxN.scala 72:15:@45533.4]
  assign io_out_bits_wstrb_40 = io_in_bits_0_wstrb_40; // @[MuxN.scala 72:15:@45534.4]
  assign io_out_bits_wstrb_41 = io_in_bits_0_wstrb_41; // @[MuxN.scala 72:15:@45535.4]
  assign io_out_bits_wstrb_42 = io_in_bits_0_wstrb_42; // @[MuxN.scala 72:15:@45536.4]
  assign io_out_bits_wstrb_43 = io_in_bits_0_wstrb_43; // @[MuxN.scala 72:15:@45537.4]
  assign io_out_bits_wstrb_44 = io_in_bits_0_wstrb_44; // @[MuxN.scala 72:15:@45538.4]
  assign io_out_bits_wstrb_45 = io_in_bits_0_wstrb_45; // @[MuxN.scala 72:15:@45539.4]
  assign io_out_bits_wstrb_46 = io_in_bits_0_wstrb_46; // @[MuxN.scala 72:15:@45540.4]
  assign io_out_bits_wstrb_47 = io_in_bits_0_wstrb_47; // @[MuxN.scala 72:15:@45541.4]
  assign io_out_bits_wstrb_48 = io_in_bits_0_wstrb_48; // @[MuxN.scala 72:15:@45542.4]
  assign io_out_bits_wstrb_49 = io_in_bits_0_wstrb_49; // @[MuxN.scala 72:15:@45543.4]
  assign io_out_bits_wstrb_50 = io_in_bits_0_wstrb_50; // @[MuxN.scala 72:15:@45544.4]
  assign io_out_bits_wstrb_51 = io_in_bits_0_wstrb_51; // @[MuxN.scala 72:15:@45545.4]
  assign io_out_bits_wstrb_52 = io_in_bits_0_wstrb_52; // @[MuxN.scala 72:15:@45546.4]
  assign io_out_bits_wstrb_53 = io_in_bits_0_wstrb_53; // @[MuxN.scala 72:15:@45547.4]
  assign io_out_bits_wstrb_54 = io_in_bits_0_wstrb_54; // @[MuxN.scala 72:15:@45548.4]
  assign io_out_bits_wstrb_55 = io_in_bits_0_wstrb_55; // @[MuxN.scala 72:15:@45549.4]
  assign io_out_bits_wstrb_56 = io_in_bits_0_wstrb_56; // @[MuxN.scala 72:15:@45550.4]
  assign io_out_bits_wstrb_57 = io_in_bits_0_wstrb_57; // @[MuxN.scala 72:15:@45551.4]
  assign io_out_bits_wstrb_58 = io_in_bits_0_wstrb_58; // @[MuxN.scala 72:15:@45552.4]
  assign io_out_bits_wstrb_59 = io_in_bits_0_wstrb_59; // @[MuxN.scala 72:15:@45553.4]
  assign io_out_bits_wstrb_60 = io_in_bits_0_wstrb_60; // @[MuxN.scala 72:15:@45554.4]
  assign io_out_bits_wstrb_61 = io_in_bits_0_wstrb_61; // @[MuxN.scala 72:15:@45555.4]
  assign io_out_bits_wstrb_62 = io_in_bits_0_wstrb_62; // @[MuxN.scala 72:15:@45556.4]
  assign io_out_bits_wstrb_63 = io_in_bits_0_wstrb_63; // @[MuxN.scala 72:15:@45557.4]
endmodule
module ElementCounter( // @[:@45575.2]
  input         clock, // @[:@45576.4]
  input         reset, // @[:@45577.4]
  input         io_reset, // @[:@45578.4]
  input         io_enable, // @[:@45578.4]
  output [31:0] io_out // @[:@45578.4]
);
  reg [31:0] count; // @[Counter.scala 37:22:@45580.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_14; // @[Counter.scala 39:24:@45581.4]
  wire [31:0] newCount; // @[Counter.scala 39:24:@45582.4]
  wire [31:0] _GEN_0; // @[Counter.scala 43:26:@45587.6]
  wire [31:0] _GEN_1; // @[Counter.scala 41:18:@45583.4]
  assign _T_14 = count + 32'h1; // @[Counter.scala 39:24:@45581.4]
  assign newCount = count + 32'h1; // @[Counter.scala 39:24:@45582.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 43:26:@45587.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 41:18:@45583.4]
  assign io_out = count; // @[Counter.scala 47:10:@45590.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module StreamArbiter( // @[:@45592.2]
  input         clock, // @[:@45593.4]
  input         reset, // @[:@45594.4]
  output        io_app_0_cmd_ready, // @[:@45595.4]
  input         io_app_0_cmd_valid, // @[:@45595.4]
  input  [63:0] io_app_0_cmd_bits_addr, // @[:@45595.4]
  input  [31:0] io_app_0_cmd_bits_size, // @[:@45595.4]
  input         io_app_0_cmd_bits_isWr, // @[:@45595.4]
  input  [31:0] io_app_0_cmd_bits_tag, // @[:@45595.4]
  output        io_app_0_wdata_ready, // @[:@45595.4]
  input         io_app_0_wdata_valid, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_0, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_1, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_2, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_3, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_4, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_5, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_6, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_7, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_8, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_9, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_10, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_11, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_12, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_13, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_14, // @[:@45595.4]
  input  [31:0] io_app_0_wdata_bits_wdata_15, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_0, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_1, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_2, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_3, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_4, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_5, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_6, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_7, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_8, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_9, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_10, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_11, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_12, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_13, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_14, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_15, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_16, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_17, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_18, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_19, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_20, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_21, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_22, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_23, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_24, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_25, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_26, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_27, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_28, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_29, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_30, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_31, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_32, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_33, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_34, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_35, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_36, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_37, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_38, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_39, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_40, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_41, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_42, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_43, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_44, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_45, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_46, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_47, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_48, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_49, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_50, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_51, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_52, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_53, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_54, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_55, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_56, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_57, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_58, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_59, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_60, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_61, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_62, // @[:@45595.4]
  input         io_app_0_wdata_bits_wstrb_63, // @[:@45595.4]
  input         io_app_0_rresp_ready, // @[:@45595.4]
  input         io_app_0_wresp_ready, // @[:@45595.4]
  output        io_app_0_wresp_valid, // @[:@45595.4]
  input         io_dram_cmd_ready, // @[:@45595.4]
  output        io_dram_cmd_valid, // @[:@45595.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@45595.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@45595.4]
  output        io_dram_cmd_bits_isWr, // @[:@45595.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@45595.4]
  input         io_dram_wdata_ready, // @[:@45595.4]
  output        io_dram_wdata_valid, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@45595.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@45595.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@45595.4]
  output        io_dram_rresp_ready, // @[:@45595.4]
  output        io_dram_wresp_ready, // @[:@45595.4]
  input         io_dram_wresp_valid, // @[:@45595.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@45595.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@45824.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@45824.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@45824.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@45824.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@45824.4]
  wire  RetimeWrapper_1_clock; // @[package.scala 93:22:@45831.4]
  wire  RetimeWrapper_1_reset; // @[package.scala 93:22:@45831.4]
  wire  RetimeWrapper_1_io_flow; // @[package.scala 93:22:@45831.4]
  wire  RetimeWrapper_1_io_in; // @[package.scala 93:22:@45831.4]
  wire  RetimeWrapper_1_io_out; // @[package.scala 93:22:@45831.4]
  wire  cmdMux_io_in_ready; // @[StreamArbiter.scala 25:22:@45841.4]
  wire  cmdMux_io_in_valid; // @[StreamArbiter.scala 25:22:@45841.4]
  wire [63:0] cmdMux_io_in_bits_0_addr; // @[StreamArbiter.scala 25:22:@45841.4]
  wire [31:0] cmdMux_io_in_bits_0_size; // @[StreamArbiter.scala 25:22:@45841.4]
  wire  cmdMux_io_in_bits_0_isWr; // @[StreamArbiter.scala 25:22:@45841.4]
  wire [31:0] cmdMux_io_in_bits_0_tag; // @[StreamArbiter.scala 25:22:@45841.4]
  wire  cmdMux_io_out_ready; // @[StreamArbiter.scala 25:22:@45841.4]
  wire  cmdMux_io_out_valid; // @[StreamArbiter.scala 25:22:@45841.4]
  wire [63:0] cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 25:22:@45841.4]
  wire [31:0] cmdMux_io_out_bits_size; // @[StreamArbiter.scala 25:22:@45841.4]
  wire  cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 25:22:@45841.4]
  wire [31:0] cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 25:22:@45841.4]
  wire  wdataMux_io_in_ready; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_valid; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_0; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_1; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_2; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_3; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_4; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_5; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_6; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_7; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_8; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_9; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_10; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_11; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_12; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_13; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_14; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_in_bits_0_wdata_15; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_0; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_1; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_2; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_3; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_4; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_5; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_6; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_7; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_8; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_9; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_10; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_11; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_12; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_13; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_14; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_15; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_16; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_17; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_18; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_19; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_20; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_21; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_22; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_23; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_24; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_25; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_26; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_27; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_28; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_29; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_30; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_31; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_32; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_33; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_34; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_35; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_36; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_37; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_38; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_39; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_40; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_41; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_42; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_43; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_44; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_45; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_46; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_47; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_48; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_49; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_50; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_51; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_52; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_53; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_54; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_55; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_56; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_57; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_58; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_59; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_60; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_61; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_62; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_in_bits_0_wstrb_63; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_ready; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_valid; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 35:24:@45864.4]
  wire [31:0] wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 35:24:@45864.4]
  wire  elementCtr_clock; // @[StreamArbiter.scala 36:26:@45867.4]
  wire  elementCtr_reset; // @[StreamArbiter.scala 36:26:@45867.4]
  wire  elementCtr_io_reset; // @[StreamArbiter.scala 36:26:@45867.4]
  wire  elementCtr_io_enable; // @[StreamArbiter.scala 36:26:@45867.4]
  wire [31:0] elementCtr_io_out; // @[StreamArbiter.scala 36:26:@45867.4]
  wire  _T_346; // @[package.scala 96:25:@45836.4 package.scala 96:25:@45837.4]
  wire  cmdIdx; // @[StreamArbiter.scala 21:16:@45838.4]
  wire [1:0] cmdInDecoder; // @[OneHot.scala 45:35:@45840.4]
  wire  _T_355; // @[FringeBundles.scala 114:28:@45856.4]
  wire [22:0] _T_356; // @[FringeBundles.scala 114:28:@45858.4]
  wire [23:0] _T_358; // @[FringeBundles.scala 115:37:@45861.4]
  wire  _T_360; // @[StreamArbiter.scala 37:49:@45870.4]
  wire [31:0] _T_365; // @[:@45874.4 :@45875.4]
  wire [7:0] _T_366; // @[FringeBundles.scala 114:28:@45876.4]
  wire [255:0] cmdOutDecoder; // @[OneHot.scala 45:35:@45882.4]
  wire  _T_379; // @[StreamArbiter.scala 42:78:@45885.4]
  wire  _T_380; // @[StreamArbiter.scala 42:121:@45886.4]
  wire [7:0] _T_395; // @[FringeBundles.scala 140:28:@46073.4]
  wire [255:0] wrespDecoder; // @[OneHot.scala 45:35:@46080.4]
  wire  _T_400; // @[StreamArbiter.scala 61:55:@46085.4]
  wire  _T_403; // @[StreamArbiter.scala 62:85:@46089.4]
  wire  _T_404; // @[StreamArbiter.scala 62:70:@46090.4]
  wire  _T_409; // @[StreamArbiter.scala 67:58:@46114.4]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@45824.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  RetimeWrapper RetimeWrapper_1 ( // @[package.scala 93:22:@45831.4]
    .clock(RetimeWrapper_1_clock),
    .reset(RetimeWrapper_1_reset),
    .io_flow(RetimeWrapper_1_io_flow),
    .io_in(RetimeWrapper_1_io_in),
    .io_out(RetimeWrapper_1_io_out)
  );
  MuxPipe cmdMux ( // @[StreamArbiter.scala 25:22:@45841.4]
    .io_in_ready(cmdMux_io_in_ready),
    .io_in_valid(cmdMux_io_in_valid),
    .io_in_bits_0_addr(cmdMux_io_in_bits_0_addr),
    .io_in_bits_0_size(cmdMux_io_in_bits_0_size),
    .io_in_bits_0_isWr(cmdMux_io_in_bits_0_isWr),
    .io_in_bits_0_tag(cmdMux_io_in_bits_0_tag),
    .io_out_ready(cmdMux_io_out_ready),
    .io_out_valid(cmdMux_io_out_valid),
    .io_out_bits_addr(cmdMux_io_out_bits_addr),
    .io_out_bits_size(cmdMux_io_out_bits_size),
    .io_out_bits_isWr(cmdMux_io_out_bits_isWr),
    .io_out_bits_tag(cmdMux_io_out_bits_tag)
  );
  MuxPipe_1 wdataMux ( // @[StreamArbiter.scala 35:24:@45864.4]
    .io_in_ready(wdataMux_io_in_ready),
    .io_in_valid(wdataMux_io_in_valid),
    .io_in_bits_0_wdata_0(wdataMux_io_in_bits_0_wdata_0),
    .io_in_bits_0_wdata_1(wdataMux_io_in_bits_0_wdata_1),
    .io_in_bits_0_wdata_2(wdataMux_io_in_bits_0_wdata_2),
    .io_in_bits_0_wdata_3(wdataMux_io_in_bits_0_wdata_3),
    .io_in_bits_0_wdata_4(wdataMux_io_in_bits_0_wdata_4),
    .io_in_bits_0_wdata_5(wdataMux_io_in_bits_0_wdata_5),
    .io_in_bits_0_wdata_6(wdataMux_io_in_bits_0_wdata_6),
    .io_in_bits_0_wdata_7(wdataMux_io_in_bits_0_wdata_7),
    .io_in_bits_0_wdata_8(wdataMux_io_in_bits_0_wdata_8),
    .io_in_bits_0_wdata_9(wdataMux_io_in_bits_0_wdata_9),
    .io_in_bits_0_wdata_10(wdataMux_io_in_bits_0_wdata_10),
    .io_in_bits_0_wdata_11(wdataMux_io_in_bits_0_wdata_11),
    .io_in_bits_0_wdata_12(wdataMux_io_in_bits_0_wdata_12),
    .io_in_bits_0_wdata_13(wdataMux_io_in_bits_0_wdata_13),
    .io_in_bits_0_wdata_14(wdataMux_io_in_bits_0_wdata_14),
    .io_in_bits_0_wdata_15(wdataMux_io_in_bits_0_wdata_15),
    .io_in_bits_0_wstrb_0(wdataMux_io_in_bits_0_wstrb_0),
    .io_in_bits_0_wstrb_1(wdataMux_io_in_bits_0_wstrb_1),
    .io_in_bits_0_wstrb_2(wdataMux_io_in_bits_0_wstrb_2),
    .io_in_bits_0_wstrb_3(wdataMux_io_in_bits_0_wstrb_3),
    .io_in_bits_0_wstrb_4(wdataMux_io_in_bits_0_wstrb_4),
    .io_in_bits_0_wstrb_5(wdataMux_io_in_bits_0_wstrb_5),
    .io_in_bits_0_wstrb_6(wdataMux_io_in_bits_0_wstrb_6),
    .io_in_bits_0_wstrb_7(wdataMux_io_in_bits_0_wstrb_7),
    .io_in_bits_0_wstrb_8(wdataMux_io_in_bits_0_wstrb_8),
    .io_in_bits_0_wstrb_9(wdataMux_io_in_bits_0_wstrb_9),
    .io_in_bits_0_wstrb_10(wdataMux_io_in_bits_0_wstrb_10),
    .io_in_bits_0_wstrb_11(wdataMux_io_in_bits_0_wstrb_11),
    .io_in_bits_0_wstrb_12(wdataMux_io_in_bits_0_wstrb_12),
    .io_in_bits_0_wstrb_13(wdataMux_io_in_bits_0_wstrb_13),
    .io_in_bits_0_wstrb_14(wdataMux_io_in_bits_0_wstrb_14),
    .io_in_bits_0_wstrb_15(wdataMux_io_in_bits_0_wstrb_15),
    .io_in_bits_0_wstrb_16(wdataMux_io_in_bits_0_wstrb_16),
    .io_in_bits_0_wstrb_17(wdataMux_io_in_bits_0_wstrb_17),
    .io_in_bits_0_wstrb_18(wdataMux_io_in_bits_0_wstrb_18),
    .io_in_bits_0_wstrb_19(wdataMux_io_in_bits_0_wstrb_19),
    .io_in_bits_0_wstrb_20(wdataMux_io_in_bits_0_wstrb_20),
    .io_in_bits_0_wstrb_21(wdataMux_io_in_bits_0_wstrb_21),
    .io_in_bits_0_wstrb_22(wdataMux_io_in_bits_0_wstrb_22),
    .io_in_bits_0_wstrb_23(wdataMux_io_in_bits_0_wstrb_23),
    .io_in_bits_0_wstrb_24(wdataMux_io_in_bits_0_wstrb_24),
    .io_in_bits_0_wstrb_25(wdataMux_io_in_bits_0_wstrb_25),
    .io_in_bits_0_wstrb_26(wdataMux_io_in_bits_0_wstrb_26),
    .io_in_bits_0_wstrb_27(wdataMux_io_in_bits_0_wstrb_27),
    .io_in_bits_0_wstrb_28(wdataMux_io_in_bits_0_wstrb_28),
    .io_in_bits_0_wstrb_29(wdataMux_io_in_bits_0_wstrb_29),
    .io_in_bits_0_wstrb_30(wdataMux_io_in_bits_0_wstrb_30),
    .io_in_bits_0_wstrb_31(wdataMux_io_in_bits_0_wstrb_31),
    .io_in_bits_0_wstrb_32(wdataMux_io_in_bits_0_wstrb_32),
    .io_in_bits_0_wstrb_33(wdataMux_io_in_bits_0_wstrb_33),
    .io_in_bits_0_wstrb_34(wdataMux_io_in_bits_0_wstrb_34),
    .io_in_bits_0_wstrb_35(wdataMux_io_in_bits_0_wstrb_35),
    .io_in_bits_0_wstrb_36(wdataMux_io_in_bits_0_wstrb_36),
    .io_in_bits_0_wstrb_37(wdataMux_io_in_bits_0_wstrb_37),
    .io_in_bits_0_wstrb_38(wdataMux_io_in_bits_0_wstrb_38),
    .io_in_bits_0_wstrb_39(wdataMux_io_in_bits_0_wstrb_39),
    .io_in_bits_0_wstrb_40(wdataMux_io_in_bits_0_wstrb_40),
    .io_in_bits_0_wstrb_41(wdataMux_io_in_bits_0_wstrb_41),
    .io_in_bits_0_wstrb_42(wdataMux_io_in_bits_0_wstrb_42),
    .io_in_bits_0_wstrb_43(wdataMux_io_in_bits_0_wstrb_43),
    .io_in_bits_0_wstrb_44(wdataMux_io_in_bits_0_wstrb_44),
    .io_in_bits_0_wstrb_45(wdataMux_io_in_bits_0_wstrb_45),
    .io_in_bits_0_wstrb_46(wdataMux_io_in_bits_0_wstrb_46),
    .io_in_bits_0_wstrb_47(wdataMux_io_in_bits_0_wstrb_47),
    .io_in_bits_0_wstrb_48(wdataMux_io_in_bits_0_wstrb_48),
    .io_in_bits_0_wstrb_49(wdataMux_io_in_bits_0_wstrb_49),
    .io_in_bits_0_wstrb_50(wdataMux_io_in_bits_0_wstrb_50),
    .io_in_bits_0_wstrb_51(wdataMux_io_in_bits_0_wstrb_51),
    .io_in_bits_0_wstrb_52(wdataMux_io_in_bits_0_wstrb_52),
    .io_in_bits_0_wstrb_53(wdataMux_io_in_bits_0_wstrb_53),
    .io_in_bits_0_wstrb_54(wdataMux_io_in_bits_0_wstrb_54),
    .io_in_bits_0_wstrb_55(wdataMux_io_in_bits_0_wstrb_55),
    .io_in_bits_0_wstrb_56(wdataMux_io_in_bits_0_wstrb_56),
    .io_in_bits_0_wstrb_57(wdataMux_io_in_bits_0_wstrb_57),
    .io_in_bits_0_wstrb_58(wdataMux_io_in_bits_0_wstrb_58),
    .io_in_bits_0_wstrb_59(wdataMux_io_in_bits_0_wstrb_59),
    .io_in_bits_0_wstrb_60(wdataMux_io_in_bits_0_wstrb_60),
    .io_in_bits_0_wstrb_61(wdataMux_io_in_bits_0_wstrb_61),
    .io_in_bits_0_wstrb_62(wdataMux_io_in_bits_0_wstrb_62),
    .io_in_bits_0_wstrb_63(wdataMux_io_in_bits_0_wstrb_63),
    .io_out_ready(wdataMux_io_out_ready),
    .io_out_valid(wdataMux_io_out_valid),
    .io_out_bits_wdata_0(wdataMux_io_out_bits_wdata_0),
    .io_out_bits_wdata_1(wdataMux_io_out_bits_wdata_1),
    .io_out_bits_wdata_2(wdataMux_io_out_bits_wdata_2),
    .io_out_bits_wdata_3(wdataMux_io_out_bits_wdata_3),
    .io_out_bits_wdata_4(wdataMux_io_out_bits_wdata_4),
    .io_out_bits_wdata_5(wdataMux_io_out_bits_wdata_5),
    .io_out_bits_wdata_6(wdataMux_io_out_bits_wdata_6),
    .io_out_bits_wdata_7(wdataMux_io_out_bits_wdata_7),
    .io_out_bits_wdata_8(wdataMux_io_out_bits_wdata_8),
    .io_out_bits_wdata_9(wdataMux_io_out_bits_wdata_9),
    .io_out_bits_wdata_10(wdataMux_io_out_bits_wdata_10),
    .io_out_bits_wdata_11(wdataMux_io_out_bits_wdata_11),
    .io_out_bits_wdata_12(wdataMux_io_out_bits_wdata_12),
    .io_out_bits_wdata_13(wdataMux_io_out_bits_wdata_13),
    .io_out_bits_wdata_14(wdataMux_io_out_bits_wdata_14),
    .io_out_bits_wdata_15(wdataMux_io_out_bits_wdata_15),
    .io_out_bits_wstrb_0(wdataMux_io_out_bits_wstrb_0),
    .io_out_bits_wstrb_1(wdataMux_io_out_bits_wstrb_1),
    .io_out_bits_wstrb_2(wdataMux_io_out_bits_wstrb_2),
    .io_out_bits_wstrb_3(wdataMux_io_out_bits_wstrb_3),
    .io_out_bits_wstrb_4(wdataMux_io_out_bits_wstrb_4),
    .io_out_bits_wstrb_5(wdataMux_io_out_bits_wstrb_5),
    .io_out_bits_wstrb_6(wdataMux_io_out_bits_wstrb_6),
    .io_out_bits_wstrb_7(wdataMux_io_out_bits_wstrb_7),
    .io_out_bits_wstrb_8(wdataMux_io_out_bits_wstrb_8),
    .io_out_bits_wstrb_9(wdataMux_io_out_bits_wstrb_9),
    .io_out_bits_wstrb_10(wdataMux_io_out_bits_wstrb_10),
    .io_out_bits_wstrb_11(wdataMux_io_out_bits_wstrb_11),
    .io_out_bits_wstrb_12(wdataMux_io_out_bits_wstrb_12),
    .io_out_bits_wstrb_13(wdataMux_io_out_bits_wstrb_13),
    .io_out_bits_wstrb_14(wdataMux_io_out_bits_wstrb_14),
    .io_out_bits_wstrb_15(wdataMux_io_out_bits_wstrb_15),
    .io_out_bits_wstrb_16(wdataMux_io_out_bits_wstrb_16),
    .io_out_bits_wstrb_17(wdataMux_io_out_bits_wstrb_17),
    .io_out_bits_wstrb_18(wdataMux_io_out_bits_wstrb_18),
    .io_out_bits_wstrb_19(wdataMux_io_out_bits_wstrb_19),
    .io_out_bits_wstrb_20(wdataMux_io_out_bits_wstrb_20),
    .io_out_bits_wstrb_21(wdataMux_io_out_bits_wstrb_21),
    .io_out_bits_wstrb_22(wdataMux_io_out_bits_wstrb_22),
    .io_out_bits_wstrb_23(wdataMux_io_out_bits_wstrb_23),
    .io_out_bits_wstrb_24(wdataMux_io_out_bits_wstrb_24),
    .io_out_bits_wstrb_25(wdataMux_io_out_bits_wstrb_25),
    .io_out_bits_wstrb_26(wdataMux_io_out_bits_wstrb_26),
    .io_out_bits_wstrb_27(wdataMux_io_out_bits_wstrb_27),
    .io_out_bits_wstrb_28(wdataMux_io_out_bits_wstrb_28),
    .io_out_bits_wstrb_29(wdataMux_io_out_bits_wstrb_29),
    .io_out_bits_wstrb_30(wdataMux_io_out_bits_wstrb_30),
    .io_out_bits_wstrb_31(wdataMux_io_out_bits_wstrb_31),
    .io_out_bits_wstrb_32(wdataMux_io_out_bits_wstrb_32),
    .io_out_bits_wstrb_33(wdataMux_io_out_bits_wstrb_33),
    .io_out_bits_wstrb_34(wdataMux_io_out_bits_wstrb_34),
    .io_out_bits_wstrb_35(wdataMux_io_out_bits_wstrb_35),
    .io_out_bits_wstrb_36(wdataMux_io_out_bits_wstrb_36),
    .io_out_bits_wstrb_37(wdataMux_io_out_bits_wstrb_37),
    .io_out_bits_wstrb_38(wdataMux_io_out_bits_wstrb_38),
    .io_out_bits_wstrb_39(wdataMux_io_out_bits_wstrb_39),
    .io_out_bits_wstrb_40(wdataMux_io_out_bits_wstrb_40),
    .io_out_bits_wstrb_41(wdataMux_io_out_bits_wstrb_41),
    .io_out_bits_wstrb_42(wdataMux_io_out_bits_wstrb_42),
    .io_out_bits_wstrb_43(wdataMux_io_out_bits_wstrb_43),
    .io_out_bits_wstrb_44(wdataMux_io_out_bits_wstrb_44),
    .io_out_bits_wstrb_45(wdataMux_io_out_bits_wstrb_45),
    .io_out_bits_wstrb_46(wdataMux_io_out_bits_wstrb_46),
    .io_out_bits_wstrb_47(wdataMux_io_out_bits_wstrb_47),
    .io_out_bits_wstrb_48(wdataMux_io_out_bits_wstrb_48),
    .io_out_bits_wstrb_49(wdataMux_io_out_bits_wstrb_49),
    .io_out_bits_wstrb_50(wdataMux_io_out_bits_wstrb_50),
    .io_out_bits_wstrb_51(wdataMux_io_out_bits_wstrb_51),
    .io_out_bits_wstrb_52(wdataMux_io_out_bits_wstrb_52),
    .io_out_bits_wstrb_53(wdataMux_io_out_bits_wstrb_53),
    .io_out_bits_wstrb_54(wdataMux_io_out_bits_wstrb_54),
    .io_out_bits_wstrb_55(wdataMux_io_out_bits_wstrb_55),
    .io_out_bits_wstrb_56(wdataMux_io_out_bits_wstrb_56),
    .io_out_bits_wstrb_57(wdataMux_io_out_bits_wstrb_57),
    .io_out_bits_wstrb_58(wdataMux_io_out_bits_wstrb_58),
    .io_out_bits_wstrb_59(wdataMux_io_out_bits_wstrb_59),
    .io_out_bits_wstrb_60(wdataMux_io_out_bits_wstrb_60),
    .io_out_bits_wstrb_61(wdataMux_io_out_bits_wstrb_61),
    .io_out_bits_wstrb_62(wdataMux_io_out_bits_wstrb_62),
    .io_out_bits_wstrb_63(wdataMux_io_out_bits_wstrb_63)
  );
  ElementCounter elementCtr ( // @[StreamArbiter.scala 36:26:@45867.4]
    .clock(elementCtr_clock),
    .reset(elementCtr_reset),
    .io_reset(elementCtr_io_reset),
    .io_enable(elementCtr_io_enable),
    .io_out(elementCtr_io_out)
  );
  assign _T_346 = RetimeWrapper_1_io_out; // @[package.scala 96:25:@45836.4 package.scala 96:25:@45837.4]
  assign cmdIdx = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[StreamArbiter.scala 21:16:@45838.4]
  assign cmdInDecoder = 2'h1 << cmdIdx; // @[OneHot.scala 45:35:@45840.4]
  assign _T_355 = io_app_0_cmd_bits_tag[8]; // @[FringeBundles.scala 114:28:@45856.4]
  assign _T_356 = io_app_0_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@45858.4]
  assign _T_358 = {_T_356,_T_355}; // @[FringeBundles.scala 115:37:@45861.4]
  assign _T_360 = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:49:@45870.4]
  assign _T_365 = cmdMux_io_out_bits_tag; // @[:@45874.4 :@45875.4]
  assign _T_366 = _T_365[7:0]; // @[FringeBundles.scala 114:28:@45876.4]
  assign cmdOutDecoder = 256'h1 << _T_366; // @[OneHot.scala 45:35:@45882.4]
  assign _T_379 = io_app_0_wdata_valid & cmdMux_io_out_valid; // @[StreamArbiter.scala 42:78:@45885.4]
  assign _T_380 = elementCtr_io_out < cmdMux_io_out_bits_size; // @[StreamArbiter.scala 42:121:@45886.4]
  assign _T_395 = io_dram_wresp_bits_tag[7:0]; // @[FringeBundles.scala 140:28:@46073.4]
  assign wrespDecoder = 256'h1 << _T_395; // @[OneHot.scala 45:35:@46080.4]
  assign _T_400 = cmdInDecoder[0]; // @[StreamArbiter.scala 61:55:@46085.4]
  assign _T_403 = cmdOutDecoder[0]; // @[StreamArbiter.scala 62:85:@46089.4]
  assign _T_404 = _T_360 & _T_403; // @[StreamArbiter.scala 62:70:@46090.4]
  assign _T_409 = wrespDecoder[0]; // @[StreamArbiter.scala 67:58:@46114.4]
  assign io_app_0_cmd_ready = cmdMux_io_in_ready & _T_400; // @[StreamArbiter.scala 61:19:@46087.4]
  assign io_app_0_wdata_ready = _T_404 & _T_380; // @[StreamArbiter.scala 62:21:@46093.4]
  assign io_app_0_wresp_valid = io_dram_wresp_valid & _T_409; // @[StreamArbiter.scala 67:21:@46116.4]
  assign io_dram_cmd_valid = cmdMux_io_out_valid; // @[StreamArbiter.scala 46:15:@45976.4]
  assign io_dram_cmd_bits_addr = cmdMux_io_out_bits_addr; // @[StreamArbiter.scala 46:15:@45975.4]
  assign io_dram_cmd_bits_size = cmdMux_io_out_bits_size; // @[StreamArbiter.scala 46:15:@45974.4]
  assign io_dram_cmd_bits_isWr = cmdMux_io_out_bits_isWr; // @[StreamArbiter.scala 46:15:@45972.4]
  assign io_dram_cmd_bits_tag = cmdMux_io_out_bits_tag; // @[StreamArbiter.scala 46:15:@45971.4]
  assign io_dram_wdata_valid = wdataMux_io_out_valid; // @[StreamArbiter.scala 47:17:@46059.4]
  assign io_dram_wdata_bits_wdata_0 = wdataMux_io_out_bits_wdata_0; // @[StreamArbiter.scala 47:17:@46043.4]
  assign io_dram_wdata_bits_wdata_1 = wdataMux_io_out_bits_wdata_1; // @[StreamArbiter.scala 47:17:@46044.4]
  assign io_dram_wdata_bits_wdata_2 = wdataMux_io_out_bits_wdata_2; // @[StreamArbiter.scala 47:17:@46045.4]
  assign io_dram_wdata_bits_wdata_3 = wdataMux_io_out_bits_wdata_3; // @[StreamArbiter.scala 47:17:@46046.4]
  assign io_dram_wdata_bits_wdata_4 = wdataMux_io_out_bits_wdata_4; // @[StreamArbiter.scala 47:17:@46047.4]
  assign io_dram_wdata_bits_wdata_5 = wdataMux_io_out_bits_wdata_5; // @[StreamArbiter.scala 47:17:@46048.4]
  assign io_dram_wdata_bits_wdata_6 = wdataMux_io_out_bits_wdata_6; // @[StreamArbiter.scala 47:17:@46049.4]
  assign io_dram_wdata_bits_wdata_7 = wdataMux_io_out_bits_wdata_7; // @[StreamArbiter.scala 47:17:@46050.4]
  assign io_dram_wdata_bits_wdata_8 = wdataMux_io_out_bits_wdata_8; // @[StreamArbiter.scala 47:17:@46051.4]
  assign io_dram_wdata_bits_wdata_9 = wdataMux_io_out_bits_wdata_9; // @[StreamArbiter.scala 47:17:@46052.4]
  assign io_dram_wdata_bits_wdata_10 = wdataMux_io_out_bits_wdata_10; // @[StreamArbiter.scala 47:17:@46053.4]
  assign io_dram_wdata_bits_wdata_11 = wdataMux_io_out_bits_wdata_11; // @[StreamArbiter.scala 47:17:@46054.4]
  assign io_dram_wdata_bits_wdata_12 = wdataMux_io_out_bits_wdata_12; // @[StreamArbiter.scala 47:17:@46055.4]
  assign io_dram_wdata_bits_wdata_13 = wdataMux_io_out_bits_wdata_13; // @[StreamArbiter.scala 47:17:@46056.4]
  assign io_dram_wdata_bits_wdata_14 = wdataMux_io_out_bits_wdata_14; // @[StreamArbiter.scala 47:17:@46057.4]
  assign io_dram_wdata_bits_wdata_15 = wdataMux_io_out_bits_wdata_15; // @[StreamArbiter.scala 47:17:@46058.4]
  assign io_dram_wdata_bits_wstrb_0 = wdataMux_io_out_bits_wstrb_0; // @[StreamArbiter.scala 47:17:@45979.4]
  assign io_dram_wdata_bits_wstrb_1 = wdataMux_io_out_bits_wstrb_1; // @[StreamArbiter.scala 47:17:@45980.4]
  assign io_dram_wdata_bits_wstrb_2 = wdataMux_io_out_bits_wstrb_2; // @[StreamArbiter.scala 47:17:@45981.4]
  assign io_dram_wdata_bits_wstrb_3 = wdataMux_io_out_bits_wstrb_3; // @[StreamArbiter.scala 47:17:@45982.4]
  assign io_dram_wdata_bits_wstrb_4 = wdataMux_io_out_bits_wstrb_4; // @[StreamArbiter.scala 47:17:@45983.4]
  assign io_dram_wdata_bits_wstrb_5 = wdataMux_io_out_bits_wstrb_5; // @[StreamArbiter.scala 47:17:@45984.4]
  assign io_dram_wdata_bits_wstrb_6 = wdataMux_io_out_bits_wstrb_6; // @[StreamArbiter.scala 47:17:@45985.4]
  assign io_dram_wdata_bits_wstrb_7 = wdataMux_io_out_bits_wstrb_7; // @[StreamArbiter.scala 47:17:@45986.4]
  assign io_dram_wdata_bits_wstrb_8 = wdataMux_io_out_bits_wstrb_8; // @[StreamArbiter.scala 47:17:@45987.4]
  assign io_dram_wdata_bits_wstrb_9 = wdataMux_io_out_bits_wstrb_9; // @[StreamArbiter.scala 47:17:@45988.4]
  assign io_dram_wdata_bits_wstrb_10 = wdataMux_io_out_bits_wstrb_10; // @[StreamArbiter.scala 47:17:@45989.4]
  assign io_dram_wdata_bits_wstrb_11 = wdataMux_io_out_bits_wstrb_11; // @[StreamArbiter.scala 47:17:@45990.4]
  assign io_dram_wdata_bits_wstrb_12 = wdataMux_io_out_bits_wstrb_12; // @[StreamArbiter.scala 47:17:@45991.4]
  assign io_dram_wdata_bits_wstrb_13 = wdataMux_io_out_bits_wstrb_13; // @[StreamArbiter.scala 47:17:@45992.4]
  assign io_dram_wdata_bits_wstrb_14 = wdataMux_io_out_bits_wstrb_14; // @[StreamArbiter.scala 47:17:@45993.4]
  assign io_dram_wdata_bits_wstrb_15 = wdataMux_io_out_bits_wstrb_15; // @[StreamArbiter.scala 47:17:@45994.4]
  assign io_dram_wdata_bits_wstrb_16 = wdataMux_io_out_bits_wstrb_16; // @[StreamArbiter.scala 47:17:@45995.4]
  assign io_dram_wdata_bits_wstrb_17 = wdataMux_io_out_bits_wstrb_17; // @[StreamArbiter.scala 47:17:@45996.4]
  assign io_dram_wdata_bits_wstrb_18 = wdataMux_io_out_bits_wstrb_18; // @[StreamArbiter.scala 47:17:@45997.4]
  assign io_dram_wdata_bits_wstrb_19 = wdataMux_io_out_bits_wstrb_19; // @[StreamArbiter.scala 47:17:@45998.4]
  assign io_dram_wdata_bits_wstrb_20 = wdataMux_io_out_bits_wstrb_20; // @[StreamArbiter.scala 47:17:@45999.4]
  assign io_dram_wdata_bits_wstrb_21 = wdataMux_io_out_bits_wstrb_21; // @[StreamArbiter.scala 47:17:@46000.4]
  assign io_dram_wdata_bits_wstrb_22 = wdataMux_io_out_bits_wstrb_22; // @[StreamArbiter.scala 47:17:@46001.4]
  assign io_dram_wdata_bits_wstrb_23 = wdataMux_io_out_bits_wstrb_23; // @[StreamArbiter.scala 47:17:@46002.4]
  assign io_dram_wdata_bits_wstrb_24 = wdataMux_io_out_bits_wstrb_24; // @[StreamArbiter.scala 47:17:@46003.4]
  assign io_dram_wdata_bits_wstrb_25 = wdataMux_io_out_bits_wstrb_25; // @[StreamArbiter.scala 47:17:@46004.4]
  assign io_dram_wdata_bits_wstrb_26 = wdataMux_io_out_bits_wstrb_26; // @[StreamArbiter.scala 47:17:@46005.4]
  assign io_dram_wdata_bits_wstrb_27 = wdataMux_io_out_bits_wstrb_27; // @[StreamArbiter.scala 47:17:@46006.4]
  assign io_dram_wdata_bits_wstrb_28 = wdataMux_io_out_bits_wstrb_28; // @[StreamArbiter.scala 47:17:@46007.4]
  assign io_dram_wdata_bits_wstrb_29 = wdataMux_io_out_bits_wstrb_29; // @[StreamArbiter.scala 47:17:@46008.4]
  assign io_dram_wdata_bits_wstrb_30 = wdataMux_io_out_bits_wstrb_30; // @[StreamArbiter.scala 47:17:@46009.4]
  assign io_dram_wdata_bits_wstrb_31 = wdataMux_io_out_bits_wstrb_31; // @[StreamArbiter.scala 47:17:@46010.4]
  assign io_dram_wdata_bits_wstrb_32 = wdataMux_io_out_bits_wstrb_32; // @[StreamArbiter.scala 47:17:@46011.4]
  assign io_dram_wdata_bits_wstrb_33 = wdataMux_io_out_bits_wstrb_33; // @[StreamArbiter.scala 47:17:@46012.4]
  assign io_dram_wdata_bits_wstrb_34 = wdataMux_io_out_bits_wstrb_34; // @[StreamArbiter.scala 47:17:@46013.4]
  assign io_dram_wdata_bits_wstrb_35 = wdataMux_io_out_bits_wstrb_35; // @[StreamArbiter.scala 47:17:@46014.4]
  assign io_dram_wdata_bits_wstrb_36 = wdataMux_io_out_bits_wstrb_36; // @[StreamArbiter.scala 47:17:@46015.4]
  assign io_dram_wdata_bits_wstrb_37 = wdataMux_io_out_bits_wstrb_37; // @[StreamArbiter.scala 47:17:@46016.4]
  assign io_dram_wdata_bits_wstrb_38 = wdataMux_io_out_bits_wstrb_38; // @[StreamArbiter.scala 47:17:@46017.4]
  assign io_dram_wdata_bits_wstrb_39 = wdataMux_io_out_bits_wstrb_39; // @[StreamArbiter.scala 47:17:@46018.4]
  assign io_dram_wdata_bits_wstrb_40 = wdataMux_io_out_bits_wstrb_40; // @[StreamArbiter.scala 47:17:@46019.4]
  assign io_dram_wdata_bits_wstrb_41 = wdataMux_io_out_bits_wstrb_41; // @[StreamArbiter.scala 47:17:@46020.4]
  assign io_dram_wdata_bits_wstrb_42 = wdataMux_io_out_bits_wstrb_42; // @[StreamArbiter.scala 47:17:@46021.4]
  assign io_dram_wdata_bits_wstrb_43 = wdataMux_io_out_bits_wstrb_43; // @[StreamArbiter.scala 47:17:@46022.4]
  assign io_dram_wdata_bits_wstrb_44 = wdataMux_io_out_bits_wstrb_44; // @[StreamArbiter.scala 47:17:@46023.4]
  assign io_dram_wdata_bits_wstrb_45 = wdataMux_io_out_bits_wstrb_45; // @[StreamArbiter.scala 47:17:@46024.4]
  assign io_dram_wdata_bits_wstrb_46 = wdataMux_io_out_bits_wstrb_46; // @[StreamArbiter.scala 47:17:@46025.4]
  assign io_dram_wdata_bits_wstrb_47 = wdataMux_io_out_bits_wstrb_47; // @[StreamArbiter.scala 47:17:@46026.4]
  assign io_dram_wdata_bits_wstrb_48 = wdataMux_io_out_bits_wstrb_48; // @[StreamArbiter.scala 47:17:@46027.4]
  assign io_dram_wdata_bits_wstrb_49 = wdataMux_io_out_bits_wstrb_49; // @[StreamArbiter.scala 47:17:@46028.4]
  assign io_dram_wdata_bits_wstrb_50 = wdataMux_io_out_bits_wstrb_50; // @[StreamArbiter.scala 47:17:@46029.4]
  assign io_dram_wdata_bits_wstrb_51 = wdataMux_io_out_bits_wstrb_51; // @[StreamArbiter.scala 47:17:@46030.4]
  assign io_dram_wdata_bits_wstrb_52 = wdataMux_io_out_bits_wstrb_52; // @[StreamArbiter.scala 47:17:@46031.4]
  assign io_dram_wdata_bits_wstrb_53 = wdataMux_io_out_bits_wstrb_53; // @[StreamArbiter.scala 47:17:@46032.4]
  assign io_dram_wdata_bits_wstrb_54 = wdataMux_io_out_bits_wstrb_54; // @[StreamArbiter.scala 47:17:@46033.4]
  assign io_dram_wdata_bits_wstrb_55 = wdataMux_io_out_bits_wstrb_55; // @[StreamArbiter.scala 47:17:@46034.4]
  assign io_dram_wdata_bits_wstrb_56 = wdataMux_io_out_bits_wstrb_56; // @[StreamArbiter.scala 47:17:@46035.4]
  assign io_dram_wdata_bits_wstrb_57 = wdataMux_io_out_bits_wstrb_57; // @[StreamArbiter.scala 47:17:@46036.4]
  assign io_dram_wdata_bits_wstrb_58 = wdataMux_io_out_bits_wstrb_58; // @[StreamArbiter.scala 47:17:@46037.4]
  assign io_dram_wdata_bits_wstrb_59 = wdataMux_io_out_bits_wstrb_59; // @[StreamArbiter.scala 47:17:@46038.4]
  assign io_dram_wdata_bits_wstrb_60 = wdataMux_io_out_bits_wstrb_60; // @[StreamArbiter.scala 47:17:@46039.4]
  assign io_dram_wdata_bits_wstrb_61 = wdataMux_io_out_bits_wstrb_61; // @[StreamArbiter.scala 47:17:@46040.4]
  assign io_dram_wdata_bits_wstrb_62 = wdataMux_io_out_bits_wstrb_62; // @[StreamArbiter.scala 47:17:@46041.4]
  assign io_dram_wdata_bits_wstrb_63 = wdataMux_io_out_bits_wstrb_63; // @[StreamArbiter.scala 47:17:@46042.4]
  assign io_dram_rresp_ready = io_app_0_rresp_ready; // @[StreamArbiter.scala 72:23:@46120.4]
  assign io_dram_wresp_ready = io_app_0_wresp_ready; // @[StreamArbiter.scala 73:23:@46123.4]
  assign RetimeWrapper_clock = clock; // @[:@45825.4]
  assign RetimeWrapper_reset = reset; // @[:@45826.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@45828.4]
  assign RetimeWrapper_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@45827.4]
  assign RetimeWrapper_1_clock = clock; // @[:@45832.4]
  assign RetimeWrapper_1_reset = reset; // @[:@45833.4]
  assign RetimeWrapper_1_io_flow = 1'h1; // @[package.scala 95:18:@45835.4]
  assign RetimeWrapper_1_io_in = io_app_0_cmd_valid ? _T_346 : 1'h0; // @[package.scala 94:16:@45834.4]
  assign cmdMux_io_in_valid = io_app_0_cmd_valid; // @[StreamArbiter.scala 26:22:@45844.4]
  assign cmdMux_io_in_bits_0_addr = io_app_0_cmd_bits_addr; // @[StreamArbiter.scala 29:9:@45850.4]
  assign cmdMux_io_in_bits_0_size = io_app_0_cmd_bits_size; // @[StreamArbiter.scala 29:9:@45849.4]
  assign cmdMux_io_in_bits_0_isWr = io_app_0_cmd_bits_isWr; // @[StreamArbiter.scala 29:9:@45847.4]
  assign cmdMux_io_in_bits_0_tag = {_T_358,8'h0}; // @[StreamArbiter.scala 29:9:@45846.4 FringeBundles.scala 115:32:@45863.4]
  assign cmdMux_io_out_ready = io_dram_cmd_valid & io_dram_cmd_ready; // @[StreamArbiter.scala 46:15:@45977.4 StreamArbiter.scala 57:23:@46083.4]
  assign wdataMux_io_in_valid = _T_379 & _T_380; // @[StreamArbiter.scala 42:24:@45888.4]
  assign wdataMux_io_in_bits_0_wdata_0 = io_app_0_wdata_bits_wdata_0; // @[StreamArbiter.scala 44:23:@45955.4]
  assign wdataMux_io_in_bits_0_wdata_1 = io_app_0_wdata_bits_wdata_1; // @[StreamArbiter.scala 44:23:@45956.4]
  assign wdataMux_io_in_bits_0_wdata_2 = io_app_0_wdata_bits_wdata_2; // @[StreamArbiter.scala 44:23:@45957.4]
  assign wdataMux_io_in_bits_0_wdata_3 = io_app_0_wdata_bits_wdata_3; // @[StreamArbiter.scala 44:23:@45958.4]
  assign wdataMux_io_in_bits_0_wdata_4 = io_app_0_wdata_bits_wdata_4; // @[StreamArbiter.scala 44:23:@45959.4]
  assign wdataMux_io_in_bits_0_wdata_5 = io_app_0_wdata_bits_wdata_5; // @[StreamArbiter.scala 44:23:@45960.4]
  assign wdataMux_io_in_bits_0_wdata_6 = io_app_0_wdata_bits_wdata_6; // @[StreamArbiter.scala 44:23:@45961.4]
  assign wdataMux_io_in_bits_0_wdata_7 = io_app_0_wdata_bits_wdata_7; // @[StreamArbiter.scala 44:23:@45962.4]
  assign wdataMux_io_in_bits_0_wdata_8 = io_app_0_wdata_bits_wdata_8; // @[StreamArbiter.scala 44:23:@45963.4]
  assign wdataMux_io_in_bits_0_wdata_9 = io_app_0_wdata_bits_wdata_9; // @[StreamArbiter.scala 44:23:@45964.4]
  assign wdataMux_io_in_bits_0_wdata_10 = io_app_0_wdata_bits_wdata_10; // @[StreamArbiter.scala 44:23:@45965.4]
  assign wdataMux_io_in_bits_0_wdata_11 = io_app_0_wdata_bits_wdata_11; // @[StreamArbiter.scala 44:23:@45966.4]
  assign wdataMux_io_in_bits_0_wdata_12 = io_app_0_wdata_bits_wdata_12; // @[StreamArbiter.scala 44:23:@45967.4]
  assign wdataMux_io_in_bits_0_wdata_13 = io_app_0_wdata_bits_wdata_13; // @[StreamArbiter.scala 44:23:@45968.4]
  assign wdataMux_io_in_bits_0_wdata_14 = io_app_0_wdata_bits_wdata_14; // @[StreamArbiter.scala 44:23:@45969.4]
  assign wdataMux_io_in_bits_0_wdata_15 = io_app_0_wdata_bits_wdata_15; // @[StreamArbiter.scala 44:23:@45970.4]
  assign wdataMux_io_in_bits_0_wstrb_0 = io_app_0_wdata_bits_wstrb_0; // @[StreamArbiter.scala 44:23:@45891.4]
  assign wdataMux_io_in_bits_0_wstrb_1 = io_app_0_wdata_bits_wstrb_1; // @[StreamArbiter.scala 44:23:@45892.4]
  assign wdataMux_io_in_bits_0_wstrb_2 = io_app_0_wdata_bits_wstrb_2; // @[StreamArbiter.scala 44:23:@45893.4]
  assign wdataMux_io_in_bits_0_wstrb_3 = io_app_0_wdata_bits_wstrb_3; // @[StreamArbiter.scala 44:23:@45894.4]
  assign wdataMux_io_in_bits_0_wstrb_4 = io_app_0_wdata_bits_wstrb_4; // @[StreamArbiter.scala 44:23:@45895.4]
  assign wdataMux_io_in_bits_0_wstrb_5 = io_app_0_wdata_bits_wstrb_5; // @[StreamArbiter.scala 44:23:@45896.4]
  assign wdataMux_io_in_bits_0_wstrb_6 = io_app_0_wdata_bits_wstrb_6; // @[StreamArbiter.scala 44:23:@45897.4]
  assign wdataMux_io_in_bits_0_wstrb_7 = io_app_0_wdata_bits_wstrb_7; // @[StreamArbiter.scala 44:23:@45898.4]
  assign wdataMux_io_in_bits_0_wstrb_8 = io_app_0_wdata_bits_wstrb_8; // @[StreamArbiter.scala 44:23:@45899.4]
  assign wdataMux_io_in_bits_0_wstrb_9 = io_app_0_wdata_bits_wstrb_9; // @[StreamArbiter.scala 44:23:@45900.4]
  assign wdataMux_io_in_bits_0_wstrb_10 = io_app_0_wdata_bits_wstrb_10; // @[StreamArbiter.scala 44:23:@45901.4]
  assign wdataMux_io_in_bits_0_wstrb_11 = io_app_0_wdata_bits_wstrb_11; // @[StreamArbiter.scala 44:23:@45902.4]
  assign wdataMux_io_in_bits_0_wstrb_12 = io_app_0_wdata_bits_wstrb_12; // @[StreamArbiter.scala 44:23:@45903.4]
  assign wdataMux_io_in_bits_0_wstrb_13 = io_app_0_wdata_bits_wstrb_13; // @[StreamArbiter.scala 44:23:@45904.4]
  assign wdataMux_io_in_bits_0_wstrb_14 = io_app_0_wdata_bits_wstrb_14; // @[StreamArbiter.scala 44:23:@45905.4]
  assign wdataMux_io_in_bits_0_wstrb_15 = io_app_0_wdata_bits_wstrb_15; // @[StreamArbiter.scala 44:23:@45906.4]
  assign wdataMux_io_in_bits_0_wstrb_16 = io_app_0_wdata_bits_wstrb_16; // @[StreamArbiter.scala 44:23:@45907.4]
  assign wdataMux_io_in_bits_0_wstrb_17 = io_app_0_wdata_bits_wstrb_17; // @[StreamArbiter.scala 44:23:@45908.4]
  assign wdataMux_io_in_bits_0_wstrb_18 = io_app_0_wdata_bits_wstrb_18; // @[StreamArbiter.scala 44:23:@45909.4]
  assign wdataMux_io_in_bits_0_wstrb_19 = io_app_0_wdata_bits_wstrb_19; // @[StreamArbiter.scala 44:23:@45910.4]
  assign wdataMux_io_in_bits_0_wstrb_20 = io_app_0_wdata_bits_wstrb_20; // @[StreamArbiter.scala 44:23:@45911.4]
  assign wdataMux_io_in_bits_0_wstrb_21 = io_app_0_wdata_bits_wstrb_21; // @[StreamArbiter.scala 44:23:@45912.4]
  assign wdataMux_io_in_bits_0_wstrb_22 = io_app_0_wdata_bits_wstrb_22; // @[StreamArbiter.scala 44:23:@45913.4]
  assign wdataMux_io_in_bits_0_wstrb_23 = io_app_0_wdata_bits_wstrb_23; // @[StreamArbiter.scala 44:23:@45914.4]
  assign wdataMux_io_in_bits_0_wstrb_24 = io_app_0_wdata_bits_wstrb_24; // @[StreamArbiter.scala 44:23:@45915.4]
  assign wdataMux_io_in_bits_0_wstrb_25 = io_app_0_wdata_bits_wstrb_25; // @[StreamArbiter.scala 44:23:@45916.4]
  assign wdataMux_io_in_bits_0_wstrb_26 = io_app_0_wdata_bits_wstrb_26; // @[StreamArbiter.scala 44:23:@45917.4]
  assign wdataMux_io_in_bits_0_wstrb_27 = io_app_0_wdata_bits_wstrb_27; // @[StreamArbiter.scala 44:23:@45918.4]
  assign wdataMux_io_in_bits_0_wstrb_28 = io_app_0_wdata_bits_wstrb_28; // @[StreamArbiter.scala 44:23:@45919.4]
  assign wdataMux_io_in_bits_0_wstrb_29 = io_app_0_wdata_bits_wstrb_29; // @[StreamArbiter.scala 44:23:@45920.4]
  assign wdataMux_io_in_bits_0_wstrb_30 = io_app_0_wdata_bits_wstrb_30; // @[StreamArbiter.scala 44:23:@45921.4]
  assign wdataMux_io_in_bits_0_wstrb_31 = io_app_0_wdata_bits_wstrb_31; // @[StreamArbiter.scala 44:23:@45922.4]
  assign wdataMux_io_in_bits_0_wstrb_32 = io_app_0_wdata_bits_wstrb_32; // @[StreamArbiter.scala 44:23:@45923.4]
  assign wdataMux_io_in_bits_0_wstrb_33 = io_app_0_wdata_bits_wstrb_33; // @[StreamArbiter.scala 44:23:@45924.4]
  assign wdataMux_io_in_bits_0_wstrb_34 = io_app_0_wdata_bits_wstrb_34; // @[StreamArbiter.scala 44:23:@45925.4]
  assign wdataMux_io_in_bits_0_wstrb_35 = io_app_0_wdata_bits_wstrb_35; // @[StreamArbiter.scala 44:23:@45926.4]
  assign wdataMux_io_in_bits_0_wstrb_36 = io_app_0_wdata_bits_wstrb_36; // @[StreamArbiter.scala 44:23:@45927.4]
  assign wdataMux_io_in_bits_0_wstrb_37 = io_app_0_wdata_bits_wstrb_37; // @[StreamArbiter.scala 44:23:@45928.4]
  assign wdataMux_io_in_bits_0_wstrb_38 = io_app_0_wdata_bits_wstrb_38; // @[StreamArbiter.scala 44:23:@45929.4]
  assign wdataMux_io_in_bits_0_wstrb_39 = io_app_0_wdata_bits_wstrb_39; // @[StreamArbiter.scala 44:23:@45930.4]
  assign wdataMux_io_in_bits_0_wstrb_40 = io_app_0_wdata_bits_wstrb_40; // @[StreamArbiter.scala 44:23:@45931.4]
  assign wdataMux_io_in_bits_0_wstrb_41 = io_app_0_wdata_bits_wstrb_41; // @[StreamArbiter.scala 44:23:@45932.4]
  assign wdataMux_io_in_bits_0_wstrb_42 = io_app_0_wdata_bits_wstrb_42; // @[StreamArbiter.scala 44:23:@45933.4]
  assign wdataMux_io_in_bits_0_wstrb_43 = io_app_0_wdata_bits_wstrb_43; // @[StreamArbiter.scala 44:23:@45934.4]
  assign wdataMux_io_in_bits_0_wstrb_44 = io_app_0_wdata_bits_wstrb_44; // @[StreamArbiter.scala 44:23:@45935.4]
  assign wdataMux_io_in_bits_0_wstrb_45 = io_app_0_wdata_bits_wstrb_45; // @[StreamArbiter.scala 44:23:@45936.4]
  assign wdataMux_io_in_bits_0_wstrb_46 = io_app_0_wdata_bits_wstrb_46; // @[StreamArbiter.scala 44:23:@45937.4]
  assign wdataMux_io_in_bits_0_wstrb_47 = io_app_0_wdata_bits_wstrb_47; // @[StreamArbiter.scala 44:23:@45938.4]
  assign wdataMux_io_in_bits_0_wstrb_48 = io_app_0_wdata_bits_wstrb_48; // @[StreamArbiter.scala 44:23:@45939.4]
  assign wdataMux_io_in_bits_0_wstrb_49 = io_app_0_wdata_bits_wstrb_49; // @[StreamArbiter.scala 44:23:@45940.4]
  assign wdataMux_io_in_bits_0_wstrb_50 = io_app_0_wdata_bits_wstrb_50; // @[StreamArbiter.scala 44:23:@45941.4]
  assign wdataMux_io_in_bits_0_wstrb_51 = io_app_0_wdata_bits_wstrb_51; // @[StreamArbiter.scala 44:23:@45942.4]
  assign wdataMux_io_in_bits_0_wstrb_52 = io_app_0_wdata_bits_wstrb_52; // @[StreamArbiter.scala 44:23:@45943.4]
  assign wdataMux_io_in_bits_0_wstrb_53 = io_app_0_wdata_bits_wstrb_53; // @[StreamArbiter.scala 44:23:@45944.4]
  assign wdataMux_io_in_bits_0_wstrb_54 = io_app_0_wdata_bits_wstrb_54; // @[StreamArbiter.scala 44:23:@45945.4]
  assign wdataMux_io_in_bits_0_wstrb_55 = io_app_0_wdata_bits_wstrb_55; // @[StreamArbiter.scala 44:23:@45946.4]
  assign wdataMux_io_in_bits_0_wstrb_56 = io_app_0_wdata_bits_wstrb_56; // @[StreamArbiter.scala 44:23:@45947.4]
  assign wdataMux_io_in_bits_0_wstrb_57 = io_app_0_wdata_bits_wstrb_57; // @[StreamArbiter.scala 44:23:@45948.4]
  assign wdataMux_io_in_bits_0_wstrb_58 = io_app_0_wdata_bits_wstrb_58; // @[StreamArbiter.scala 44:23:@45949.4]
  assign wdataMux_io_in_bits_0_wstrb_59 = io_app_0_wdata_bits_wstrb_59; // @[StreamArbiter.scala 44:23:@45950.4]
  assign wdataMux_io_in_bits_0_wstrb_60 = io_app_0_wdata_bits_wstrb_60; // @[StreamArbiter.scala 44:23:@45951.4]
  assign wdataMux_io_in_bits_0_wstrb_61 = io_app_0_wdata_bits_wstrb_61; // @[StreamArbiter.scala 44:23:@45952.4]
  assign wdataMux_io_in_bits_0_wstrb_62 = io_app_0_wdata_bits_wstrb_62; // @[StreamArbiter.scala 44:23:@45953.4]
  assign wdataMux_io_in_bits_0_wstrb_63 = io_app_0_wdata_bits_wstrb_63; // @[StreamArbiter.scala 44:23:@45954.4]
  assign wdataMux_io_out_ready = io_dram_wdata_valid & io_dram_wdata_ready; // @[StreamArbiter.scala 47:17:@46060.4 StreamArbiter.scala 58:25:@46084.4]
  assign elementCtr_clock = clock; // @[:@45868.4]
  assign elementCtr_reset = reset; // @[:@45869.4]
  assign elementCtr_io_reset = cmdMux_io_out_ready; // @[StreamArbiter.scala 38:23:@45872.4]
  assign elementCtr_io_enable = wdataMux_io_in_ready & wdataMux_io_in_valid; // @[StreamArbiter.scala 37:24:@45871.4]
endmodule
module Counter_72( // @[:@46125.2]
  input         clock, // @[:@46126.4]
  input         reset, // @[:@46127.4]
  input         io_reset, // @[:@46128.4]
  input         io_enable, // @[:@46128.4]
  input  [31:0] io_stride, // @[:@46128.4]
  output [31:0] io_out, // @[:@46128.4]
  output [31:0] io_next // @[:@46128.4]
);
  reg [31:0] count; // @[Counter.scala 15:22:@46130.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_17; // @[Counter.scala 17:24:@46131.4]
  wire [31:0] newCount; // @[Counter.scala 17:24:@46132.4]
  wire [31:0] _GEN_0; // @[Counter.scala 21:26:@46137.6]
  wire [31:0] _GEN_1; // @[Counter.scala 19:18:@46133.4]
  assign _T_17 = count + io_stride; // @[Counter.scala 17:24:@46131.4]
  assign newCount = count + io_stride; // @[Counter.scala 17:24:@46132.4]
  assign _GEN_0 = io_enable ? newCount : count; // @[Counter.scala 21:26:@46137.6]
  assign _GEN_1 = io_reset ? 32'h0 : _GEN_0; // @[Counter.scala 19:18:@46133.4]
  assign io_out = count; // @[Counter.scala 25:10:@46140.4]
  assign io_next = count + io_stride; // @[Counter.scala 26:11:@46141.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  count = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      count <= 32'h0;
    end else begin
      if (io_reset) begin
        count <= 32'h0;
      end else begin
        if (io_enable) begin
          count <= newCount;
        end
      end
    end
  end
endmodule
module AXICmdSplit( // @[:@46143.2]
  input         clock, // @[:@46144.4]
  input         reset, // @[:@46145.4]
  output        io_in_cmd_ready, // @[:@46146.4]
  input         io_in_cmd_valid, // @[:@46146.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@46146.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@46146.4]
  input         io_in_cmd_bits_isWr, // @[:@46146.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@46146.4]
  output        io_in_wdata_ready, // @[:@46146.4]
  input         io_in_wdata_valid, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@46146.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@46146.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@46146.4]
  input         io_in_rresp_ready, // @[:@46146.4]
  input         io_in_wresp_ready, // @[:@46146.4]
  output        io_in_wresp_valid, // @[:@46146.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@46146.4]
  input         io_out_cmd_ready, // @[:@46146.4]
  output        io_out_cmd_valid, // @[:@46146.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@46146.4]
  output [31:0] io_out_cmd_bits_size, // @[:@46146.4]
  output        io_out_cmd_bits_isWr, // @[:@46146.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@46146.4]
  input         io_out_wdata_ready, // @[:@46146.4]
  output        io_out_wdata_valid, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@46146.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@46146.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@46146.4]
  output        io_out_rresp_ready, // @[:@46146.4]
  output        io_out_wresp_ready, // @[:@46146.4]
  input         io_out_wresp_valid, // @[:@46146.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@46146.4]
);
  wire  cmdSizeCounter_clock; // @[AXIProtocol.scala 18:30:@46260.4]
  wire  cmdSizeCounter_reset; // @[AXIProtocol.scala 18:30:@46260.4]
  wire  cmdSizeCounter_io_reset; // @[AXIProtocol.scala 18:30:@46260.4]
  wire  cmdSizeCounter_io_enable; // @[AXIProtocol.scala 18:30:@46260.4]
  wire [31:0] cmdSizeCounter_io_stride; // @[AXIProtocol.scala 18:30:@46260.4]
  wire [31:0] cmdSizeCounter_io_out; // @[AXIProtocol.scala 18:30:@46260.4]
  wire [31:0] cmdSizeCounter_io_next; // @[AXIProtocol.scala 18:30:@46260.4]
  wire [32:0] _T_199; // @[AXIProtocol.scala 20:46:@46263.4]
  wire [32:0] _T_200; // @[AXIProtocol.scala 20:46:@46264.4]
  wire [31:0] cmdSizeRemaining; // @[AXIProtocol.scala 20:46:@46265.4]
  wire  lastCmd; // @[AXIProtocol.scala 23:35:@46266.4]
  wire [37:0] _GEN_0; // @[AXIProtocol.scala 27:47:@46269.4]
  wire [37:0] addrOffsetBytes; // @[AXIProtocol.scala 27:47:@46269.4]
  wire [63:0] _GEN_1; // @[AXIProtocol.scala 28:49:@46270.4]
  wire [64:0] _T_201; // @[AXIProtocol.scala 28:49:@46270.4]
  wire [63:0] cmdAddr_bits; // @[AXIProtocol.scala 28:49:@46271.4]
  wire [57:0] _T_204; // @[FringeBundles.scala 158:22:@46274.4]
  wire [7:0] cmdTag_streamID; // @[FringeBundles.scala 114:28:@46281.4]
  wire [22:0] cmdTag_uid; // @[FringeBundles.scala 114:28:@46285.4]
  wire [23:0] _T_214; // @[FringeBundles.scala 115:37:@46288.4]
  wire  cmdIssue; // @[AXIProtocol.scala 36:35:@46291.4]
  wire  _T_223; // @[FringeBundles.scala 140:28:@46302.4]
  Counter_72 cmdSizeCounter ( // @[AXIProtocol.scala 18:30:@46260.4]
    .clock(cmdSizeCounter_clock),
    .reset(cmdSizeCounter_reset),
    .io_reset(cmdSizeCounter_io_reset),
    .io_enable(cmdSizeCounter_io_enable),
    .io_stride(cmdSizeCounter_io_stride),
    .io_out(cmdSizeCounter_io_out),
    .io_next(cmdSizeCounter_io_next)
  );
  assign _T_199 = io_in_cmd_bits_size - cmdSizeCounter_io_out; // @[AXIProtocol.scala 20:46:@46263.4]
  assign _T_200 = $unsigned(_T_199); // @[AXIProtocol.scala 20:46:@46264.4]
  assign cmdSizeRemaining = _T_200[31:0]; // @[AXIProtocol.scala 20:46:@46265.4]
  assign lastCmd = cmdSizeRemaining <= 32'h100; // @[AXIProtocol.scala 23:35:@46266.4]
  assign _GEN_0 = {{6'd0}, cmdSizeCounter_io_out}; // @[AXIProtocol.scala 27:47:@46269.4]
  assign addrOffsetBytes = _GEN_0 << 6; // @[AXIProtocol.scala 27:47:@46269.4]
  assign _GEN_1 = {{26'd0}, addrOffsetBytes}; // @[AXIProtocol.scala 28:49:@46270.4]
  assign _T_201 = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@46270.4]
  assign cmdAddr_bits = io_in_cmd_bits_addr + _GEN_1; // @[AXIProtocol.scala 28:49:@46271.4]
  assign _T_204 = cmdAddr_bits[63:6]; // @[FringeBundles.scala 158:22:@46274.4]
  assign cmdTag_streamID = io_in_cmd_bits_tag[7:0]; // @[FringeBundles.scala 114:28:@46281.4]
  assign cmdTag_uid = io_in_cmd_bits_tag[31:9]; // @[FringeBundles.scala 114:28:@46285.4]
  assign _T_214 = {cmdTag_uid,lastCmd}; // @[FringeBundles.scala 115:37:@46288.4]
  assign cmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 36:35:@46291.4]
  assign _T_223 = io_out_wresp_bits_tag[8]; // @[FringeBundles.scala 140:28:@46302.4]
  assign io_in_cmd_ready = lastCmd & cmdIssue; // @[AXIProtocol.scala 15:10:@46259.4 AXIProtocol.scala 38:19:@46293.4]
  assign io_in_wdata_ready = io_out_wdata_ready; // @[AXIProtocol.scala 15:10:@46252.4]
  assign io_in_wresp_valid = io_out_wresp_valid & _T_223; // @[AXIProtocol.scala 15:10:@46149.4 AXIProtocol.scala 46:21:@46307.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 15:10:@46148.4]
  assign io_out_cmd_valid = io_in_cmd_valid; // @[AXIProtocol.scala 15:10:@46258.4]
  assign io_out_cmd_bits_addr = {_T_204,6'h0}; // @[AXIProtocol.scala 15:10:@46257.4 AXIProtocol.scala 29:24:@46276.4]
  assign io_out_cmd_bits_size = lastCmd ? cmdSizeRemaining : 32'h100; // @[AXIProtocol.scala 15:10:@46256.4 AXIProtocol.scala 25:24:@46268.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 15:10:@46254.4]
  assign io_out_cmd_bits_tag = {_T_214,cmdTag_streamID}; // @[AXIProtocol.scala 15:10:@46253.4 FringeBundles.scala 115:32:@46290.4]
  assign io_out_wdata_valid = io_in_wdata_valid; // @[AXIProtocol.scala 15:10:@46251.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 15:10:@46235.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 15:10:@46236.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 15:10:@46237.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 15:10:@46238.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 15:10:@46239.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 15:10:@46240.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 15:10:@46241.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 15:10:@46242.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 15:10:@46243.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 15:10:@46244.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 15:10:@46245.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 15:10:@46246.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 15:10:@46247.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 15:10:@46248.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 15:10:@46249.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 15:10:@46250.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 15:10:@46171.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 15:10:@46172.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 15:10:@46173.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 15:10:@46174.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 15:10:@46175.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 15:10:@46176.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 15:10:@46177.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 15:10:@46178.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 15:10:@46179.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 15:10:@46180.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 15:10:@46181.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 15:10:@46182.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 15:10:@46183.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 15:10:@46184.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 15:10:@46185.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 15:10:@46186.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 15:10:@46187.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 15:10:@46188.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 15:10:@46189.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 15:10:@46190.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 15:10:@46191.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 15:10:@46192.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 15:10:@46193.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 15:10:@46194.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 15:10:@46195.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 15:10:@46196.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 15:10:@46197.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 15:10:@46198.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 15:10:@46199.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 15:10:@46200.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 15:10:@46201.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 15:10:@46202.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 15:10:@46203.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 15:10:@46204.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 15:10:@46205.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 15:10:@46206.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 15:10:@46207.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 15:10:@46208.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 15:10:@46209.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 15:10:@46210.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 15:10:@46211.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 15:10:@46212.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 15:10:@46213.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 15:10:@46214.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 15:10:@46215.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 15:10:@46216.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 15:10:@46217.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 15:10:@46218.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 15:10:@46219.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 15:10:@46220.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 15:10:@46221.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 15:10:@46222.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 15:10:@46223.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 15:10:@46224.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 15:10:@46225.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 15:10:@46226.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 15:10:@46227.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 15:10:@46228.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 15:10:@46229.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 15:10:@46230.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 15:10:@46231.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 15:10:@46232.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 15:10:@46233.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 15:10:@46234.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 15:10:@46169.4]
  assign io_out_wresp_ready = _T_223 ? io_in_wresp_ready : 1'h1; // @[AXIProtocol.scala 15:10:@46150.4 AXIProtocol.scala 47:22:@46309.4]
  assign cmdSizeCounter_clock = clock; // @[:@46261.4]
  assign cmdSizeCounter_reset = reset; // @[:@46262.4]
  assign cmdSizeCounter_io_reset = lastCmd & cmdIssue; // @[AXIProtocol.scala 40:27:@46294.4]
  assign cmdSizeCounter_io_enable = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 41:28:@46295.4]
  assign cmdSizeCounter_io_stride = 32'h100; // @[AXIProtocol.scala 42:28:@46296.4]
endmodule
module AXICmdIssue( // @[:@46329.2]
  input         clock, // @[:@46330.4]
  input         reset, // @[:@46331.4]
  output        io_in_cmd_ready, // @[:@46332.4]
  input         io_in_cmd_valid, // @[:@46332.4]
  input  [63:0] io_in_cmd_bits_addr, // @[:@46332.4]
  input  [31:0] io_in_cmd_bits_size, // @[:@46332.4]
  input         io_in_cmd_bits_isWr, // @[:@46332.4]
  input  [31:0] io_in_cmd_bits_tag, // @[:@46332.4]
  output        io_in_wdata_ready, // @[:@46332.4]
  input         io_in_wdata_valid, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_0, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_1, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_2, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_3, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_4, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_5, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_6, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_7, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_8, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_9, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_10, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_11, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_12, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_13, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_14, // @[:@46332.4]
  input  [31:0] io_in_wdata_bits_wdata_15, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_0, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_1, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_2, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_3, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_4, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_5, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_6, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_7, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_8, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_9, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_10, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_11, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_12, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_13, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_14, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_15, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_16, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_17, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_18, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_19, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_20, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_21, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_22, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_23, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_24, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_25, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_26, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_27, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_28, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_29, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_30, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_31, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_32, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_33, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_34, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_35, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_36, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_37, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_38, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_39, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_40, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_41, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_42, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_43, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_44, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_45, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_46, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_47, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_48, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_49, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_50, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_51, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_52, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_53, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_54, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_55, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_56, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_57, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_58, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_59, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_60, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_61, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_62, // @[:@46332.4]
  input         io_in_wdata_bits_wstrb_63, // @[:@46332.4]
  input         io_in_rresp_ready, // @[:@46332.4]
  input         io_in_wresp_ready, // @[:@46332.4]
  output        io_in_wresp_valid, // @[:@46332.4]
  output [31:0] io_in_wresp_bits_tag, // @[:@46332.4]
  input         io_out_cmd_ready, // @[:@46332.4]
  output        io_out_cmd_valid, // @[:@46332.4]
  output [63:0] io_out_cmd_bits_addr, // @[:@46332.4]
  output [31:0] io_out_cmd_bits_size, // @[:@46332.4]
  output        io_out_cmd_bits_isWr, // @[:@46332.4]
  output [31:0] io_out_cmd_bits_tag, // @[:@46332.4]
  input         io_out_wdata_ready, // @[:@46332.4]
  output        io_out_wdata_valid, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_0, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_1, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_2, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_3, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_4, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_5, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_6, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_7, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_8, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_9, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_10, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_11, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_12, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_13, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_14, // @[:@46332.4]
  output [31:0] io_out_wdata_bits_wdata_15, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_0, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_1, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_2, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_3, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_4, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_5, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_6, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_7, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_8, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_9, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_10, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_11, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_12, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_13, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_14, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_15, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_16, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_17, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_18, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_19, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_20, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_21, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_22, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_23, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_24, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_25, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_26, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_27, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_28, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_29, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_30, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_31, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_32, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_33, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_34, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_35, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_36, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_37, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_38, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_39, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_40, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_41, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_42, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_43, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_44, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_45, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_46, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_47, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_48, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_49, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_50, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_51, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_52, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_53, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_54, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_55, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_56, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_57, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_58, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_59, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_60, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_61, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_62, // @[:@46332.4]
  output        io_out_wdata_bits_wstrb_63, // @[:@46332.4]
  output        io_out_wdata_bits_wlast, // @[:@46332.4]
  output        io_out_rresp_ready, // @[:@46332.4]
  output        io_out_wresp_ready, // @[:@46332.4]
  input         io_out_wresp_valid, // @[:@46332.4]
  input  [31:0] io_out_wresp_bits_tag // @[:@46332.4]
);
  wire  wdataCounter_clock; // @[AXIProtocol.scala 59:28:@46446.4]
  wire  wdataCounter_reset; // @[AXIProtocol.scala 59:28:@46446.4]
  wire  wdataCounter_io_reset; // @[AXIProtocol.scala 59:28:@46446.4]
  wire  wdataCounter_io_enable; // @[AXIProtocol.scala 59:28:@46446.4]
  wire [31:0] wdataCounter_io_stride; // @[AXIProtocol.scala 59:28:@46446.4]
  wire [31:0] wdataCounter_io_out; // @[AXIProtocol.scala 59:28:@46446.4]
  wire [31:0] wdataCounter_io_next; // @[AXIProtocol.scala 59:28:@46446.4]
  reg  writeIssued; // @[AXIProtocol.scala 61:28:@46449.4]
  reg [31:0] _RAND_0;
  wire  dramCmdIssue; // @[AXIProtocol.scala 63:39:@46450.4]
  wire  dramWriteIssue; // @[AXIProtocol.scala 64:43:@46451.4]
  wire  _T_201; // @[AXIProtocol.scala 68:54:@46452.4]
  wire  wlast; // @[AXIProtocol.scala 68:30:@46453.4]
  wire  _T_203; // @[AXIProtocol.scala 72:28:@46459.6]
  wire  _GEN_0; // @[AXIProtocol.scala 72:40:@46460.6]
  wire  _GEN_1; // @[AXIProtocol.scala 70:15:@46455.4]
  wire  _T_208; // @[AXIProtocol.scala 84:55:@46469.4]
  wire  _T_210; // @[AXIProtocol.scala 84:44:@46470.4]
  Counter_72 wdataCounter ( // @[AXIProtocol.scala 59:28:@46446.4]
    .clock(wdataCounter_clock),
    .reset(wdataCounter_reset),
    .io_reset(wdataCounter_io_reset),
    .io_enable(wdataCounter_io_enable),
    .io_stride(wdataCounter_io_stride),
    .io_out(wdataCounter_io_out),
    .io_next(wdataCounter_io_next)
  );
  assign dramCmdIssue = io_out_cmd_valid & io_out_cmd_ready; // @[AXIProtocol.scala 63:39:@46450.4]
  assign dramWriteIssue = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 64:43:@46451.4]
  assign _T_201 = wdataCounter_io_next == io_in_cmd_bits_size; // @[AXIProtocol.scala 68:54:@46452.4]
  assign wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 68:30:@46453.4]
  assign _T_203 = dramCmdIssue & io_in_cmd_bits_isWr; // @[AXIProtocol.scala 72:28:@46459.6]
  assign _GEN_0 = _T_203 ? 1'h1 : writeIssued; // @[AXIProtocol.scala 72:40:@46460.6]
  assign _GEN_1 = wlast ? 1'h0 : _GEN_0; // @[AXIProtocol.scala 70:15:@46455.4]
  assign _T_208 = writeIssued == 1'h0; // @[AXIProtocol.scala 84:55:@46469.4]
  assign _T_210 = io_in_cmd_bits_isWr ? _T_208 : 1'h1; // @[AXIProtocol.scala 84:44:@46470.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? wlast : dramCmdIssue; // @[AXIProtocol.scala 56:10:@46445.4 AXIProtocol.scala 81:19:@46467.4]
  assign io_in_wdata_ready = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 56:10:@46438.4 AXIProtocol.scala 82:21:@46468.4]
  assign io_in_wresp_valid = io_out_wresp_valid; // @[AXIProtocol.scala 56:10:@46335.4]
  assign io_in_wresp_bits_tag = io_out_wresp_bits_tag; // @[AXIProtocol.scala 56:10:@46334.4]
  assign io_out_cmd_valid = io_in_cmd_valid & _T_210; // @[AXIProtocol.scala 56:10:@46444.4 AXIProtocol.scala 84:20:@46472.4]
  assign io_out_cmd_bits_addr = io_in_cmd_bits_addr; // @[AXIProtocol.scala 56:10:@46443.4]
  assign io_out_cmd_bits_size = io_in_cmd_bits_size; // @[AXIProtocol.scala 56:10:@46442.4]
  assign io_out_cmd_bits_isWr = io_in_cmd_bits_isWr; // @[AXIProtocol.scala 56:10:@46440.4]
  assign io_out_cmd_bits_tag = io_in_cmd_bits_tag; // @[AXIProtocol.scala 56:10:@46439.4]
  assign io_out_wdata_valid = io_in_wdata_valid & writeIssued; // @[AXIProtocol.scala 56:10:@46437.4 AXIProtocol.scala 86:22:@46474.4]
  assign io_out_wdata_bits_wdata_0 = io_in_wdata_bits_wdata_0; // @[AXIProtocol.scala 56:10:@46421.4]
  assign io_out_wdata_bits_wdata_1 = io_in_wdata_bits_wdata_1; // @[AXIProtocol.scala 56:10:@46422.4]
  assign io_out_wdata_bits_wdata_2 = io_in_wdata_bits_wdata_2; // @[AXIProtocol.scala 56:10:@46423.4]
  assign io_out_wdata_bits_wdata_3 = io_in_wdata_bits_wdata_3; // @[AXIProtocol.scala 56:10:@46424.4]
  assign io_out_wdata_bits_wdata_4 = io_in_wdata_bits_wdata_4; // @[AXIProtocol.scala 56:10:@46425.4]
  assign io_out_wdata_bits_wdata_5 = io_in_wdata_bits_wdata_5; // @[AXIProtocol.scala 56:10:@46426.4]
  assign io_out_wdata_bits_wdata_6 = io_in_wdata_bits_wdata_6; // @[AXIProtocol.scala 56:10:@46427.4]
  assign io_out_wdata_bits_wdata_7 = io_in_wdata_bits_wdata_7; // @[AXIProtocol.scala 56:10:@46428.4]
  assign io_out_wdata_bits_wdata_8 = io_in_wdata_bits_wdata_8; // @[AXIProtocol.scala 56:10:@46429.4]
  assign io_out_wdata_bits_wdata_9 = io_in_wdata_bits_wdata_9; // @[AXIProtocol.scala 56:10:@46430.4]
  assign io_out_wdata_bits_wdata_10 = io_in_wdata_bits_wdata_10; // @[AXIProtocol.scala 56:10:@46431.4]
  assign io_out_wdata_bits_wdata_11 = io_in_wdata_bits_wdata_11; // @[AXIProtocol.scala 56:10:@46432.4]
  assign io_out_wdata_bits_wdata_12 = io_in_wdata_bits_wdata_12; // @[AXIProtocol.scala 56:10:@46433.4]
  assign io_out_wdata_bits_wdata_13 = io_in_wdata_bits_wdata_13; // @[AXIProtocol.scala 56:10:@46434.4]
  assign io_out_wdata_bits_wdata_14 = io_in_wdata_bits_wdata_14; // @[AXIProtocol.scala 56:10:@46435.4]
  assign io_out_wdata_bits_wdata_15 = io_in_wdata_bits_wdata_15; // @[AXIProtocol.scala 56:10:@46436.4]
  assign io_out_wdata_bits_wstrb_0 = io_in_wdata_bits_wstrb_0; // @[AXIProtocol.scala 56:10:@46357.4]
  assign io_out_wdata_bits_wstrb_1 = io_in_wdata_bits_wstrb_1; // @[AXIProtocol.scala 56:10:@46358.4]
  assign io_out_wdata_bits_wstrb_2 = io_in_wdata_bits_wstrb_2; // @[AXIProtocol.scala 56:10:@46359.4]
  assign io_out_wdata_bits_wstrb_3 = io_in_wdata_bits_wstrb_3; // @[AXIProtocol.scala 56:10:@46360.4]
  assign io_out_wdata_bits_wstrb_4 = io_in_wdata_bits_wstrb_4; // @[AXIProtocol.scala 56:10:@46361.4]
  assign io_out_wdata_bits_wstrb_5 = io_in_wdata_bits_wstrb_5; // @[AXIProtocol.scala 56:10:@46362.4]
  assign io_out_wdata_bits_wstrb_6 = io_in_wdata_bits_wstrb_6; // @[AXIProtocol.scala 56:10:@46363.4]
  assign io_out_wdata_bits_wstrb_7 = io_in_wdata_bits_wstrb_7; // @[AXIProtocol.scala 56:10:@46364.4]
  assign io_out_wdata_bits_wstrb_8 = io_in_wdata_bits_wstrb_8; // @[AXIProtocol.scala 56:10:@46365.4]
  assign io_out_wdata_bits_wstrb_9 = io_in_wdata_bits_wstrb_9; // @[AXIProtocol.scala 56:10:@46366.4]
  assign io_out_wdata_bits_wstrb_10 = io_in_wdata_bits_wstrb_10; // @[AXIProtocol.scala 56:10:@46367.4]
  assign io_out_wdata_bits_wstrb_11 = io_in_wdata_bits_wstrb_11; // @[AXIProtocol.scala 56:10:@46368.4]
  assign io_out_wdata_bits_wstrb_12 = io_in_wdata_bits_wstrb_12; // @[AXIProtocol.scala 56:10:@46369.4]
  assign io_out_wdata_bits_wstrb_13 = io_in_wdata_bits_wstrb_13; // @[AXIProtocol.scala 56:10:@46370.4]
  assign io_out_wdata_bits_wstrb_14 = io_in_wdata_bits_wstrb_14; // @[AXIProtocol.scala 56:10:@46371.4]
  assign io_out_wdata_bits_wstrb_15 = io_in_wdata_bits_wstrb_15; // @[AXIProtocol.scala 56:10:@46372.4]
  assign io_out_wdata_bits_wstrb_16 = io_in_wdata_bits_wstrb_16; // @[AXIProtocol.scala 56:10:@46373.4]
  assign io_out_wdata_bits_wstrb_17 = io_in_wdata_bits_wstrb_17; // @[AXIProtocol.scala 56:10:@46374.4]
  assign io_out_wdata_bits_wstrb_18 = io_in_wdata_bits_wstrb_18; // @[AXIProtocol.scala 56:10:@46375.4]
  assign io_out_wdata_bits_wstrb_19 = io_in_wdata_bits_wstrb_19; // @[AXIProtocol.scala 56:10:@46376.4]
  assign io_out_wdata_bits_wstrb_20 = io_in_wdata_bits_wstrb_20; // @[AXIProtocol.scala 56:10:@46377.4]
  assign io_out_wdata_bits_wstrb_21 = io_in_wdata_bits_wstrb_21; // @[AXIProtocol.scala 56:10:@46378.4]
  assign io_out_wdata_bits_wstrb_22 = io_in_wdata_bits_wstrb_22; // @[AXIProtocol.scala 56:10:@46379.4]
  assign io_out_wdata_bits_wstrb_23 = io_in_wdata_bits_wstrb_23; // @[AXIProtocol.scala 56:10:@46380.4]
  assign io_out_wdata_bits_wstrb_24 = io_in_wdata_bits_wstrb_24; // @[AXIProtocol.scala 56:10:@46381.4]
  assign io_out_wdata_bits_wstrb_25 = io_in_wdata_bits_wstrb_25; // @[AXIProtocol.scala 56:10:@46382.4]
  assign io_out_wdata_bits_wstrb_26 = io_in_wdata_bits_wstrb_26; // @[AXIProtocol.scala 56:10:@46383.4]
  assign io_out_wdata_bits_wstrb_27 = io_in_wdata_bits_wstrb_27; // @[AXIProtocol.scala 56:10:@46384.4]
  assign io_out_wdata_bits_wstrb_28 = io_in_wdata_bits_wstrb_28; // @[AXIProtocol.scala 56:10:@46385.4]
  assign io_out_wdata_bits_wstrb_29 = io_in_wdata_bits_wstrb_29; // @[AXIProtocol.scala 56:10:@46386.4]
  assign io_out_wdata_bits_wstrb_30 = io_in_wdata_bits_wstrb_30; // @[AXIProtocol.scala 56:10:@46387.4]
  assign io_out_wdata_bits_wstrb_31 = io_in_wdata_bits_wstrb_31; // @[AXIProtocol.scala 56:10:@46388.4]
  assign io_out_wdata_bits_wstrb_32 = io_in_wdata_bits_wstrb_32; // @[AXIProtocol.scala 56:10:@46389.4]
  assign io_out_wdata_bits_wstrb_33 = io_in_wdata_bits_wstrb_33; // @[AXIProtocol.scala 56:10:@46390.4]
  assign io_out_wdata_bits_wstrb_34 = io_in_wdata_bits_wstrb_34; // @[AXIProtocol.scala 56:10:@46391.4]
  assign io_out_wdata_bits_wstrb_35 = io_in_wdata_bits_wstrb_35; // @[AXIProtocol.scala 56:10:@46392.4]
  assign io_out_wdata_bits_wstrb_36 = io_in_wdata_bits_wstrb_36; // @[AXIProtocol.scala 56:10:@46393.4]
  assign io_out_wdata_bits_wstrb_37 = io_in_wdata_bits_wstrb_37; // @[AXIProtocol.scala 56:10:@46394.4]
  assign io_out_wdata_bits_wstrb_38 = io_in_wdata_bits_wstrb_38; // @[AXIProtocol.scala 56:10:@46395.4]
  assign io_out_wdata_bits_wstrb_39 = io_in_wdata_bits_wstrb_39; // @[AXIProtocol.scala 56:10:@46396.4]
  assign io_out_wdata_bits_wstrb_40 = io_in_wdata_bits_wstrb_40; // @[AXIProtocol.scala 56:10:@46397.4]
  assign io_out_wdata_bits_wstrb_41 = io_in_wdata_bits_wstrb_41; // @[AXIProtocol.scala 56:10:@46398.4]
  assign io_out_wdata_bits_wstrb_42 = io_in_wdata_bits_wstrb_42; // @[AXIProtocol.scala 56:10:@46399.4]
  assign io_out_wdata_bits_wstrb_43 = io_in_wdata_bits_wstrb_43; // @[AXIProtocol.scala 56:10:@46400.4]
  assign io_out_wdata_bits_wstrb_44 = io_in_wdata_bits_wstrb_44; // @[AXIProtocol.scala 56:10:@46401.4]
  assign io_out_wdata_bits_wstrb_45 = io_in_wdata_bits_wstrb_45; // @[AXIProtocol.scala 56:10:@46402.4]
  assign io_out_wdata_bits_wstrb_46 = io_in_wdata_bits_wstrb_46; // @[AXIProtocol.scala 56:10:@46403.4]
  assign io_out_wdata_bits_wstrb_47 = io_in_wdata_bits_wstrb_47; // @[AXIProtocol.scala 56:10:@46404.4]
  assign io_out_wdata_bits_wstrb_48 = io_in_wdata_bits_wstrb_48; // @[AXIProtocol.scala 56:10:@46405.4]
  assign io_out_wdata_bits_wstrb_49 = io_in_wdata_bits_wstrb_49; // @[AXIProtocol.scala 56:10:@46406.4]
  assign io_out_wdata_bits_wstrb_50 = io_in_wdata_bits_wstrb_50; // @[AXIProtocol.scala 56:10:@46407.4]
  assign io_out_wdata_bits_wstrb_51 = io_in_wdata_bits_wstrb_51; // @[AXIProtocol.scala 56:10:@46408.4]
  assign io_out_wdata_bits_wstrb_52 = io_in_wdata_bits_wstrb_52; // @[AXIProtocol.scala 56:10:@46409.4]
  assign io_out_wdata_bits_wstrb_53 = io_in_wdata_bits_wstrb_53; // @[AXIProtocol.scala 56:10:@46410.4]
  assign io_out_wdata_bits_wstrb_54 = io_in_wdata_bits_wstrb_54; // @[AXIProtocol.scala 56:10:@46411.4]
  assign io_out_wdata_bits_wstrb_55 = io_in_wdata_bits_wstrb_55; // @[AXIProtocol.scala 56:10:@46412.4]
  assign io_out_wdata_bits_wstrb_56 = io_in_wdata_bits_wstrb_56; // @[AXIProtocol.scala 56:10:@46413.4]
  assign io_out_wdata_bits_wstrb_57 = io_in_wdata_bits_wstrb_57; // @[AXIProtocol.scala 56:10:@46414.4]
  assign io_out_wdata_bits_wstrb_58 = io_in_wdata_bits_wstrb_58; // @[AXIProtocol.scala 56:10:@46415.4]
  assign io_out_wdata_bits_wstrb_59 = io_in_wdata_bits_wstrb_59; // @[AXIProtocol.scala 56:10:@46416.4]
  assign io_out_wdata_bits_wstrb_60 = io_in_wdata_bits_wstrb_60; // @[AXIProtocol.scala 56:10:@46417.4]
  assign io_out_wdata_bits_wstrb_61 = io_in_wdata_bits_wstrb_61; // @[AXIProtocol.scala 56:10:@46418.4]
  assign io_out_wdata_bits_wstrb_62 = io_in_wdata_bits_wstrb_62; // @[AXIProtocol.scala 56:10:@46419.4]
  assign io_out_wdata_bits_wstrb_63 = io_in_wdata_bits_wstrb_63; // @[AXIProtocol.scala 56:10:@46420.4]
  assign io_out_wdata_bits_wlast = dramWriteIssue & _T_201; // @[AXIProtocol.scala 56:10:@46356.4 AXIProtocol.scala 87:27:@46475.4]
  assign io_out_rresp_ready = io_in_rresp_ready; // @[AXIProtocol.scala 56:10:@46355.4]
  assign io_out_wresp_ready = io_in_wresp_ready; // @[AXIProtocol.scala 56:10:@46336.4]
  assign wdataCounter_clock = clock; // @[:@46447.4]
  assign wdataCounter_reset = reset; // @[:@46448.4]
  assign wdataCounter_io_reset = dramWriteIssue & _T_201; // @[AXIProtocol.scala 76:25:@46463.4]
  assign wdataCounter_io_enable = io_out_wdata_valid & io_out_wdata_ready; // @[AXIProtocol.scala 77:26:@46464.4]
  assign wdataCounter_io_stride = 32'h1; // @[AXIProtocol.scala 78:26:@46465.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeIssued = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      writeIssued <= 1'h0;
    end else begin
      if (wlast) begin
        writeIssued <= 1'h0;
      end else begin
        if (_T_203) begin
          writeIssued <= 1'h1;
        end
      end
    end
  end
endmodule
module DRAMArbiter( // @[:@46477.2]
  input         clock, // @[:@46478.4]
  input         reset, // @[:@46479.4]
  input         io_enable, // @[:@46480.4]
  output        io_app_stores_0_cmd_ready, // @[:@46480.4]
  input         io_app_stores_0_cmd_valid, // @[:@46480.4]
  input  [63:0] io_app_stores_0_cmd_bits_addr, // @[:@46480.4]
  input  [31:0] io_app_stores_0_cmd_bits_size, // @[:@46480.4]
  output        io_app_stores_0_data_ready, // @[:@46480.4]
  input         io_app_stores_0_data_valid, // @[:@46480.4]
  input  [31:0] io_app_stores_0_data_bits_wdata_0, // @[:@46480.4]
  input         io_app_stores_0_data_bits_wstrb, // @[:@46480.4]
  input         io_app_stores_0_wresp_ready, // @[:@46480.4]
  output        io_app_stores_0_wresp_valid, // @[:@46480.4]
  output        io_app_stores_0_wresp_bits, // @[:@46480.4]
  input         io_dram_cmd_ready, // @[:@46480.4]
  output        io_dram_cmd_valid, // @[:@46480.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@46480.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@46480.4]
  output        io_dram_cmd_bits_isWr, // @[:@46480.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@46480.4]
  input         io_dram_wdata_ready, // @[:@46480.4]
  output        io_dram_wdata_valid, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@46480.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@46480.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@46480.4]
  output        io_dram_wdata_bits_wlast, // @[:@46480.4]
  output        io_dram_rresp_ready, // @[:@46480.4]
  output        io_dram_wresp_ready, // @[:@46480.4]
  input         io_dram_wresp_valid, // @[:@46480.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@46480.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@47366.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@47380.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@47608.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@47723.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@47723.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@47366.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@47380.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@47608.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@47723.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_app_stores_0_cmd_ready = StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 68:18:@47379.4]
  assign io_app_stores_0_data_ready = StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 68:18:@47375.4]
  assign io_app_stores_0_wresp_valid = StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 68:18:@47370.4]
  assign io_app_stores_0_wresp_bits = StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 68:18:@47369.4]
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@47948.4 DRAMArbiter.scala 100:23:@47951.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@47947.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@47946.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@47944.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@47943.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@47941.4 DRAMArbiter.scala 101:25:@47953.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@47925.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@47926.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@47927.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@47928.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@47929.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@47930.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@47931.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@47932.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@47933.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@47934.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@47935.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@47936.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@47937.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@47938.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@47939.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@47940.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@47861.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@47862.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@47863.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@47864.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@47865.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@47866.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@47867.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@47868.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@47869.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@47870.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@47871.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@47872.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@47873.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@47874.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@47875.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@47876.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@47877.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@47878.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@47879.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@47880.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@47881.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@47882.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@47883.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@47884.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@47885.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@47886.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@47887.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@47888.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@47889.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@47890.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@47891.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@47892.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@47893.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@47894.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@47895.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@47896.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@47897.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@47898.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@47899.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@47900.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@47901.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@47902.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@47903.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@47904.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@47905.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@47906.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@47907.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@47908.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@47909.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@47910.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@47911.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@47912.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@47913.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@47914.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@47915.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@47916.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@47917.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@47918.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@47919.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@47920.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@47921.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@47922.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@47923.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@47924.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@47860.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@47859.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@47840.4]
  assign StreamControllerStore_clock = clock; // @[:@47367.4]
  assign StreamControllerStore_reset = reset; // @[:@47368.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@47495.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@47488.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@47385.4]
  assign StreamControllerStore_io_store_cmd_valid = io_app_stores_0_cmd_valid; // @[DRAMArbiter.scala 68:18:@47378.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = io_app_stores_0_cmd_bits_addr; // @[DRAMArbiter.scala 68:18:@47377.4]
  assign StreamControllerStore_io_store_cmd_bits_size = io_app_stores_0_cmd_bits_size; // @[DRAMArbiter.scala 68:18:@47376.4]
  assign StreamControllerStore_io_store_data_valid = io_app_stores_0_data_valid; // @[DRAMArbiter.scala 68:18:@47374.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = io_app_stores_0_data_bits_wdata_0; // @[DRAMArbiter.scala 68:18:@47373.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = io_app_stores_0_data_bits_wstrb; // @[DRAMArbiter.scala 68:18:@47372.4]
  assign StreamControllerStore_io_store_wresp_ready = io_app_stores_0_wresp_ready; // @[DRAMArbiter.scala 68:18:@47371.4]
  assign StreamArbiter_clock = clock; // @[:@47381.4]
  assign StreamArbiter_reset = reset; // @[:@47382.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@47606.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@47605.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@47604.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@47602.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@47601.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@47599.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@47583.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@47584.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@47585.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@47586.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@47587.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@47588.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@47589.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@47590.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@47591.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@47592.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@47593.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@47594.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@47595.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@47596.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@47597.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@47598.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@47519.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@47520.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@47521.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@47522.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@47523.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@47524.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@47525.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@47526.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@47527.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@47528.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@47529.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@47530.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@47531.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@47532.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@47533.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@47534.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@47535.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@47536.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@47537.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@47538.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@47539.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@47540.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@47541.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@47542.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@47543.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@47544.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@47545.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@47546.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@47547.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@47548.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@47549.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@47550.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@47551.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@47552.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@47553.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@47554.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@47555.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@47556.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@47557.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@47558.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@47559.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@47560.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@47561.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@47562.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@47563.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@47564.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@47565.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@47566.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@47567.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@47568.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@47569.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@47570.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@47571.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@47572.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@47573.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@47574.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@47575.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@47576.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@47577.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@47578.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@47579.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@47580.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@47581.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@47582.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@47517.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@47498.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@47722.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@47715.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@47612.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@47611.4]
  assign AXICmdSplit_clock = clock; // @[:@47609.4]
  assign AXICmdSplit_reset = reset; // @[:@47610.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@47721.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@47720.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@47719.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@47717.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@47716.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@47714.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@47698.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@47699.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@47700.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@47701.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@47702.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@47703.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@47704.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@47705.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@47706.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@47707.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@47708.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@47709.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@47710.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@47711.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@47712.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@47713.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@47634.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@47635.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@47636.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@47637.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@47638.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@47639.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@47640.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@47641.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@47642.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@47643.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@47644.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@47645.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@47646.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@47647.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@47648.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@47649.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@47650.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@47651.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@47652.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@47653.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@47654.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@47655.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@47656.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@47657.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@47658.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@47659.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@47660.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@47661.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@47662.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@47663.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@47664.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@47665.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@47666.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@47667.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@47668.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@47669.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@47670.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@47671.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@47672.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@47673.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@47674.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@47675.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@47676.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@47677.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@47678.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@47679.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@47680.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@47681.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@47682.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@47683.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@47684.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@47685.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@47686.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@47687.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@47688.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@47689.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@47690.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@47691.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@47692.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@47693.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@47694.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@47695.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@47696.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@47697.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@47632.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@47613.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@47837.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@47830.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@47727.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@47726.4]
  assign AXICmdIssue_clock = clock; // @[:@47724.4]
  assign AXICmdIssue_reset = reset; // @[:@47725.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@47836.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@47835.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@47834.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@47832.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@47831.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@47829.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@47813.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@47814.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@47815.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@47816.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@47817.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@47818.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@47819.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@47820.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@47821.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@47822.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@47823.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@47824.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@47825.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@47826.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@47827.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@47828.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@47749.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@47750.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@47751.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@47752.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@47753.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@47754.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@47755.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@47756.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@47757.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@47758.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@47759.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@47760.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@47761.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@47762.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@47763.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@47764.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@47765.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@47766.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@47767.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@47768.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@47769.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@47770.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@47771.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@47772.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@47773.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@47774.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@47775.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@47776.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@47777.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@47778.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@47779.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@47780.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@47781.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@47782.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@47783.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@47784.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@47785.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@47786.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@47787.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@47788.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@47789.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@47790.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@47791.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@47792.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@47793.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@47794.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@47795.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@47796.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@47797.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@47798.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@47799.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@47800.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@47801.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@47802.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@47803.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@47804.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@47805.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@47806.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@47807.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@47808.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@47809.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@47810.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@47811.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@47812.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@47747.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@47728.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@47949.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@47942.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@47839.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@47838.4]
endmodule
module DRAMArbiter_1( // @[:@62178.2]
  input         clock, // @[:@62179.4]
  input         reset, // @[:@62180.4]
  input         io_enable, // @[:@62181.4]
  input         io_dram_cmd_ready, // @[:@62181.4]
  output        io_dram_cmd_valid, // @[:@62181.4]
  output [63:0] io_dram_cmd_bits_addr, // @[:@62181.4]
  output [31:0] io_dram_cmd_bits_size, // @[:@62181.4]
  output        io_dram_cmd_bits_isWr, // @[:@62181.4]
  output [31:0] io_dram_cmd_bits_tag, // @[:@62181.4]
  input         io_dram_wdata_ready, // @[:@62181.4]
  output        io_dram_wdata_valid, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_0, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_1, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_2, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_3, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_4, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_5, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_6, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_7, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_8, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_9, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_10, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_11, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_12, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_13, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_14, // @[:@62181.4]
  output [31:0] io_dram_wdata_bits_wdata_15, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_0, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_1, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_2, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_3, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_4, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_5, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_6, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_7, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_8, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_9, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_10, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_11, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_12, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_13, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_14, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_15, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_16, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_17, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_18, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_19, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_20, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_21, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_22, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_23, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_24, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_25, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_26, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_27, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_28, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_29, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_30, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_31, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_32, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_33, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_34, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_35, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_36, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_37, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_38, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_39, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_40, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_41, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_42, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_43, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_44, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_45, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_46, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_47, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_48, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_49, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_50, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_51, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_52, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_53, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_54, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_55, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_56, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_57, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_58, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_59, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_60, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_61, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_62, // @[:@62181.4]
  output        io_dram_wdata_bits_wstrb_63, // @[:@62181.4]
  output        io_dram_wdata_bits_wlast, // @[:@62181.4]
  output        io_dram_rresp_ready, // @[:@62181.4]
  output        io_dram_wresp_ready, // @[:@62181.4]
  input         io_dram_wresp_valid, // @[:@62181.4]
  input  [31:0] io_dram_wresp_bits_tag // @[:@62181.4]
);
  wire  StreamControllerStore_clock; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_reset; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_cmd_ready; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [63:0] StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_ready; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_dram_wresp_valid; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_store_cmd_ready; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_store_cmd_valid; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [63:0] StreamControllerStore_io_store_cmd_bits_addr; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_store_cmd_bits_size; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_store_data_ready; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_store_data_valid; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire [31:0] StreamControllerStore_io_store_data_bits_wdata_0; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_store_data_bits_wstrb; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_store_wresp_ready; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_store_wresp_valid; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamControllerStore_io_store_wresp_bits; // @[DRAMArbiter.scala 67:21:@63067.4]
  wire  StreamArbiter_clock; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_reset; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_cmd_valid; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [63:0] StreamArbiter_io_app_0_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_valid; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_app_0_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_rresp_ready; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wresp_ready; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_cmd_ready; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [63:0] StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_ready; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  StreamArbiter_io_dram_wresp_valid; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire [31:0] StreamArbiter_io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 86:27:@63081.4]
  wire  AXICmdSplit_clock; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_reset; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_cmd_valid; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [63:0] AXICmdSplit_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_valid; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_rresp_ready; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wresp_ready; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_cmd_ready; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [63:0] AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_ready; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdSplit_io_out_wresp_valid; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire [31:0] AXICmdSplit_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 94:26:@63309.4]
  wire  AXICmdIssue_clock; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_reset; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_cmd_valid; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [63:0] AXICmdIssue_io_in_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_valid; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_rresp_ready; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wresp_ready; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_cmd_ready; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [63:0] AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_ready; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire  AXICmdIssue_io_out_wresp_valid; // @[DRAMArbiter.scala 97:26:@63424.4]
  wire [31:0] AXICmdIssue_io_out_wresp_bits_tag; // @[DRAMArbiter.scala 97:26:@63424.4]
  StreamControllerStore StreamControllerStore ( // @[DRAMArbiter.scala 67:21:@63067.4]
    .clock(StreamControllerStore_clock),
    .reset(StreamControllerStore_reset),
    .io_dram_cmd_ready(StreamControllerStore_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamControllerStore_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamControllerStore_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamControllerStore_io_dram_cmd_bits_size),
    .io_dram_wdata_ready(StreamControllerStore_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamControllerStore_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamControllerStore_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamControllerStore_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamControllerStore_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamControllerStore_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamControllerStore_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamControllerStore_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamControllerStore_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamControllerStore_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamControllerStore_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamControllerStore_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamControllerStore_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamControllerStore_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamControllerStore_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamControllerStore_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamControllerStore_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamControllerStore_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamControllerStore_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamControllerStore_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamControllerStore_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamControllerStore_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamControllerStore_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamControllerStore_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamControllerStore_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamControllerStore_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamControllerStore_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamControllerStore_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamControllerStore_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamControllerStore_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamControllerStore_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamControllerStore_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamControllerStore_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamControllerStore_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamControllerStore_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamControllerStore_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamControllerStore_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamControllerStore_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamControllerStore_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamControllerStore_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamControllerStore_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamControllerStore_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamControllerStore_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamControllerStore_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamControllerStore_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamControllerStore_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamControllerStore_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamControllerStore_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamControllerStore_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamControllerStore_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamControllerStore_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamControllerStore_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamControllerStore_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamControllerStore_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamControllerStore_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamControllerStore_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamControllerStore_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamControllerStore_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamControllerStore_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamControllerStore_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamControllerStore_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamControllerStore_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamControllerStore_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamControllerStore_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamControllerStore_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamControllerStore_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamControllerStore_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamControllerStore_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamControllerStore_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamControllerStore_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamControllerStore_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamControllerStore_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamControllerStore_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamControllerStore_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamControllerStore_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamControllerStore_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamControllerStore_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamControllerStore_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamControllerStore_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamControllerStore_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamControllerStore_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamControllerStore_io_dram_wdata_bits_wstrb_63),
    .io_dram_wresp_ready(StreamControllerStore_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamControllerStore_io_dram_wresp_valid),
    .io_store_cmd_ready(StreamControllerStore_io_store_cmd_ready),
    .io_store_cmd_valid(StreamControllerStore_io_store_cmd_valid),
    .io_store_cmd_bits_addr(StreamControllerStore_io_store_cmd_bits_addr),
    .io_store_cmd_bits_size(StreamControllerStore_io_store_cmd_bits_size),
    .io_store_data_ready(StreamControllerStore_io_store_data_ready),
    .io_store_data_valid(StreamControllerStore_io_store_data_valid),
    .io_store_data_bits_wdata_0(StreamControllerStore_io_store_data_bits_wdata_0),
    .io_store_data_bits_wstrb(StreamControllerStore_io_store_data_bits_wstrb),
    .io_store_wresp_ready(StreamControllerStore_io_store_wresp_ready),
    .io_store_wresp_valid(StreamControllerStore_io_store_wresp_valid),
    .io_store_wresp_bits(StreamControllerStore_io_store_wresp_bits)
  );
  StreamArbiter StreamArbiter ( // @[DRAMArbiter.scala 86:27:@63081.4]
    .clock(StreamArbiter_clock),
    .reset(StreamArbiter_reset),
    .io_app_0_cmd_ready(StreamArbiter_io_app_0_cmd_ready),
    .io_app_0_cmd_valid(StreamArbiter_io_app_0_cmd_valid),
    .io_app_0_cmd_bits_addr(StreamArbiter_io_app_0_cmd_bits_addr),
    .io_app_0_cmd_bits_size(StreamArbiter_io_app_0_cmd_bits_size),
    .io_app_0_cmd_bits_isWr(StreamArbiter_io_app_0_cmd_bits_isWr),
    .io_app_0_cmd_bits_tag(StreamArbiter_io_app_0_cmd_bits_tag),
    .io_app_0_wdata_ready(StreamArbiter_io_app_0_wdata_ready),
    .io_app_0_wdata_valid(StreamArbiter_io_app_0_wdata_valid),
    .io_app_0_wdata_bits_wdata_0(StreamArbiter_io_app_0_wdata_bits_wdata_0),
    .io_app_0_wdata_bits_wdata_1(StreamArbiter_io_app_0_wdata_bits_wdata_1),
    .io_app_0_wdata_bits_wdata_2(StreamArbiter_io_app_0_wdata_bits_wdata_2),
    .io_app_0_wdata_bits_wdata_3(StreamArbiter_io_app_0_wdata_bits_wdata_3),
    .io_app_0_wdata_bits_wdata_4(StreamArbiter_io_app_0_wdata_bits_wdata_4),
    .io_app_0_wdata_bits_wdata_5(StreamArbiter_io_app_0_wdata_bits_wdata_5),
    .io_app_0_wdata_bits_wdata_6(StreamArbiter_io_app_0_wdata_bits_wdata_6),
    .io_app_0_wdata_bits_wdata_7(StreamArbiter_io_app_0_wdata_bits_wdata_7),
    .io_app_0_wdata_bits_wdata_8(StreamArbiter_io_app_0_wdata_bits_wdata_8),
    .io_app_0_wdata_bits_wdata_9(StreamArbiter_io_app_0_wdata_bits_wdata_9),
    .io_app_0_wdata_bits_wdata_10(StreamArbiter_io_app_0_wdata_bits_wdata_10),
    .io_app_0_wdata_bits_wdata_11(StreamArbiter_io_app_0_wdata_bits_wdata_11),
    .io_app_0_wdata_bits_wdata_12(StreamArbiter_io_app_0_wdata_bits_wdata_12),
    .io_app_0_wdata_bits_wdata_13(StreamArbiter_io_app_0_wdata_bits_wdata_13),
    .io_app_0_wdata_bits_wdata_14(StreamArbiter_io_app_0_wdata_bits_wdata_14),
    .io_app_0_wdata_bits_wdata_15(StreamArbiter_io_app_0_wdata_bits_wdata_15),
    .io_app_0_wdata_bits_wstrb_0(StreamArbiter_io_app_0_wdata_bits_wstrb_0),
    .io_app_0_wdata_bits_wstrb_1(StreamArbiter_io_app_0_wdata_bits_wstrb_1),
    .io_app_0_wdata_bits_wstrb_2(StreamArbiter_io_app_0_wdata_bits_wstrb_2),
    .io_app_0_wdata_bits_wstrb_3(StreamArbiter_io_app_0_wdata_bits_wstrb_3),
    .io_app_0_wdata_bits_wstrb_4(StreamArbiter_io_app_0_wdata_bits_wstrb_4),
    .io_app_0_wdata_bits_wstrb_5(StreamArbiter_io_app_0_wdata_bits_wstrb_5),
    .io_app_0_wdata_bits_wstrb_6(StreamArbiter_io_app_0_wdata_bits_wstrb_6),
    .io_app_0_wdata_bits_wstrb_7(StreamArbiter_io_app_0_wdata_bits_wstrb_7),
    .io_app_0_wdata_bits_wstrb_8(StreamArbiter_io_app_0_wdata_bits_wstrb_8),
    .io_app_0_wdata_bits_wstrb_9(StreamArbiter_io_app_0_wdata_bits_wstrb_9),
    .io_app_0_wdata_bits_wstrb_10(StreamArbiter_io_app_0_wdata_bits_wstrb_10),
    .io_app_0_wdata_bits_wstrb_11(StreamArbiter_io_app_0_wdata_bits_wstrb_11),
    .io_app_0_wdata_bits_wstrb_12(StreamArbiter_io_app_0_wdata_bits_wstrb_12),
    .io_app_0_wdata_bits_wstrb_13(StreamArbiter_io_app_0_wdata_bits_wstrb_13),
    .io_app_0_wdata_bits_wstrb_14(StreamArbiter_io_app_0_wdata_bits_wstrb_14),
    .io_app_0_wdata_bits_wstrb_15(StreamArbiter_io_app_0_wdata_bits_wstrb_15),
    .io_app_0_wdata_bits_wstrb_16(StreamArbiter_io_app_0_wdata_bits_wstrb_16),
    .io_app_0_wdata_bits_wstrb_17(StreamArbiter_io_app_0_wdata_bits_wstrb_17),
    .io_app_0_wdata_bits_wstrb_18(StreamArbiter_io_app_0_wdata_bits_wstrb_18),
    .io_app_0_wdata_bits_wstrb_19(StreamArbiter_io_app_0_wdata_bits_wstrb_19),
    .io_app_0_wdata_bits_wstrb_20(StreamArbiter_io_app_0_wdata_bits_wstrb_20),
    .io_app_0_wdata_bits_wstrb_21(StreamArbiter_io_app_0_wdata_bits_wstrb_21),
    .io_app_0_wdata_bits_wstrb_22(StreamArbiter_io_app_0_wdata_bits_wstrb_22),
    .io_app_0_wdata_bits_wstrb_23(StreamArbiter_io_app_0_wdata_bits_wstrb_23),
    .io_app_0_wdata_bits_wstrb_24(StreamArbiter_io_app_0_wdata_bits_wstrb_24),
    .io_app_0_wdata_bits_wstrb_25(StreamArbiter_io_app_0_wdata_bits_wstrb_25),
    .io_app_0_wdata_bits_wstrb_26(StreamArbiter_io_app_0_wdata_bits_wstrb_26),
    .io_app_0_wdata_bits_wstrb_27(StreamArbiter_io_app_0_wdata_bits_wstrb_27),
    .io_app_0_wdata_bits_wstrb_28(StreamArbiter_io_app_0_wdata_bits_wstrb_28),
    .io_app_0_wdata_bits_wstrb_29(StreamArbiter_io_app_0_wdata_bits_wstrb_29),
    .io_app_0_wdata_bits_wstrb_30(StreamArbiter_io_app_0_wdata_bits_wstrb_30),
    .io_app_0_wdata_bits_wstrb_31(StreamArbiter_io_app_0_wdata_bits_wstrb_31),
    .io_app_0_wdata_bits_wstrb_32(StreamArbiter_io_app_0_wdata_bits_wstrb_32),
    .io_app_0_wdata_bits_wstrb_33(StreamArbiter_io_app_0_wdata_bits_wstrb_33),
    .io_app_0_wdata_bits_wstrb_34(StreamArbiter_io_app_0_wdata_bits_wstrb_34),
    .io_app_0_wdata_bits_wstrb_35(StreamArbiter_io_app_0_wdata_bits_wstrb_35),
    .io_app_0_wdata_bits_wstrb_36(StreamArbiter_io_app_0_wdata_bits_wstrb_36),
    .io_app_0_wdata_bits_wstrb_37(StreamArbiter_io_app_0_wdata_bits_wstrb_37),
    .io_app_0_wdata_bits_wstrb_38(StreamArbiter_io_app_0_wdata_bits_wstrb_38),
    .io_app_0_wdata_bits_wstrb_39(StreamArbiter_io_app_0_wdata_bits_wstrb_39),
    .io_app_0_wdata_bits_wstrb_40(StreamArbiter_io_app_0_wdata_bits_wstrb_40),
    .io_app_0_wdata_bits_wstrb_41(StreamArbiter_io_app_0_wdata_bits_wstrb_41),
    .io_app_0_wdata_bits_wstrb_42(StreamArbiter_io_app_0_wdata_bits_wstrb_42),
    .io_app_0_wdata_bits_wstrb_43(StreamArbiter_io_app_0_wdata_bits_wstrb_43),
    .io_app_0_wdata_bits_wstrb_44(StreamArbiter_io_app_0_wdata_bits_wstrb_44),
    .io_app_0_wdata_bits_wstrb_45(StreamArbiter_io_app_0_wdata_bits_wstrb_45),
    .io_app_0_wdata_bits_wstrb_46(StreamArbiter_io_app_0_wdata_bits_wstrb_46),
    .io_app_0_wdata_bits_wstrb_47(StreamArbiter_io_app_0_wdata_bits_wstrb_47),
    .io_app_0_wdata_bits_wstrb_48(StreamArbiter_io_app_0_wdata_bits_wstrb_48),
    .io_app_0_wdata_bits_wstrb_49(StreamArbiter_io_app_0_wdata_bits_wstrb_49),
    .io_app_0_wdata_bits_wstrb_50(StreamArbiter_io_app_0_wdata_bits_wstrb_50),
    .io_app_0_wdata_bits_wstrb_51(StreamArbiter_io_app_0_wdata_bits_wstrb_51),
    .io_app_0_wdata_bits_wstrb_52(StreamArbiter_io_app_0_wdata_bits_wstrb_52),
    .io_app_0_wdata_bits_wstrb_53(StreamArbiter_io_app_0_wdata_bits_wstrb_53),
    .io_app_0_wdata_bits_wstrb_54(StreamArbiter_io_app_0_wdata_bits_wstrb_54),
    .io_app_0_wdata_bits_wstrb_55(StreamArbiter_io_app_0_wdata_bits_wstrb_55),
    .io_app_0_wdata_bits_wstrb_56(StreamArbiter_io_app_0_wdata_bits_wstrb_56),
    .io_app_0_wdata_bits_wstrb_57(StreamArbiter_io_app_0_wdata_bits_wstrb_57),
    .io_app_0_wdata_bits_wstrb_58(StreamArbiter_io_app_0_wdata_bits_wstrb_58),
    .io_app_0_wdata_bits_wstrb_59(StreamArbiter_io_app_0_wdata_bits_wstrb_59),
    .io_app_0_wdata_bits_wstrb_60(StreamArbiter_io_app_0_wdata_bits_wstrb_60),
    .io_app_0_wdata_bits_wstrb_61(StreamArbiter_io_app_0_wdata_bits_wstrb_61),
    .io_app_0_wdata_bits_wstrb_62(StreamArbiter_io_app_0_wdata_bits_wstrb_62),
    .io_app_0_wdata_bits_wstrb_63(StreamArbiter_io_app_0_wdata_bits_wstrb_63),
    .io_app_0_rresp_ready(StreamArbiter_io_app_0_rresp_ready),
    .io_app_0_wresp_ready(StreamArbiter_io_app_0_wresp_ready),
    .io_app_0_wresp_valid(StreamArbiter_io_app_0_wresp_valid),
    .io_dram_cmd_ready(StreamArbiter_io_dram_cmd_ready),
    .io_dram_cmd_valid(StreamArbiter_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(StreamArbiter_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(StreamArbiter_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(StreamArbiter_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(StreamArbiter_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(StreamArbiter_io_dram_wdata_ready),
    .io_dram_wdata_valid(StreamArbiter_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(StreamArbiter_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(StreamArbiter_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(StreamArbiter_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(StreamArbiter_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(StreamArbiter_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(StreamArbiter_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(StreamArbiter_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(StreamArbiter_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(StreamArbiter_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(StreamArbiter_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(StreamArbiter_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(StreamArbiter_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(StreamArbiter_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(StreamArbiter_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(StreamArbiter_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(StreamArbiter_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(StreamArbiter_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(StreamArbiter_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(StreamArbiter_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(StreamArbiter_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(StreamArbiter_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(StreamArbiter_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(StreamArbiter_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(StreamArbiter_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(StreamArbiter_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(StreamArbiter_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(StreamArbiter_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(StreamArbiter_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(StreamArbiter_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(StreamArbiter_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(StreamArbiter_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(StreamArbiter_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(StreamArbiter_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(StreamArbiter_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(StreamArbiter_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(StreamArbiter_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(StreamArbiter_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(StreamArbiter_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(StreamArbiter_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(StreamArbiter_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(StreamArbiter_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(StreamArbiter_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(StreamArbiter_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(StreamArbiter_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(StreamArbiter_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(StreamArbiter_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(StreamArbiter_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(StreamArbiter_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(StreamArbiter_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(StreamArbiter_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(StreamArbiter_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(StreamArbiter_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(StreamArbiter_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(StreamArbiter_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(StreamArbiter_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(StreamArbiter_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(StreamArbiter_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(StreamArbiter_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(StreamArbiter_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(StreamArbiter_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(StreamArbiter_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(StreamArbiter_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(StreamArbiter_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(StreamArbiter_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(StreamArbiter_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(StreamArbiter_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(StreamArbiter_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(StreamArbiter_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(StreamArbiter_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(StreamArbiter_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(StreamArbiter_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(StreamArbiter_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(StreamArbiter_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(StreamArbiter_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(StreamArbiter_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(StreamArbiter_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(StreamArbiter_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(StreamArbiter_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(StreamArbiter_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(StreamArbiter_io_dram_wdata_bits_wstrb_63),
    .io_dram_rresp_ready(StreamArbiter_io_dram_rresp_ready),
    .io_dram_wresp_ready(StreamArbiter_io_dram_wresp_ready),
    .io_dram_wresp_valid(StreamArbiter_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(StreamArbiter_io_dram_wresp_bits_tag)
  );
  AXICmdSplit AXICmdSplit ( // @[DRAMArbiter.scala 94:26:@63309.4]
    .clock(AXICmdSplit_clock),
    .reset(AXICmdSplit_reset),
    .io_in_cmd_ready(AXICmdSplit_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdSplit_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdSplit_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdSplit_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdSplit_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdSplit_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdSplit_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdSplit_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdSplit_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdSplit_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdSplit_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdSplit_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdSplit_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdSplit_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdSplit_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdSplit_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdSplit_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdSplit_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdSplit_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdSplit_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdSplit_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdSplit_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdSplit_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdSplit_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdSplit_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdSplit_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdSplit_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdSplit_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdSplit_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdSplit_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdSplit_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdSplit_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdSplit_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdSplit_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdSplit_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdSplit_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdSplit_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdSplit_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdSplit_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdSplit_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdSplit_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdSplit_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdSplit_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdSplit_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdSplit_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdSplit_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdSplit_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdSplit_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdSplit_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdSplit_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdSplit_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdSplit_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdSplit_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdSplit_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdSplit_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdSplit_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdSplit_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdSplit_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdSplit_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdSplit_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdSplit_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdSplit_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdSplit_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdSplit_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdSplit_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdSplit_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdSplit_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdSplit_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdSplit_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdSplit_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdSplit_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdSplit_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdSplit_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdSplit_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdSplit_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdSplit_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdSplit_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdSplit_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdSplit_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdSplit_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdSplit_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdSplit_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdSplit_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdSplit_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdSplit_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdSplit_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdSplit_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdSplit_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdSplit_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdSplit_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdSplit_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdSplit_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdSplit_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdSplit_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdSplit_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdSplit_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdSplit_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdSplit_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdSplit_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdSplit_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdSplit_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdSplit_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdSplit_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdSplit_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdSplit_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdSplit_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdSplit_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdSplit_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdSplit_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdSplit_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdSplit_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdSplit_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdSplit_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdSplit_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdSplit_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdSplit_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdSplit_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdSplit_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdSplit_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdSplit_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdSplit_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdSplit_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdSplit_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdSplit_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdSplit_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdSplit_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdSplit_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdSplit_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdSplit_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdSplit_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdSplit_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdSplit_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdSplit_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdSplit_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdSplit_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdSplit_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdSplit_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdSplit_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdSplit_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdSplit_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdSplit_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdSplit_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdSplit_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdSplit_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdSplit_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdSplit_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdSplit_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdSplit_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdSplit_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdSplit_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdSplit_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdSplit_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdSplit_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdSplit_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdSplit_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdSplit_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdSplit_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdSplit_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdSplit_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdSplit_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdSplit_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdSplit_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdSplit_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdSplit_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdSplit_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdSplit_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdSplit_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdSplit_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdSplit_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdSplit_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdSplit_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdSplit_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdSplit_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdSplit_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdSplit_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdSplit_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdSplit_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdSplit_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdSplit_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdSplit_io_out_wdata_bits_wstrb_63),
    .io_out_rresp_ready(AXICmdSplit_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdSplit_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdSplit_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdSplit_io_out_wresp_bits_tag)
  );
  AXICmdIssue AXICmdIssue ( // @[DRAMArbiter.scala 97:26:@63424.4]
    .clock(AXICmdIssue_clock),
    .reset(AXICmdIssue_reset),
    .io_in_cmd_ready(AXICmdIssue_io_in_cmd_ready),
    .io_in_cmd_valid(AXICmdIssue_io_in_cmd_valid),
    .io_in_cmd_bits_addr(AXICmdIssue_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(AXICmdIssue_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(AXICmdIssue_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(AXICmdIssue_io_in_cmd_bits_tag),
    .io_in_wdata_ready(AXICmdIssue_io_in_wdata_ready),
    .io_in_wdata_valid(AXICmdIssue_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(AXICmdIssue_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(AXICmdIssue_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(AXICmdIssue_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(AXICmdIssue_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(AXICmdIssue_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(AXICmdIssue_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(AXICmdIssue_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(AXICmdIssue_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(AXICmdIssue_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(AXICmdIssue_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(AXICmdIssue_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(AXICmdIssue_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(AXICmdIssue_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(AXICmdIssue_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(AXICmdIssue_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(AXICmdIssue_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(AXICmdIssue_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(AXICmdIssue_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(AXICmdIssue_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(AXICmdIssue_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(AXICmdIssue_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(AXICmdIssue_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(AXICmdIssue_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(AXICmdIssue_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(AXICmdIssue_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(AXICmdIssue_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(AXICmdIssue_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(AXICmdIssue_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(AXICmdIssue_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(AXICmdIssue_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(AXICmdIssue_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(AXICmdIssue_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(AXICmdIssue_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(AXICmdIssue_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(AXICmdIssue_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(AXICmdIssue_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(AXICmdIssue_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(AXICmdIssue_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(AXICmdIssue_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(AXICmdIssue_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(AXICmdIssue_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(AXICmdIssue_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(AXICmdIssue_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(AXICmdIssue_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(AXICmdIssue_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(AXICmdIssue_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(AXICmdIssue_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(AXICmdIssue_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(AXICmdIssue_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(AXICmdIssue_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(AXICmdIssue_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(AXICmdIssue_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(AXICmdIssue_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(AXICmdIssue_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(AXICmdIssue_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(AXICmdIssue_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(AXICmdIssue_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(AXICmdIssue_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(AXICmdIssue_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(AXICmdIssue_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(AXICmdIssue_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(AXICmdIssue_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(AXICmdIssue_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(AXICmdIssue_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(AXICmdIssue_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(AXICmdIssue_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(AXICmdIssue_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(AXICmdIssue_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(AXICmdIssue_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(AXICmdIssue_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(AXICmdIssue_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(AXICmdIssue_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(AXICmdIssue_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(AXICmdIssue_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(AXICmdIssue_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(AXICmdIssue_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(AXICmdIssue_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(AXICmdIssue_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(AXICmdIssue_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(AXICmdIssue_io_in_wdata_bits_wstrb_63),
    .io_in_rresp_ready(AXICmdIssue_io_in_rresp_ready),
    .io_in_wresp_ready(AXICmdIssue_io_in_wresp_ready),
    .io_in_wresp_valid(AXICmdIssue_io_in_wresp_valid),
    .io_in_wresp_bits_tag(AXICmdIssue_io_in_wresp_bits_tag),
    .io_out_cmd_ready(AXICmdIssue_io_out_cmd_ready),
    .io_out_cmd_valid(AXICmdIssue_io_out_cmd_valid),
    .io_out_cmd_bits_addr(AXICmdIssue_io_out_cmd_bits_addr),
    .io_out_cmd_bits_size(AXICmdIssue_io_out_cmd_bits_size),
    .io_out_cmd_bits_isWr(AXICmdIssue_io_out_cmd_bits_isWr),
    .io_out_cmd_bits_tag(AXICmdIssue_io_out_cmd_bits_tag),
    .io_out_wdata_ready(AXICmdIssue_io_out_wdata_ready),
    .io_out_wdata_valid(AXICmdIssue_io_out_wdata_valid),
    .io_out_wdata_bits_wdata_0(AXICmdIssue_io_out_wdata_bits_wdata_0),
    .io_out_wdata_bits_wdata_1(AXICmdIssue_io_out_wdata_bits_wdata_1),
    .io_out_wdata_bits_wdata_2(AXICmdIssue_io_out_wdata_bits_wdata_2),
    .io_out_wdata_bits_wdata_3(AXICmdIssue_io_out_wdata_bits_wdata_3),
    .io_out_wdata_bits_wdata_4(AXICmdIssue_io_out_wdata_bits_wdata_4),
    .io_out_wdata_bits_wdata_5(AXICmdIssue_io_out_wdata_bits_wdata_5),
    .io_out_wdata_bits_wdata_6(AXICmdIssue_io_out_wdata_bits_wdata_6),
    .io_out_wdata_bits_wdata_7(AXICmdIssue_io_out_wdata_bits_wdata_7),
    .io_out_wdata_bits_wdata_8(AXICmdIssue_io_out_wdata_bits_wdata_8),
    .io_out_wdata_bits_wdata_9(AXICmdIssue_io_out_wdata_bits_wdata_9),
    .io_out_wdata_bits_wdata_10(AXICmdIssue_io_out_wdata_bits_wdata_10),
    .io_out_wdata_bits_wdata_11(AXICmdIssue_io_out_wdata_bits_wdata_11),
    .io_out_wdata_bits_wdata_12(AXICmdIssue_io_out_wdata_bits_wdata_12),
    .io_out_wdata_bits_wdata_13(AXICmdIssue_io_out_wdata_bits_wdata_13),
    .io_out_wdata_bits_wdata_14(AXICmdIssue_io_out_wdata_bits_wdata_14),
    .io_out_wdata_bits_wdata_15(AXICmdIssue_io_out_wdata_bits_wdata_15),
    .io_out_wdata_bits_wstrb_0(AXICmdIssue_io_out_wdata_bits_wstrb_0),
    .io_out_wdata_bits_wstrb_1(AXICmdIssue_io_out_wdata_bits_wstrb_1),
    .io_out_wdata_bits_wstrb_2(AXICmdIssue_io_out_wdata_bits_wstrb_2),
    .io_out_wdata_bits_wstrb_3(AXICmdIssue_io_out_wdata_bits_wstrb_3),
    .io_out_wdata_bits_wstrb_4(AXICmdIssue_io_out_wdata_bits_wstrb_4),
    .io_out_wdata_bits_wstrb_5(AXICmdIssue_io_out_wdata_bits_wstrb_5),
    .io_out_wdata_bits_wstrb_6(AXICmdIssue_io_out_wdata_bits_wstrb_6),
    .io_out_wdata_bits_wstrb_7(AXICmdIssue_io_out_wdata_bits_wstrb_7),
    .io_out_wdata_bits_wstrb_8(AXICmdIssue_io_out_wdata_bits_wstrb_8),
    .io_out_wdata_bits_wstrb_9(AXICmdIssue_io_out_wdata_bits_wstrb_9),
    .io_out_wdata_bits_wstrb_10(AXICmdIssue_io_out_wdata_bits_wstrb_10),
    .io_out_wdata_bits_wstrb_11(AXICmdIssue_io_out_wdata_bits_wstrb_11),
    .io_out_wdata_bits_wstrb_12(AXICmdIssue_io_out_wdata_bits_wstrb_12),
    .io_out_wdata_bits_wstrb_13(AXICmdIssue_io_out_wdata_bits_wstrb_13),
    .io_out_wdata_bits_wstrb_14(AXICmdIssue_io_out_wdata_bits_wstrb_14),
    .io_out_wdata_bits_wstrb_15(AXICmdIssue_io_out_wdata_bits_wstrb_15),
    .io_out_wdata_bits_wstrb_16(AXICmdIssue_io_out_wdata_bits_wstrb_16),
    .io_out_wdata_bits_wstrb_17(AXICmdIssue_io_out_wdata_bits_wstrb_17),
    .io_out_wdata_bits_wstrb_18(AXICmdIssue_io_out_wdata_bits_wstrb_18),
    .io_out_wdata_bits_wstrb_19(AXICmdIssue_io_out_wdata_bits_wstrb_19),
    .io_out_wdata_bits_wstrb_20(AXICmdIssue_io_out_wdata_bits_wstrb_20),
    .io_out_wdata_bits_wstrb_21(AXICmdIssue_io_out_wdata_bits_wstrb_21),
    .io_out_wdata_bits_wstrb_22(AXICmdIssue_io_out_wdata_bits_wstrb_22),
    .io_out_wdata_bits_wstrb_23(AXICmdIssue_io_out_wdata_bits_wstrb_23),
    .io_out_wdata_bits_wstrb_24(AXICmdIssue_io_out_wdata_bits_wstrb_24),
    .io_out_wdata_bits_wstrb_25(AXICmdIssue_io_out_wdata_bits_wstrb_25),
    .io_out_wdata_bits_wstrb_26(AXICmdIssue_io_out_wdata_bits_wstrb_26),
    .io_out_wdata_bits_wstrb_27(AXICmdIssue_io_out_wdata_bits_wstrb_27),
    .io_out_wdata_bits_wstrb_28(AXICmdIssue_io_out_wdata_bits_wstrb_28),
    .io_out_wdata_bits_wstrb_29(AXICmdIssue_io_out_wdata_bits_wstrb_29),
    .io_out_wdata_bits_wstrb_30(AXICmdIssue_io_out_wdata_bits_wstrb_30),
    .io_out_wdata_bits_wstrb_31(AXICmdIssue_io_out_wdata_bits_wstrb_31),
    .io_out_wdata_bits_wstrb_32(AXICmdIssue_io_out_wdata_bits_wstrb_32),
    .io_out_wdata_bits_wstrb_33(AXICmdIssue_io_out_wdata_bits_wstrb_33),
    .io_out_wdata_bits_wstrb_34(AXICmdIssue_io_out_wdata_bits_wstrb_34),
    .io_out_wdata_bits_wstrb_35(AXICmdIssue_io_out_wdata_bits_wstrb_35),
    .io_out_wdata_bits_wstrb_36(AXICmdIssue_io_out_wdata_bits_wstrb_36),
    .io_out_wdata_bits_wstrb_37(AXICmdIssue_io_out_wdata_bits_wstrb_37),
    .io_out_wdata_bits_wstrb_38(AXICmdIssue_io_out_wdata_bits_wstrb_38),
    .io_out_wdata_bits_wstrb_39(AXICmdIssue_io_out_wdata_bits_wstrb_39),
    .io_out_wdata_bits_wstrb_40(AXICmdIssue_io_out_wdata_bits_wstrb_40),
    .io_out_wdata_bits_wstrb_41(AXICmdIssue_io_out_wdata_bits_wstrb_41),
    .io_out_wdata_bits_wstrb_42(AXICmdIssue_io_out_wdata_bits_wstrb_42),
    .io_out_wdata_bits_wstrb_43(AXICmdIssue_io_out_wdata_bits_wstrb_43),
    .io_out_wdata_bits_wstrb_44(AXICmdIssue_io_out_wdata_bits_wstrb_44),
    .io_out_wdata_bits_wstrb_45(AXICmdIssue_io_out_wdata_bits_wstrb_45),
    .io_out_wdata_bits_wstrb_46(AXICmdIssue_io_out_wdata_bits_wstrb_46),
    .io_out_wdata_bits_wstrb_47(AXICmdIssue_io_out_wdata_bits_wstrb_47),
    .io_out_wdata_bits_wstrb_48(AXICmdIssue_io_out_wdata_bits_wstrb_48),
    .io_out_wdata_bits_wstrb_49(AXICmdIssue_io_out_wdata_bits_wstrb_49),
    .io_out_wdata_bits_wstrb_50(AXICmdIssue_io_out_wdata_bits_wstrb_50),
    .io_out_wdata_bits_wstrb_51(AXICmdIssue_io_out_wdata_bits_wstrb_51),
    .io_out_wdata_bits_wstrb_52(AXICmdIssue_io_out_wdata_bits_wstrb_52),
    .io_out_wdata_bits_wstrb_53(AXICmdIssue_io_out_wdata_bits_wstrb_53),
    .io_out_wdata_bits_wstrb_54(AXICmdIssue_io_out_wdata_bits_wstrb_54),
    .io_out_wdata_bits_wstrb_55(AXICmdIssue_io_out_wdata_bits_wstrb_55),
    .io_out_wdata_bits_wstrb_56(AXICmdIssue_io_out_wdata_bits_wstrb_56),
    .io_out_wdata_bits_wstrb_57(AXICmdIssue_io_out_wdata_bits_wstrb_57),
    .io_out_wdata_bits_wstrb_58(AXICmdIssue_io_out_wdata_bits_wstrb_58),
    .io_out_wdata_bits_wstrb_59(AXICmdIssue_io_out_wdata_bits_wstrb_59),
    .io_out_wdata_bits_wstrb_60(AXICmdIssue_io_out_wdata_bits_wstrb_60),
    .io_out_wdata_bits_wstrb_61(AXICmdIssue_io_out_wdata_bits_wstrb_61),
    .io_out_wdata_bits_wstrb_62(AXICmdIssue_io_out_wdata_bits_wstrb_62),
    .io_out_wdata_bits_wstrb_63(AXICmdIssue_io_out_wdata_bits_wstrb_63),
    .io_out_wdata_bits_wlast(AXICmdIssue_io_out_wdata_bits_wlast),
    .io_out_rresp_ready(AXICmdIssue_io_out_rresp_ready),
    .io_out_wresp_ready(AXICmdIssue_io_out_wresp_ready),
    .io_out_wresp_valid(AXICmdIssue_io_out_wresp_valid),
    .io_out_wresp_bits_tag(AXICmdIssue_io_out_wresp_bits_tag)
  );
  assign io_dram_cmd_valid = io_enable & AXICmdIssue_io_out_cmd_valid; // @[DRAMArbiter.scala 99:13:@63649.4 DRAMArbiter.scala 100:23:@63652.4]
  assign io_dram_cmd_bits_addr = AXICmdIssue_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 99:13:@63648.4]
  assign io_dram_cmd_bits_size = AXICmdIssue_io_out_cmd_bits_size; // @[DRAMArbiter.scala 99:13:@63647.4]
  assign io_dram_cmd_bits_isWr = AXICmdIssue_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 99:13:@63645.4]
  assign io_dram_cmd_bits_tag = AXICmdIssue_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 99:13:@63644.4]
  assign io_dram_wdata_valid = io_enable & AXICmdIssue_io_out_wdata_valid; // @[DRAMArbiter.scala 99:13:@63642.4 DRAMArbiter.scala 101:25:@63654.4]
  assign io_dram_wdata_bits_wdata_0 = AXICmdIssue_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 99:13:@63626.4]
  assign io_dram_wdata_bits_wdata_1 = AXICmdIssue_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 99:13:@63627.4]
  assign io_dram_wdata_bits_wdata_2 = AXICmdIssue_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 99:13:@63628.4]
  assign io_dram_wdata_bits_wdata_3 = AXICmdIssue_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 99:13:@63629.4]
  assign io_dram_wdata_bits_wdata_4 = AXICmdIssue_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 99:13:@63630.4]
  assign io_dram_wdata_bits_wdata_5 = AXICmdIssue_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 99:13:@63631.4]
  assign io_dram_wdata_bits_wdata_6 = AXICmdIssue_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 99:13:@63632.4]
  assign io_dram_wdata_bits_wdata_7 = AXICmdIssue_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 99:13:@63633.4]
  assign io_dram_wdata_bits_wdata_8 = AXICmdIssue_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 99:13:@63634.4]
  assign io_dram_wdata_bits_wdata_9 = AXICmdIssue_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 99:13:@63635.4]
  assign io_dram_wdata_bits_wdata_10 = AXICmdIssue_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 99:13:@63636.4]
  assign io_dram_wdata_bits_wdata_11 = AXICmdIssue_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 99:13:@63637.4]
  assign io_dram_wdata_bits_wdata_12 = AXICmdIssue_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 99:13:@63638.4]
  assign io_dram_wdata_bits_wdata_13 = AXICmdIssue_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 99:13:@63639.4]
  assign io_dram_wdata_bits_wdata_14 = AXICmdIssue_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 99:13:@63640.4]
  assign io_dram_wdata_bits_wdata_15 = AXICmdIssue_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 99:13:@63641.4]
  assign io_dram_wdata_bits_wstrb_0 = AXICmdIssue_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 99:13:@63562.4]
  assign io_dram_wdata_bits_wstrb_1 = AXICmdIssue_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 99:13:@63563.4]
  assign io_dram_wdata_bits_wstrb_2 = AXICmdIssue_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 99:13:@63564.4]
  assign io_dram_wdata_bits_wstrb_3 = AXICmdIssue_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 99:13:@63565.4]
  assign io_dram_wdata_bits_wstrb_4 = AXICmdIssue_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 99:13:@63566.4]
  assign io_dram_wdata_bits_wstrb_5 = AXICmdIssue_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 99:13:@63567.4]
  assign io_dram_wdata_bits_wstrb_6 = AXICmdIssue_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 99:13:@63568.4]
  assign io_dram_wdata_bits_wstrb_7 = AXICmdIssue_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 99:13:@63569.4]
  assign io_dram_wdata_bits_wstrb_8 = AXICmdIssue_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 99:13:@63570.4]
  assign io_dram_wdata_bits_wstrb_9 = AXICmdIssue_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 99:13:@63571.4]
  assign io_dram_wdata_bits_wstrb_10 = AXICmdIssue_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 99:13:@63572.4]
  assign io_dram_wdata_bits_wstrb_11 = AXICmdIssue_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 99:13:@63573.4]
  assign io_dram_wdata_bits_wstrb_12 = AXICmdIssue_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 99:13:@63574.4]
  assign io_dram_wdata_bits_wstrb_13 = AXICmdIssue_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 99:13:@63575.4]
  assign io_dram_wdata_bits_wstrb_14 = AXICmdIssue_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 99:13:@63576.4]
  assign io_dram_wdata_bits_wstrb_15 = AXICmdIssue_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 99:13:@63577.4]
  assign io_dram_wdata_bits_wstrb_16 = AXICmdIssue_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 99:13:@63578.4]
  assign io_dram_wdata_bits_wstrb_17 = AXICmdIssue_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 99:13:@63579.4]
  assign io_dram_wdata_bits_wstrb_18 = AXICmdIssue_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 99:13:@63580.4]
  assign io_dram_wdata_bits_wstrb_19 = AXICmdIssue_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 99:13:@63581.4]
  assign io_dram_wdata_bits_wstrb_20 = AXICmdIssue_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 99:13:@63582.4]
  assign io_dram_wdata_bits_wstrb_21 = AXICmdIssue_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 99:13:@63583.4]
  assign io_dram_wdata_bits_wstrb_22 = AXICmdIssue_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 99:13:@63584.4]
  assign io_dram_wdata_bits_wstrb_23 = AXICmdIssue_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 99:13:@63585.4]
  assign io_dram_wdata_bits_wstrb_24 = AXICmdIssue_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 99:13:@63586.4]
  assign io_dram_wdata_bits_wstrb_25 = AXICmdIssue_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 99:13:@63587.4]
  assign io_dram_wdata_bits_wstrb_26 = AXICmdIssue_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 99:13:@63588.4]
  assign io_dram_wdata_bits_wstrb_27 = AXICmdIssue_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 99:13:@63589.4]
  assign io_dram_wdata_bits_wstrb_28 = AXICmdIssue_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 99:13:@63590.4]
  assign io_dram_wdata_bits_wstrb_29 = AXICmdIssue_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 99:13:@63591.4]
  assign io_dram_wdata_bits_wstrb_30 = AXICmdIssue_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 99:13:@63592.4]
  assign io_dram_wdata_bits_wstrb_31 = AXICmdIssue_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 99:13:@63593.4]
  assign io_dram_wdata_bits_wstrb_32 = AXICmdIssue_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 99:13:@63594.4]
  assign io_dram_wdata_bits_wstrb_33 = AXICmdIssue_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 99:13:@63595.4]
  assign io_dram_wdata_bits_wstrb_34 = AXICmdIssue_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 99:13:@63596.4]
  assign io_dram_wdata_bits_wstrb_35 = AXICmdIssue_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 99:13:@63597.4]
  assign io_dram_wdata_bits_wstrb_36 = AXICmdIssue_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 99:13:@63598.4]
  assign io_dram_wdata_bits_wstrb_37 = AXICmdIssue_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 99:13:@63599.4]
  assign io_dram_wdata_bits_wstrb_38 = AXICmdIssue_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 99:13:@63600.4]
  assign io_dram_wdata_bits_wstrb_39 = AXICmdIssue_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 99:13:@63601.4]
  assign io_dram_wdata_bits_wstrb_40 = AXICmdIssue_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 99:13:@63602.4]
  assign io_dram_wdata_bits_wstrb_41 = AXICmdIssue_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 99:13:@63603.4]
  assign io_dram_wdata_bits_wstrb_42 = AXICmdIssue_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 99:13:@63604.4]
  assign io_dram_wdata_bits_wstrb_43 = AXICmdIssue_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 99:13:@63605.4]
  assign io_dram_wdata_bits_wstrb_44 = AXICmdIssue_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 99:13:@63606.4]
  assign io_dram_wdata_bits_wstrb_45 = AXICmdIssue_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 99:13:@63607.4]
  assign io_dram_wdata_bits_wstrb_46 = AXICmdIssue_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 99:13:@63608.4]
  assign io_dram_wdata_bits_wstrb_47 = AXICmdIssue_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 99:13:@63609.4]
  assign io_dram_wdata_bits_wstrb_48 = AXICmdIssue_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 99:13:@63610.4]
  assign io_dram_wdata_bits_wstrb_49 = AXICmdIssue_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 99:13:@63611.4]
  assign io_dram_wdata_bits_wstrb_50 = AXICmdIssue_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 99:13:@63612.4]
  assign io_dram_wdata_bits_wstrb_51 = AXICmdIssue_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 99:13:@63613.4]
  assign io_dram_wdata_bits_wstrb_52 = AXICmdIssue_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 99:13:@63614.4]
  assign io_dram_wdata_bits_wstrb_53 = AXICmdIssue_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 99:13:@63615.4]
  assign io_dram_wdata_bits_wstrb_54 = AXICmdIssue_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 99:13:@63616.4]
  assign io_dram_wdata_bits_wstrb_55 = AXICmdIssue_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 99:13:@63617.4]
  assign io_dram_wdata_bits_wstrb_56 = AXICmdIssue_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 99:13:@63618.4]
  assign io_dram_wdata_bits_wstrb_57 = AXICmdIssue_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 99:13:@63619.4]
  assign io_dram_wdata_bits_wstrb_58 = AXICmdIssue_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 99:13:@63620.4]
  assign io_dram_wdata_bits_wstrb_59 = AXICmdIssue_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 99:13:@63621.4]
  assign io_dram_wdata_bits_wstrb_60 = AXICmdIssue_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 99:13:@63622.4]
  assign io_dram_wdata_bits_wstrb_61 = AXICmdIssue_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 99:13:@63623.4]
  assign io_dram_wdata_bits_wstrb_62 = AXICmdIssue_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 99:13:@63624.4]
  assign io_dram_wdata_bits_wstrb_63 = AXICmdIssue_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 99:13:@63625.4]
  assign io_dram_wdata_bits_wlast = AXICmdIssue_io_out_wdata_bits_wlast; // @[DRAMArbiter.scala 99:13:@63561.4]
  assign io_dram_rresp_ready = AXICmdIssue_io_out_rresp_ready; // @[DRAMArbiter.scala 99:13:@63560.4]
  assign io_dram_wresp_ready = AXICmdIssue_io_out_wresp_ready; // @[DRAMArbiter.scala 99:13:@63541.4]
  assign StreamControllerStore_clock = clock; // @[:@63068.4]
  assign StreamControllerStore_reset = reset; // @[:@63069.4]
  assign StreamControllerStore_io_dram_cmd_ready = StreamArbiter_io_app_0_cmd_ready; // @[DRAMArbiter.scala 87:32:@63196.4]
  assign StreamControllerStore_io_dram_wdata_ready = StreamArbiter_io_app_0_wdata_ready; // @[DRAMArbiter.scala 87:32:@63189.4]
  assign StreamControllerStore_io_dram_wresp_valid = StreamArbiter_io_app_0_wresp_valid; // @[DRAMArbiter.scala 87:32:@63086.4]
  assign StreamControllerStore_io_store_cmd_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@63079.4]
  assign StreamControllerStore_io_store_cmd_bits_addr = 64'h0; // @[DRAMArbiter.scala 68:18:@63078.4]
  assign StreamControllerStore_io_store_cmd_bits_size = 32'h0; // @[DRAMArbiter.scala 68:18:@63077.4]
  assign StreamControllerStore_io_store_data_valid = 1'h0; // @[DRAMArbiter.scala 68:18:@63075.4]
  assign StreamControllerStore_io_store_data_bits_wdata_0 = 32'h0; // @[DRAMArbiter.scala 68:18:@63074.4]
  assign StreamControllerStore_io_store_data_bits_wstrb = 1'h0; // @[DRAMArbiter.scala 68:18:@63073.4]
  assign StreamControllerStore_io_store_wresp_ready = 1'h0; // @[DRAMArbiter.scala 68:18:@63072.4]
  assign StreamArbiter_clock = clock; // @[:@63082.4]
  assign StreamArbiter_reset = reset; // @[:@63083.4]
  assign StreamArbiter_io_app_0_cmd_valid = StreamControllerStore_io_dram_cmd_valid; // @[DRAMArbiter.scala 87:22:@63307.4]
  assign StreamArbiter_io_app_0_cmd_bits_addr = StreamControllerStore_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 87:22:@63306.4]
  assign StreamArbiter_io_app_0_cmd_bits_size = StreamControllerStore_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 87:22:@63305.4]
  assign StreamArbiter_io_app_0_cmd_bits_isWr = 1'h1; // @[DRAMArbiter.scala 87:22:@63303.4]
  assign StreamArbiter_io_app_0_cmd_bits_tag = 32'h0; // @[DRAMArbiter.scala 87:22:@63302.4]
  assign StreamArbiter_io_app_0_wdata_valid = StreamControllerStore_io_dram_wdata_valid; // @[DRAMArbiter.scala 87:22:@63300.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_0 = StreamControllerStore_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 87:22:@63284.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_1 = StreamControllerStore_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 87:22:@63285.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_2 = StreamControllerStore_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 87:22:@63286.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_3 = StreamControllerStore_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 87:22:@63287.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_4 = StreamControllerStore_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 87:22:@63288.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_5 = StreamControllerStore_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 87:22:@63289.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_6 = StreamControllerStore_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 87:22:@63290.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_7 = StreamControllerStore_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 87:22:@63291.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_8 = StreamControllerStore_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 87:22:@63292.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_9 = StreamControllerStore_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 87:22:@63293.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_10 = StreamControllerStore_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 87:22:@63294.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_11 = StreamControllerStore_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 87:22:@63295.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_12 = StreamControllerStore_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 87:22:@63296.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_13 = StreamControllerStore_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 87:22:@63297.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_14 = StreamControllerStore_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 87:22:@63298.4]
  assign StreamArbiter_io_app_0_wdata_bits_wdata_15 = StreamControllerStore_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 87:22:@63299.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_0 = StreamControllerStore_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 87:22:@63220.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_1 = StreamControllerStore_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 87:22:@63221.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_2 = StreamControllerStore_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 87:22:@63222.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_3 = StreamControllerStore_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 87:22:@63223.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_4 = StreamControllerStore_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 87:22:@63224.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_5 = StreamControllerStore_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 87:22:@63225.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_6 = StreamControllerStore_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 87:22:@63226.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_7 = StreamControllerStore_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 87:22:@63227.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_8 = StreamControllerStore_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 87:22:@63228.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_9 = StreamControllerStore_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 87:22:@63229.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_10 = StreamControllerStore_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 87:22:@63230.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_11 = StreamControllerStore_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 87:22:@63231.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_12 = StreamControllerStore_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 87:22:@63232.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_13 = StreamControllerStore_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 87:22:@63233.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_14 = StreamControllerStore_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 87:22:@63234.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_15 = StreamControllerStore_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 87:22:@63235.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_16 = StreamControllerStore_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 87:22:@63236.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_17 = StreamControllerStore_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 87:22:@63237.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_18 = StreamControllerStore_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 87:22:@63238.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_19 = StreamControllerStore_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 87:22:@63239.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_20 = StreamControllerStore_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 87:22:@63240.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_21 = StreamControllerStore_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 87:22:@63241.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_22 = StreamControllerStore_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 87:22:@63242.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_23 = StreamControllerStore_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 87:22:@63243.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_24 = StreamControllerStore_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 87:22:@63244.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_25 = StreamControllerStore_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 87:22:@63245.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_26 = StreamControllerStore_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 87:22:@63246.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_27 = StreamControllerStore_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 87:22:@63247.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_28 = StreamControllerStore_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 87:22:@63248.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_29 = StreamControllerStore_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 87:22:@63249.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_30 = StreamControllerStore_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 87:22:@63250.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_31 = StreamControllerStore_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 87:22:@63251.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_32 = StreamControllerStore_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 87:22:@63252.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_33 = StreamControllerStore_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 87:22:@63253.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_34 = StreamControllerStore_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 87:22:@63254.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_35 = StreamControllerStore_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 87:22:@63255.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_36 = StreamControllerStore_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 87:22:@63256.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_37 = StreamControllerStore_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 87:22:@63257.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_38 = StreamControllerStore_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 87:22:@63258.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_39 = StreamControllerStore_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 87:22:@63259.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_40 = StreamControllerStore_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 87:22:@63260.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_41 = StreamControllerStore_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 87:22:@63261.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_42 = StreamControllerStore_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 87:22:@63262.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_43 = StreamControllerStore_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 87:22:@63263.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_44 = StreamControllerStore_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 87:22:@63264.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_45 = StreamControllerStore_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 87:22:@63265.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_46 = StreamControllerStore_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 87:22:@63266.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_47 = StreamControllerStore_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 87:22:@63267.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_48 = StreamControllerStore_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 87:22:@63268.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_49 = StreamControllerStore_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 87:22:@63269.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_50 = StreamControllerStore_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 87:22:@63270.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_51 = StreamControllerStore_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 87:22:@63271.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_52 = StreamControllerStore_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 87:22:@63272.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_53 = StreamControllerStore_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 87:22:@63273.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_54 = StreamControllerStore_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 87:22:@63274.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_55 = StreamControllerStore_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 87:22:@63275.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_56 = StreamControllerStore_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 87:22:@63276.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_57 = StreamControllerStore_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 87:22:@63277.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_58 = StreamControllerStore_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 87:22:@63278.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_59 = StreamControllerStore_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 87:22:@63279.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_60 = StreamControllerStore_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 87:22:@63280.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_61 = StreamControllerStore_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 87:22:@63281.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_62 = StreamControllerStore_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 87:22:@63282.4]
  assign StreamArbiter_io_app_0_wdata_bits_wstrb_63 = StreamControllerStore_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 87:22:@63283.4]
  assign StreamArbiter_io_app_0_rresp_ready = 1'h0; // @[DRAMArbiter.scala 87:22:@63218.4]
  assign StreamArbiter_io_app_0_wresp_ready = StreamControllerStore_io_dram_wresp_ready; // @[DRAMArbiter.scala 87:22:@63199.4]
  assign StreamArbiter_io_dram_cmd_ready = AXICmdSplit_io_in_cmd_ready; // @[DRAMArbiter.scala 95:20:@63423.4]
  assign StreamArbiter_io_dram_wdata_ready = AXICmdSplit_io_in_wdata_ready; // @[DRAMArbiter.scala 95:20:@63416.4]
  assign StreamArbiter_io_dram_wresp_valid = AXICmdSplit_io_in_wresp_valid; // @[DRAMArbiter.scala 95:20:@63313.4]
  assign StreamArbiter_io_dram_wresp_bits_tag = AXICmdSplit_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 95:20:@63312.4]
  assign AXICmdSplit_clock = clock; // @[:@63310.4]
  assign AXICmdSplit_reset = reset; // @[:@63311.4]
  assign AXICmdSplit_io_in_cmd_valid = StreamArbiter_io_dram_cmd_valid; // @[DRAMArbiter.scala 95:20:@63422.4]
  assign AXICmdSplit_io_in_cmd_bits_addr = StreamArbiter_io_dram_cmd_bits_addr; // @[DRAMArbiter.scala 95:20:@63421.4]
  assign AXICmdSplit_io_in_cmd_bits_size = StreamArbiter_io_dram_cmd_bits_size; // @[DRAMArbiter.scala 95:20:@63420.4]
  assign AXICmdSplit_io_in_cmd_bits_isWr = StreamArbiter_io_dram_cmd_bits_isWr; // @[DRAMArbiter.scala 95:20:@63418.4]
  assign AXICmdSplit_io_in_cmd_bits_tag = StreamArbiter_io_dram_cmd_bits_tag; // @[DRAMArbiter.scala 95:20:@63417.4]
  assign AXICmdSplit_io_in_wdata_valid = StreamArbiter_io_dram_wdata_valid; // @[DRAMArbiter.scala 95:20:@63415.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_0 = StreamArbiter_io_dram_wdata_bits_wdata_0; // @[DRAMArbiter.scala 95:20:@63399.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_1 = StreamArbiter_io_dram_wdata_bits_wdata_1; // @[DRAMArbiter.scala 95:20:@63400.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_2 = StreamArbiter_io_dram_wdata_bits_wdata_2; // @[DRAMArbiter.scala 95:20:@63401.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_3 = StreamArbiter_io_dram_wdata_bits_wdata_3; // @[DRAMArbiter.scala 95:20:@63402.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_4 = StreamArbiter_io_dram_wdata_bits_wdata_4; // @[DRAMArbiter.scala 95:20:@63403.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_5 = StreamArbiter_io_dram_wdata_bits_wdata_5; // @[DRAMArbiter.scala 95:20:@63404.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_6 = StreamArbiter_io_dram_wdata_bits_wdata_6; // @[DRAMArbiter.scala 95:20:@63405.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_7 = StreamArbiter_io_dram_wdata_bits_wdata_7; // @[DRAMArbiter.scala 95:20:@63406.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_8 = StreamArbiter_io_dram_wdata_bits_wdata_8; // @[DRAMArbiter.scala 95:20:@63407.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_9 = StreamArbiter_io_dram_wdata_bits_wdata_9; // @[DRAMArbiter.scala 95:20:@63408.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_10 = StreamArbiter_io_dram_wdata_bits_wdata_10; // @[DRAMArbiter.scala 95:20:@63409.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_11 = StreamArbiter_io_dram_wdata_bits_wdata_11; // @[DRAMArbiter.scala 95:20:@63410.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_12 = StreamArbiter_io_dram_wdata_bits_wdata_12; // @[DRAMArbiter.scala 95:20:@63411.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_13 = StreamArbiter_io_dram_wdata_bits_wdata_13; // @[DRAMArbiter.scala 95:20:@63412.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_14 = StreamArbiter_io_dram_wdata_bits_wdata_14; // @[DRAMArbiter.scala 95:20:@63413.4]
  assign AXICmdSplit_io_in_wdata_bits_wdata_15 = StreamArbiter_io_dram_wdata_bits_wdata_15; // @[DRAMArbiter.scala 95:20:@63414.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_0 = StreamArbiter_io_dram_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 95:20:@63335.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_1 = StreamArbiter_io_dram_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 95:20:@63336.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_2 = StreamArbiter_io_dram_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 95:20:@63337.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_3 = StreamArbiter_io_dram_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 95:20:@63338.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_4 = StreamArbiter_io_dram_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 95:20:@63339.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_5 = StreamArbiter_io_dram_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 95:20:@63340.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_6 = StreamArbiter_io_dram_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 95:20:@63341.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_7 = StreamArbiter_io_dram_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 95:20:@63342.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_8 = StreamArbiter_io_dram_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 95:20:@63343.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_9 = StreamArbiter_io_dram_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 95:20:@63344.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_10 = StreamArbiter_io_dram_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 95:20:@63345.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_11 = StreamArbiter_io_dram_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 95:20:@63346.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_12 = StreamArbiter_io_dram_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 95:20:@63347.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_13 = StreamArbiter_io_dram_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 95:20:@63348.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_14 = StreamArbiter_io_dram_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 95:20:@63349.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_15 = StreamArbiter_io_dram_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 95:20:@63350.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_16 = StreamArbiter_io_dram_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 95:20:@63351.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_17 = StreamArbiter_io_dram_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 95:20:@63352.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_18 = StreamArbiter_io_dram_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 95:20:@63353.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_19 = StreamArbiter_io_dram_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 95:20:@63354.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_20 = StreamArbiter_io_dram_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 95:20:@63355.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_21 = StreamArbiter_io_dram_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 95:20:@63356.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_22 = StreamArbiter_io_dram_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 95:20:@63357.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_23 = StreamArbiter_io_dram_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 95:20:@63358.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_24 = StreamArbiter_io_dram_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 95:20:@63359.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_25 = StreamArbiter_io_dram_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 95:20:@63360.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_26 = StreamArbiter_io_dram_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 95:20:@63361.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_27 = StreamArbiter_io_dram_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 95:20:@63362.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_28 = StreamArbiter_io_dram_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 95:20:@63363.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_29 = StreamArbiter_io_dram_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 95:20:@63364.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_30 = StreamArbiter_io_dram_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 95:20:@63365.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_31 = StreamArbiter_io_dram_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 95:20:@63366.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_32 = StreamArbiter_io_dram_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 95:20:@63367.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_33 = StreamArbiter_io_dram_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 95:20:@63368.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_34 = StreamArbiter_io_dram_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 95:20:@63369.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_35 = StreamArbiter_io_dram_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 95:20:@63370.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_36 = StreamArbiter_io_dram_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 95:20:@63371.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_37 = StreamArbiter_io_dram_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 95:20:@63372.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_38 = StreamArbiter_io_dram_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 95:20:@63373.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_39 = StreamArbiter_io_dram_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 95:20:@63374.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_40 = StreamArbiter_io_dram_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 95:20:@63375.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_41 = StreamArbiter_io_dram_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 95:20:@63376.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_42 = StreamArbiter_io_dram_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 95:20:@63377.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_43 = StreamArbiter_io_dram_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 95:20:@63378.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_44 = StreamArbiter_io_dram_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 95:20:@63379.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_45 = StreamArbiter_io_dram_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 95:20:@63380.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_46 = StreamArbiter_io_dram_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 95:20:@63381.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_47 = StreamArbiter_io_dram_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 95:20:@63382.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_48 = StreamArbiter_io_dram_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 95:20:@63383.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_49 = StreamArbiter_io_dram_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 95:20:@63384.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_50 = StreamArbiter_io_dram_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 95:20:@63385.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_51 = StreamArbiter_io_dram_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 95:20:@63386.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_52 = StreamArbiter_io_dram_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 95:20:@63387.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_53 = StreamArbiter_io_dram_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 95:20:@63388.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_54 = StreamArbiter_io_dram_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 95:20:@63389.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_55 = StreamArbiter_io_dram_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 95:20:@63390.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_56 = StreamArbiter_io_dram_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 95:20:@63391.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_57 = StreamArbiter_io_dram_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 95:20:@63392.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_58 = StreamArbiter_io_dram_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 95:20:@63393.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_59 = StreamArbiter_io_dram_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 95:20:@63394.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_60 = StreamArbiter_io_dram_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 95:20:@63395.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_61 = StreamArbiter_io_dram_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 95:20:@63396.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_62 = StreamArbiter_io_dram_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 95:20:@63397.4]
  assign AXICmdSplit_io_in_wdata_bits_wstrb_63 = StreamArbiter_io_dram_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 95:20:@63398.4]
  assign AXICmdSplit_io_in_rresp_ready = StreamArbiter_io_dram_rresp_ready; // @[DRAMArbiter.scala 95:20:@63333.4]
  assign AXICmdSplit_io_in_wresp_ready = StreamArbiter_io_dram_wresp_ready; // @[DRAMArbiter.scala 95:20:@63314.4]
  assign AXICmdSplit_io_out_cmd_ready = AXICmdIssue_io_in_cmd_ready; // @[DRAMArbiter.scala 98:20:@63538.4]
  assign AXICmdSplit_io_out_wdata_ready = AXICmdIssue_io_in_wdata_ready; // @[DRAMArbiter.scala 98:20:@63531.4]
  assign AXICmdSplit_io_out_wresp_valid = AXICmdIssue_io_in_wresp_valid; // @[DRAMArbiter.scala 98:20:@63428.4]
  assign AXICmdSplit_io_out_wresp_bits_tag = AXICmdIssue_io_in_wresp_bits_tag; // @[DRAMArbiter.scala 98:20:@63427.4]
  assign AXICmdIssue_clock = clock; // @[:@63425.4]
  assign AXICmdIssue_reset = reset; // @[:@63426.4]
  assign AXICmdIssue_io_in_cmd_valid = AXICmdSplit_io_out_cmd_valid; // @[DRAMArbiter.scala 98:20:@63537.4]
  assign AXICmdIssue_io_in_cmd_bits_addr = AXICmdSplit_io_out_cmd_bits_addr; // @[DRAMArbiter.scala 98:20:@63536.4]
  assign AXICmdIssue_io_in_cmd_bits_size = AXICmdSplit_io_out_cmd_bits_size; // @[DRAMArbiter.scala 98:20:@63535.4]
  assign AXICmdIssue_io_in_cmd_bits_isWr = AXICmdSplit_io_out_cmd_bits_isWr; // @[DRAMArbiter.scala 98:20:@63533.4]
  assign AXICmdIssue_io_in_cmd_bits_tag = AXICmdSplit_io_out_cmd_bits_tag; // @[DRAMArbiter.scala 98:20:@63532.4]
  assign AXICmdIssue_io_in_wdata_valid = AXICmdSplit_io_out_wdata_valid; // @[DRAMArbiter.scala 98:20:@63530.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_0 = AXICmdSplit_io_out_wdata_bits_wdata_0; // @[DRAMArbiter.scala 98:20:@63514.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_1 = AXICmdSplit_io_out_wdata_bits_wdata_1; // @[DRAMArbiter.scala 98:20:@63515.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_2 = AXICmdSplit_io_out_wdata_bits_wdata_2; // @[DRAMArbiter.scala 98:20:@63516.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_3 = AXICmdSplit_io_out_wdata_bits_wdata_3; // @[DRAMArbiter.scala 98:20:@63517.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_4 = AXICmdSplit_io_out_wdata_bits_wdata_4; // @[DRAMArbiter.scala 98:20:@63518.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_5 = AXICmdSplit_io_out_wdata_bits_wdata_5; // @[DRAMArbiter.scala 98:20:@63519.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_6 = AXICmdSplit_io_out_wdata_bits_wdata_6; // @[DRAMArbiter.scala 98:20:@63520.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_7 = AXICmdSplit_io_out_wdata_bits_wdata_7; // @[DRAMArbiter.scala 98:20:@63521.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_8 = AXICmdSplit_io_out_wdata_bits_wdata_8; // @[DRAMArbiter.scala 98:20:@63522.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_9 = AXICmdSplit_io_out_wdata_bits_wdata_9; // @[DRAMArbiter.scala 98:20:@63523.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_10 = AXICmdSplit_io_out_wdata_bits_wdata_10; // @[DRAMArbiter.scala 98:20:@63524.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_11 = AXICmdSplit_io_out_wdata_bits_wdata_11; // @[DRAMArbiter.scala 98:20:@63525.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_12 = AXICmdSplit_io_out_wdata_bits_wdata_12; // @[DRAMArbiter.scala 98:20:@63526.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_13 = AXICmdSplit_io_out_wdata_bits_wdata_13; // @[DRAMArbiter.scala 98:20:@63527.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_14 = AXICmdSplit_io_out_wdata_bits_wdata_14; // @[DRAMArbiter.scala 98:20:@63528.4]
  assign AXICmdIssue_io_in_wdata_bits_wdata_15 = AXICmdSplit_io_out_wdata_bits_wdata_15; // @[DRAMArbiter.scala 98:20:@63529.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_0 = AXICmdSplit_io_out_wdata_bits_wstrb_0; // @[DRAMArbiter.scala 98:20:@63450.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_1 = AXICmdSplit_io_out_wdata_bits_wstrb_1; // @[DRAMArbiter.scala 98:20:@63451.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_2 = AXICmdSplit_io_out_wdata_bits_wstrb_2; // @[DRAMArbiter.scala 98:20:@63452.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_3 = AXICmdSplit_io_out_wdata_bits_wstrb_3; // @[DRAMArbiter.scala 98:20:@63453.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_4 = AXICmdSplit_io_out_wdata_bits_wstrb_4; // @[DRAMArbiter.scala 98:20:@63454.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_5 = AXICmdSplit_io_out_wdata_bits_wstrb_5; // @[DRAMArbiter.scala 98:20:@63455.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_6 = AXICmdSplit_io_out_wdata_bits_wstrb_6; // @[DRAMArbiter.scala 98:20:@63456.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_7 = AXICmdSplit_io_out_wdata_bits_wstrb_7; // @[DRAMArbiter.scala 98:20:@63457.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_8 = AXICmdSplit_io_out_wdata_bits_wstrb_8; // @[DRAMArbiter.scala 98:20:@63458.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_9 = AXICmdSplit_io_out_wdata_bits_wstrb_9; // @[DRAMArbiter.scala 98:20:@63459.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_10 = AXICmdSplit_io_out_wdata_bits_wstrb_10; // @[DRAMArbiter.scala 98:20:@63460.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_11 = AXICmdSplit_io_out_wdata_bits_wstrb_11; // @[DRAMArbiter.scala 98:20:@63461.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_12 = AXICmdSplit_io_out_wdata_bits_wstrb_12; // @[DRAMArbiter.scala 98:20:@63462.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_13 = AXICmdSplit_io_out_wdata_bits_wstrb_13; // @[DRAMArbiter.scala 98:20:@63463.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_14 = AXICmdSplit_io_out_wdata_bits_wstrb_14; // @[DRAMArbiter.scala 98:20:@63464.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_15 = AXICmdSplit_io_out_wdata_bits_wstrb_15; // @[DRAMArbiter.scala 98:20:@63465.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_16 = AXICmdSplit_io_out_wdata_bits_wstrb_16; // @[DRAMArbiter.scala 98:20:@63466.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_17 = AXICmdSplit_io_out_wdata_bits_wstrb_17; // @[DRAMArbiter.scala 98:20:@63467.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_18 = AXICmdSplit_io_out_wdata_bits_wstrb_18; // @[DRAMArbiter.scala 98:20:@63468.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_19 = AXICmdSplit_io_out_wdata_bits_wstrb_19; // @[DRAMArbiter.scala 98:20:@63469.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_20 = AXICmdSplit_io_out_wdata_bits_wstrb_20; // @[DRAMArbiter.scala 98:20:@63470.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_21 = AXICmdSplit_io_out_wdata_bits_wstrb_21; // @[DRAMArbiter.scala 98:20:@63471.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_22 = AXICmdSplit_io_out_wdata_bits_wstrb_22; // @[DRAMArbiter.scala 98:20:@63472.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_23 = AXICmdSplit_io_out_wdata_bits_wstrb_23; // @[DRAMArbiter.scala 98:20:@63473.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_24 = AXICmdSplit_io_out_wdata_bits_wstrb_24; // @[DRAMArbiter.scala 98:20:@63474.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_25 = AXICmdSplit_io_out_wdata_bits_wstrb_25; // @[DRAMArbiter.scala 98:20:@63475.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_26 = AXICmdSplit_io_out_wdata_bits_wstrb_26; // @[DRAMArbiter.scala 98:20:@63476.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_27 = AXICmdSplit_io_out_wdata_bits_wstrb_27; // @[DRAMArbiter.scala 98:20:@63477.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_28 = AXICmdSplit_io_out_wdata_bits_wstrb_28; // @[DRAMArbiter.scala 98:20:@63478.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_29 = AXICmdSplit_io_out_wdata_bits_wstrb_29; // @[DRAMArbiter.scala 98:20:@63479.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_30 = AXICmdSplit_io_out_wdata_bits_wstrb_30; // @[DRAMArbiter.scala 98:20:@63480.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_31 = AXICmdSplit_io_out_wdata_bits_wstrb_31; // @[DRAMArbiter.scala 98:20:@63481.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_32 = AXICmdSplit_io_out_wdata_bits_wstrb_32; // @[DRAMArbiter.scala 98:20:@63482.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_33 = AXICmdSplit_io_out_wdata_bits_wstrb_33; // @[DRAMArbiter.scala 98:20:@63483.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_34 = AXICmdSplit_io_out_wdata_bits_wstrb_34; // @[DRAMArbiter.scala 98:20:@63484.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_35 = AXICmdSplit_io_out_wdata_bits_wstrb_35; // @[DRAMArbiter.scala 98:20:@63485.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_36 = AXICmdSplit_io_out_wdata_bits_wstrb_36; // @[DRAMArbiter.scala 98:20:@63486.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_37 = AXICmdSplit_io_out_wdata_bits_wstrb_37; // @[DRAMArbiter.scala 98:20:@63487.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_38 = AXICmdSplit_io_out_wdata_bits_wstrb_38; // @[DRAMArbiter.scala 98:20:@63488.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_39 = AXICmdSplit_io_out_wdata_bits_wstrb_39; // @[DRAMArbiter.scala 98:20:@63489.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_40 = AXICmdSplit_io_out_wdata_bits_wstrb_40; // @[DRAMArbiter.scala 98:20:@63490.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_41 = AXICmdSplit_io_out_wdata_bits_wstrb_41; // @[DRAMArbiter.scala 98:20:@63491.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_42 = AXICmdSplit_io_out_wdata_bits_wstrb_42; // @[DRAMArbiter.scala 98:20:@63492.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_43 = AXICmdSplit_io_out_wdata_bits_wstrb_43; // @[DRAMArbiter.scala 98:20:@63493.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_44 = AXICmdSplit_io_out_wdata_bits_wstrb_44; // @[DRAMArbiter.scala 98:20:@63494.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_45 = AXICmdSplit_io_out_wdata_bits_wstrb_45; // @[DRAMArbiter.scala 98:20:@63495.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_46 = AXICmdSplit_io_out_wdata_bits_wstrb_46; // @[DRAMArbiter.scala 98:20:@63496.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_47 = AXICmdSplit_io_out_wdata_bits_wstrb_47; // @[DRAMArbiter.scala 98:20:@63497.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_48 = AXICmdSplit_io_out_wdata_bits_wstrb_48; // @[DRAMArbiter.scala 98:20:@63498.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_49 = AXICmdSplit_io_out_wdata_bits_wstrb_49; // @[DRAMArbiter.scala 98:20:@63499.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_50 = AXICmdSplit_io_out_wdata_bits_wstrb_50; // @[DRAMArbiter.scala 98:20:@63500.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_51 = AXICmdSplit_io_out_wdata_bits_wstrb_51; // @[DRAMArbiter.scala 98:20:@63501.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_52 = AXICmdSplit_io_out_wdata_bits_wstrb_52; // @[DRAMArbiter.scala 98:20:@63502.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_53 = AXICmdSplit_io_out_wdata_bits_wstrb_53; // @[DRAMArbiter.scala 98:20:@63503.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_54 = AXICmdSplit_io_out_wdata_bits_wstrb_54; // @[DRAMArbiter.scala 98:20:@63504.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_55 = AXICmdSplit_io_out_wdata_bits_wstrb_55; // @[DRAMArbiter.scala 98:20:@63505.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_56 = AXICmdSplit_io_out_wdata_bits_wstrb_56; // @[DRAMArbiter.scala 98:20:@63506.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_57 = AXICmdSplit_io_out_wdata_bits_wstrb_57; // @[DRAMArbiter.scala 98:20:@63507.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_58 = AXICmdSplit_io_out_wdata_bits_wstrb_58; // @[DRAMArbiter.scala 98:20:@63508.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_59 = AXICmdSplit_io_out_wdata_bits_wstrb_59; // @[DRAMArbiter.scala 98:20:@63509.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_60 = AXICmdSplit_io_out_wdata_bits_wstrb_60; // @[DRAMArbiter.scala 98:20:@63510.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_61 = AXICmdSplit_io_out_wdata_bits_wstrb_61; // @[DRAMArbiter.scala 98:20:@63511.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_62 = AXICmdSplit_io_out_wdata_bits_wstrb_62; // @[DRAMArbiter.scala 98:20:@63512.4]
  assign AXICmdIssue_io_in_wdata_bits_wstrb_63 = AXICmdSplit_io_out_wdata_bits_wstrb_63; // @[DRAMArbiter.scala 98:20:@63513.4]
  assign AXICmdIssue_io_in_rresp_ready = AXICmdSplit_io_out_rresp_ready; // @[DRAMArbiter.scala 98:20:@63448.4]
  assign AXICmdIssue_io_in_wresp_ready = AXICmdSplit_io_out_wresp_ready; // @[DRAMArbiter.scala 98:20:@63429.4]
  assign AXICmdIssue_io_out_cmd_ready = io_dram_cmd_ready; // @[DRAMArbiter.scala 99:13:@63650.4]
  assign AXICmdIssue_io_out_wdata_ready = io_dram_wdata_ready; // @[DRAMArbiter.scala 99:13:@63643.4]
  assign AXICmdIssue_io_out_wresp_valid = io_dram_wresp_valid; // @[DRAMArbiter.scala 99:13:@63540.4]
  assign AXICmdIssue_io_out_wresp_bits_tag = io_dram_wresp_bits_tag; // @[DRAMArbiter.scala 99:13:@63539.4]
endmodule
module DRAMHeap( // @[:@94286.2]
  input         io_accel_0_req_valid, // @[:@94289.4]
  input         io_accel_0_req_bits_allocDealloc, // @[:@94289.4]
  input  [63:0] io_accel_0_req_bits_sizeAddr, // @[:@94289.4]
  output        io_accel_0_resp_valid, // @[:@94289.4]
  output        io_accel_0_resp_bits_allocDealloc, // @[:@94289.4]
  output [63:0] io_accel_0_resp_bits_sizeAddr, // @[:@94289.4]
  output        io_host_0_req_valid, // @[:@94289.4]
  output        io_host_0_req_bits_allocDealloc, // @[:@94289.4]
  output [63:0] io_host_0_req_bits_sizeAddr, // @[:@94289.4]
  input         io_host_0_resp_valid, // @[:@94289.4]
  input         io_host_0_resp_bits_allocDealloc, // @[:@94289.4]
  input  [63:0] io_host_0_resp_bits_sizeAddr // @[:@94289.4]
);
  assign io_accel_0_resp_valid = io_host_0_resp_valid; // @[DRAMHeap.scala 24:18:@94296.4]
  assign io_accel_0_resp_bits_allocDealloc = io_host_0_resp_bits_allocDealloc; // @[DRAMHeap.scala 25:17:@94298.4]
  assign io_accel_0_resp_bits_sizeAddr = io_host_0_resp_bits_sizeAddr; // @[DRAMHeap.scala 25:17:@94297.4]
  assign io_host_0_req_valid = io_accel_0_req_valid; // @[DRAMHeap.scala 21:18:@94293.4]
  assign io_host_0_req_bits_allocDealloc = io_accel_0_req_bits_allocDealloc; // @[DRAMHeap.scala 21:18:@94292.4]
  assign io_host_0_req_bits_sizeAddr = io_accel_0_req_bits_sizeAddr; // @[DRAMHeap.scala 21:18:@94291.4]
endmodule
module FringeFF( // @[:@94332.2]
  input         clock, // @[:@94333.4]
  input         reset, // @[:@94334.4]
  input  [63:0] io_in, // @[:@94335.4]
  input         io_reset, // @[:@94335.4]
  output [63:0] io_out, // @[:@94335.4]
  input         io_enable // @[:@94335.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@94338.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@94338.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@94338.4]
  wire [63:0] RetimeWrapper_io_in; // @[package.scala 93:22:@94338.4]
  wire [63:0] RetimeWrapper_io_out; // @[package.scala 93:22:@94338.4]
  wire [63:0] _T_18; // @[package.scala 96:25:@94343.4 package.scala 96:25:@94344.4]
  wire [63:0] _GEN_0; // @[FringeFF.scala 21:27:@94349.6]
  RetimeWrapper_52 RetimeWrapper ( // @[package.scala 93:22:@94338.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@94343.4 package.scala 96:25:@94344.4]
  assign _GEN_0 = io_reset ? 64'h0 : _T_18; // @[FringeFF.scala 21:27:@94349.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@94355.4]
  assign RetimeWrapper_clock = clock; // @[:@94339.4]
  assign RetimeWrapper_reset = reset; // @[:@94340.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@94342.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@94341.4]
endmodule
module MuxN( // @[:@122971.2]
  input  [63:0] io_ins_0, // @[:@122974.4]
  input  [63:0] io_ins_1, // @[:@122974.4]
  input  [63:0] io_ins_2, // @[:@122974.4]
  input  [63:0] io_ins_3, // @[:@122974.4]
  input  [63:0] io_ins_4, // @[:@122974.4]
  input  [63:0] io_ins_5, // @[:@122974.4]
  input  [63:0] io_ins_6, // @[:@122974.4]
  input  [63:0] io_ins_7, // @[:@122974.4]
  input  [63:0] io_ins_8, // @[:@122974.4]
  input  [63:0] io_ins_9, // @[:@122974.4]
  input  [63:0] io_ins_10, // @[:@122974.4]
  input  [63:0] io_ins_11, // @[:@122974.4]
  input  [63:0] io_ins_12, // @[:@122974.4]
  input  [63:0] io_ins_13, // @[:@122974.4]
  input  [63:0] io_ins_14, // @[:@122974.4]
  input  [63:0] io_ins_15, // @[:@122974.4]
  input  [63:0] io_ins_16, // @[:@122974.4]
  input  [63:0] io_ins_17, // @[:@122974.4]
  input  [63:0] io_ins_18, // @[:@122974.4]
  input  [63:0] io_ins_19, // @[:@122974.4]
  input  [63:0] io_ins_20, // @[:@122974.4]
  input  [63:0] io_ins_21, // @[:@122974.4]
  input  [63:0] io_ins_22, // @[:@122974.4]
  input  [63:0] io_ins_23, // @[:@122974.4]
  input  [63:0] io_ins_24, // @[:@122974.4]
  input  [63:0] io_ins_25, // @[:@122974.4]
  input  [63:0] io_ins_26, // @[:@122974.4]
  input  [63:0] io_ins_27, // @[:@122974.4]
  input  [63:0] io_ins_28, // @[:@122974.4]
  input  [63:0] io_ins_29, // @[:@122974.4]
  input  [63:0] io_ins_30, // @[:@122974.4]
  input  [63:0] io_ins_31, // @[:@122974.4]
  input  [63:0] io_ins_32, // @[:@122974.4]
  input  [63:0] io_ins_33, // @[:@122974.4]
  input  [63:0] io_ins_34, // @[:@122974.4]
  input  [63:0] io_ins_35, // @[:@122974.4]
  input  [63:0] io_ins_36, // @[:@122974.4]
  input  [63:0] io_ins_37, // @[:@122974.4]
  input  [63:0] io_ins_38, // @[:@122974.4]
  input  [63:0] io_ins_39, // @[:@122974.4]
  input  [63:0] io_ins_40, // @[:@122974.4]
  input  [63:0] io_ins_41, // @[:@122974.4]
  input  [63:0] io_ins_42, // @[:@122974.4]
  input  [63:0] io_ins_43, // @[:@122974.4]
  input  [63:0] io_ins_44, // @[:@122974.4]
  input  [63:0] io_ins_45, // @[:@122974.4]
  input  [63:0] io_ins_46, // @[:@122974.4]
  input  [63:0] io_ins_47, // @[:@122974.4]
  input  [63:0] io_ins_48, // @[:@122974.4]
  input  [63:0] io_ins_49, // @[:@122974.4]
  input  [63:0] io_ins_50, // @[:@122974.4]
  input  [63:0] io_ins_51, // @[:@122974.4]
  input  [63:0] io_ins_52, // @[:@122974.4]
  input  [63:0] io_ins_53, // @[:@122974.4]
  input  [63:0] io_ins_54, // @[:@122974.4]
  input  [63:0] io_ins_55, // @[:@122974.4]
  input  [63:0] io_ins_56, // @[:@122974.4]
  input  [63:0] io_ins_57, // @[:@122974.4]
  input  [63:0] io_ins_58, // @[:@122974.4]
  input  [63:0] io_ins_59, // @[:@122974.4]
  input  [63:0] io_ins_60, // @[:@122974.4]
  input  [63:0] io_ins_61, // @[:@122974.4]
  input  [63:0] io_ins_62, // @[:@122974.4]
  input  [63:0] io_ins_63, // @[:@122974.4]
  input  [63:0] io_ins_64, // @[:@122974.4]
  input  [63:0] io_ins_65, // @[:@122974.4]
  input  [63:0] io_ins_66, // @[:@122974.4]
  input  [63:0] io_ins_67, // @[:@122974.4]
  input  [63:0] io_ins_68, // @[:@122974.4]
  input  [63:0] io_ins_69, // @[:@122974.4]
  input  [63:0] io_ins_70, // @[:@122974.4]
  input  [63:0] io_ins_71, // @[:@122974.4]
  input  [63:0] io_ins_72, // @[:@122974.4]
  input  [63:0] io_ins_73, // @[:@122974.4]
  input  [63:0] io_ins_74, // @[:@122974.4]
  input  [63:0] io_ins_75, // @[:@122974.4]
  input  [63:0] io_ins_76, // @[:@122974.4]
  input  [63:0] io_ins_77, // @[:@122974.4]
  input  [63:0] io_ins_78, // @[:@122974.4]
  input  [63:0] io_ins_79, // @[:@122974.4]
  input  [63:0] io_ins_80, // @[:@122974.4]
  input  [63:0] io_ins_81, // @[:@122974.4]
  input  [63:0] io_ins_82, // @[:@122974.4]
  input  [63:0] io_ins_83, // @[:@122974.4]
  input  [63:0] io_ins_84, // @[:@122974.4]
  input  [63:0] io_ins_85, // @[:@122974.4]
  input  [63:0] io_ins_86, // @[:@122974.4]
  input  [63:0] io_ins_87, // @[:@122974.4]
  input  [63:0] io_ins_88, // @[:@122974.4]
  input  [63:0] io_ins_89, // @[:@122974.4]
  input  [63:0] io_ins_90, // @[:@122974.4]
  input  [63:0] io_ins_91, // @[:@122974.4]
  input  [63:0] io_ins_92, // @[:@122974.4]
  input  [63:0] io_ins_93, // @[:@122974.4]
  input  [63:0] io_ins_94, // @[:@122974.4]
  input  [63:0] io_ins_95, // @[:@122974.4]
  input  [63:0] io_ins_96, // @[:@122974.4]
  input  [63:0] io_ins_97, // @[:@122974.4]
  input  [63:0] io_ins_98, // @[:@122974.4]
  input  [63:0] io_ins_99, // @[:@122974.4]
  input  [63:0] io_ins_100, // @[:@122974.4]
  input  [63:0] io_ins_101, // @[:@122974.4]
  input  [63:0] io_ins_102, // @[:@122974.4]
  input  [63:0] io_ins_103, // @[:@122974.4]
  input  [63:0] io_ins_104, // @[:@122974.4]
  input  [63:0] io_ins_105, // @[:@122974.4]
  input  [63:0] io_ins_106, // @[:@122974.4]
  input  [63:0] io_ins_107, // @[:@122974.4]
  input  [63:0] io_ins_108, // @[:@122974.4]
  input  [63:0] io_ins_109, // @[:@122974.4]
  input  [63:0] io_ins_110, // @[:@122974.4]
  input  [63:0] io_ins_111, // @[:@122974.4]
  input  [63:0] io_ins_112, // @[:@122974.4]
  input  [63:0] io_ins_113, // @[:@122974.4]
  input  [63:0] io_ins_114, // @[:@122974.4]
  input  [63:0] io_ins_115, // @[:@122974.4]
  input  [63:0] io_ins_116, // @[:@122974.4]
  input  [63:0] io_ins_117, // @[:@122974.4]
  input  [63:0] io_ins_118, // @[:@122974.4]
  input  [63:0] io_ins_119, // @[:@122974.4]
  input  [63:0] io_ins_120, // @[:@122974.4]
  input  [63:0] io_ins_121, // @[:@122974.4]
  input  [63:0] io_ins_122, // @[:@122974.4]
  input  [63:0] io_ins_123, // @[:@122974.4]
  input  [63:0] io_ins_124, // @[:@122974.4]
  input  [63:0] io_ins_125, // @[:@122974.4]
  input  [63:0] io_ins_126, // @[:@122974.4]
  input  [63:0] io_ins_127, // @[:@122974.4]
  input  [63:0] io_ins_128, // @[:@122974.4]
  input  [63:0] io_ins_129, // @[:@122974.4]
  input  [63:0] io_ins_130, // @[:@122974.4]
  input  [63:0] io_ins_131, // @[:@122974.4]
  input  [63:0] io_ins_132, // @[:@122974.4]
  input  [63:0] io_ins_133, // @[:@122974.4]
  input  [63:0] io_ins_134, // @[:@122974.4]
  input  [63:0] io_ins_135, // @[:@122974.4]
  input  [63:0] io_ins_136, // @[:@122974.4]
  input  [63:0] io_ins_137, // @[:@122974.4]
  input  [63:0] io_ins_138, // @[:@122974.4]
  input  [63:0] io_ins_139, // @[:@122974.4]
  input  [63:0] io_ins_140, // @[:@122974.4]
  input  [63:0] io_ins_141, // @[:@122974.4]
  input  [63:0] io_ins_142, // @[:@122974.4]
  input  [63:0] io_ins_143, // @[:@122974.4]
  input  [63:0] io_ins_144, // @[:@122974.4]
  input  [63:0] io_ins_145, // @[:@122974.4]
  input  [63:0] io_ins_146, // @[:@122974.4]
  input  [63:0] io_ins_147, // @[:@122974.4]
  input  [63:0] io_ins_148, // @[:@122974.4]
  input  [63:0] io_ins_149, // @[:@122974.4]
  input  [63:0] io_ins_150, // @[:@122974.4]
  input  [63:0] io_ins_151, // @[:@122974.4]
  input  [63:0] io_ins_152, // @[:@122974.4]
  input  [63:0] io_ins_153, // @[:@122974.4]
  input  [63:0] io_ins_154, // @[:@122974.4]
  input  [63:0] io_ins_155, // @[:@122974.4]
  input  [63:0] io_ins_156, // @[:@122974.4]
  input  [63:0] io_ins_157, // @[:@122974.4]
  input  [63:0] io_ins_158, // @[:@122974.4]
  input  [63:0] io_ins_159, // @[:@122974.4]
  input  [63:0] io_ins_160, // @[:@122974.4]
  input  [63:0] io_ins_161, // @[:@122974.4]
  input  [63:0] io_ins_162, // @[:@122974.4]
  input  [63:0] io_ins_163, // @[:@122974.4]
  input  [63:0] io_ins_164, // @[:@122974.4]
  input  [63:0] io_ins_165, // @[:@122974.4]
  input  [63:0] io_ins_166, // @[:@122974.4]
  input  [63:0] io_ins_167, // @[:@122974.4]
  input  [63:0] io_ins_168, // @[:@122974.4]
  input  [63:0] io_ins_169, // @[:@122974.4]
  input  [63:0] io_ins_170, // @[:@122974.4]
  input  [63:0] io_ins_171, // @[:@122974.4]
  input  [63:0] io_ins_172, // @[:@122974.4]
  input  [63:0] io_ins_173, // @[:@122974.4]
  input  [63:0] io_ins_174, // @[:@122974.4]
  input  [63:0] io_ins_175, // @[:@122974.4]
  input  [63:0] io_ins_176, // @[:@122974.4]
  input  [63:0] io_ins_177, // @[:@122974.4]
  input  [63:0] io_ins_178, // @[:@122974.4]
  input  [63:0] io_ins_179, // @[:@122974.4]
  input  [63:0] io_ins_180, // @[:@122974.4]
  input  [63:0] io_ins_181, // @[:@122974.4]
  input  [63:0] io_ins_182, // @[:@122974.4]
  input  [63:0] io_ins_183, // @[:@122974.4]
  input  [63:0] io_ins_184, // @[:@122974.4]
  input  [63:0] io_ins_185, // @[:@122974.4]
  input  [63:0] io_ins_186, // @[:@122974.4]
  input  [63:0] io_ins_187, // @[:@122974.4]
  input  [63:0] io_ins_188, // @[:@122974.4]
  input  [63:0] io_ins_189, // @[:@122974.4]
  input  [63:0] io_ins_190, // @[:@122974.4]
  input  [63:0] io_ins_191, // @[:@122974.4]
  input  [63:0] io_ins_192, // @[:@122974.4]
  input  [63:0] io_ins_193, // @[:@122974.4]
  input  [63:0] io_ins_194, // @[:@122974.4]
  input  [63:0] io_ins_195, // @[:@122974.4]
  input  [63:0] io_ins_196, // @[:@122974.4]
  input  [63:0] io_ins_197, // @[:@122974.4]
  input  [63:0] io_ins_198, // @[:@122974.4]
  input  [63:0] io_ins_199, // @[:@122974.4]
  input  [63:0] io_ins_200, // @[:@122974.4]
  input  [63:0] io_ins_201, // @[:@122974.4]
  input  [63:0] io_ins_202, // @[:@122974.4]
  input  [63:0] io_ins_203, // @[:@122974.4]
  input  [63:0] io_ins_204, // @[:@122974.4]
  input  [63:0] io_ins_205, // @[:@122974.4]
  input  [63:0] io_ins_206, // @[:@122974.4]
  input  [63:0] io_ins_207, // @[:@122974.4]
  input  [63:0] io_ins_208, // @[:@122974.4]
  input  [63:0] io_ins_209, // @[:@122974.4]
  input  [63:0] io_ins_210, // @[:@122974.4]
  input  [63:0] io_ins_211, // @[:@122974.4]
  input  [63:0] io_ins_212, // @[:@122974.4]
  input  [63:0] io_ins_213, // @[:@122974.4]
  input  [63:0] io_ins_214, // @[:@122974.4]
  input  [63:0] io_ins_215, // @[:@122974.4]
  input  [63:0] io_ins_216, // @[:@122974.4]
  input  [63:0] io_ins_217, // @[:@122974.4]
  input  [63:0] io_ins_218, // @[:@122974.4]
  input  [63:0] io_ins_219, // @[:@122974.4]
  input  [63:0] io_ins_220, // @[:@122974.4]
  input  [63:0] io_ins_221, // @[:@122974.4]
  input  [63:0] io_ins_222, // @[:@122974.4]
  input  [63:0] io_ins_223, // @[:@122974.4]
  input  [63:0] io_ins_224, // @[:@122974.4]
  input  [63:0] io_ins_225, // @[:@122974.4]
  input  [63:0] io_ins_226, // @[:@122974.4]
  input  [63:0] io_ins_227, // @[:@122974.4]
  input  [63:0] io_ins_228, // @[:@122974.4]
  input  [63:0] io_ins_229, // @[:@122974.4]
  input  [63:0] io_ins_230, // @[:@122974.4]
  input  [63:0] io_ins_231, // @[:@122974.4]
  input  [63:0] io_ins_232, // @[:@122974.4]
  input  [63:0] io_ins_233, // @[:@122974.4]
  input  [63:0] io_ins_234, // @[:@122974.4]
  input  [63:0] io_ins_235, // @[:@122974.4]
  input  [63:0] io_ins_236, // @[:@122974.4]
  input  [63:0] io_ins_237, // @[:@122974.4]
  input  [63:0] io_ins_238, // @[:@122974.4]
  input  [63:0] io_ins_239, // @[:@122974.4]
  input  [63:0] io_ins_240, // @[:@122974.4]
  input  [63:0] io_ins_241, // @[:@122974.4]
  input  [63:0] io_ins_242, // @[:@122974.4]
  input  [63:0] io_ins_243, // @[:@122974.4]
  input  [63:0] io_ins_244, // @[:@122974.4]
  input  [63:0] io_ins_245, // @[:@122974.4]
  input  [63:0] io_ins_246, // @[:@122974.4]
  input  [63:0] io_ins_247, // @[:@122974.4]
  input  [63:0] io_ins_248, // @[:@122974.4]
  input  [63:0] io_ins_249, // @[:@122974.4]
  input  [63:0] io_ins_250, // @[:@122974.4]
  input  [63:0] io_ins_251, // @[:@122974.4]
  input  [63:0] io_ins_252, // @[:@122974.4]
  input  [63:0] io_ins_253, // @[:@122974.4]
  input  [63:0] io_ins_254, // @[:@122974.4]
  input  [63:0] io_ins_255, // @[:@122974.4]
  input  [63:0] io_ins_256, // @[:@122974.4]
  input  [63:0] io_ins_257, // @[:@122974.4]
  input  [63:0] io_ins_258, // @[:@122974.4]
  input  [63:0] io_ins_259, // @[:@122974.4]
  input  [63:0] io_ins_260, // @[:@122974.4]
  input  [63:0] io_ins_261, // @[:@122974.4]
  input  [63:0] io_ins_262, // @[:@122974.4]
  input  [63:0] io_ins_263, // @[:@122974.4]
  input  [63:0] io_ins_264, // @[:@122974.4]
  input  [63:0] io_ins_265, // @[:@122974.4]
  input  [63:0] io_ins_266, // @[:@122974.4]
  input  [63:0] io_ins_267, // @[:@122974.4]
  input  [63:0] io_ins_268, // @[:@122974.4]
  input  [63:0] io_ins_269, // @[:@122974.4]
  input  [63:0] io_ins_270, // @[:@122974.4]
  input  [63:0] io_ins_271, // @[:@122974.4]
  input  [63:0] io_ins_272, // @[:@122974.4]
  input  [63:0] io_ins_273, // @[:@122974.4]
  input  [63:0] io_ins_274, // @[:@122974.4]
  input  [63:0] io_ins_275, // @[:@122974.4]
  input  [63:0] io_ins_276, // @[:@122974.4]
  input  [63:0] io_ins_277, // @[:@122974.4]
  input  [63:0] io_ins_278, // @[:@122974.4]
  input  [63:0] io_ins_279, // @[:@122974.4]
  input  [63:0] io_ins_280, // @[:@122974.4]
  input  [63:0] io_ins_281, // @[:@122974.4]
  input  [63:0] io_ins_282, // @[:@122974.4]
  input  [63:0] io_ins_283, // @[:@122974.4]
  input  [63:0] io_ins_284, // @[:@122974.4]
  input  [63:0] io_ins_285, // @[:@122974.4]
  input  [63:0] io_ins_286, // @[:@122974.4]
  input  [63:0] io_ins_287, // @[:@122974.4]
  input  [63:0] io_ins_288, // @[:@122974.4]
  input  [63:0] io_ins_289, // @[:@122974.4]
  input  [63:0] io_ins_290, // @[:@122974.4]
  input  [63:0] io_ins_291, // @[:@122974.4]
  input  [63:0] io_ins_292, // @[:@122974.4]
  input  [63:0] io_ins_293, // @[:@122974.4]
  input  [63:0] io_ins_294, // @[:@122974.4]
  input  [63:0] io_ins_295, // @[:@122974.4]
  input  [63:0] io_ins_296, // @[:@122974.4]
  input  [63:0] io_ins_297, // @[:@122974.4]
  input  [63:0] io_ins_298, // @[:@122974.4]
  input  [63:0] io_ins_299, // @[:@122974.4]
  input  [63:0] io_ins_300, // @[:@122974.4]
  input  [63:0] io_ins_301, // @[:@122974.4]
  input  [63:0] io_ins_302, // @[:@122974.4]
  input  [63:0] io_ins_303, // @[:@122974.4]
  input  [63:0] io_ins_304, // @[:@122974.4]
  input  [63:0] io_ins_305, // @[:@122974.4]
  input  [63:0] io_ins_306, // @[:@122974.4]
  input  [63:0] io_ins_307, // @[:@122974.4]
  input  [63:0] io_ins_308, // @[:@122974.4]
  input  [63:0] io_ins_309, // @[:@122974.4]
  input  [63:0] io_ins_310, // @[:@122974.4]
  input  [63:0] io_ins_311, // @[:@122974.4]
  input  [63:0] io_ins_312, // @[:@122974.4]
  input  [63:0] io_ins_313, // @[:@122974.4]
  input  [63:0] io_ins_314, // @[:@122974.4]
  input  [63:0] io_ins_315, // @[:@122974.4]
  input  [63:0] io_ins_316, // @[:@122974.4]
  input  [63:0] io_ins_317, // @[:@122974.4]
  input  [63:0] io_ins_318, // @[:@122974.4]
  input  [63:0] io_ins_319, // @[:@122974.4]
  input  [63:0] io_ins_320, // @[:@122974.4]
  input  [63:0] io_ins_321, // @[:@122974.4]
  input  [63:0] io_ins_322, // @[:@122974.4]
  input  [63:0] io_ins_323, // @[:@122974.4]
  input  [63:0] io_ins_324, // @[:@122974.4]
  input  [63:0] io_ins_325, // @[:@122974.4]
  input  [63:0] io_ins_326, // @[:@122974.4]
  input  [63:0] io_ins_327, // @[:@122974.4]
  input  [63:0] io_ins_328, // @[:@122974.4]
  input  [63:0] io_ins_329, // @[:@122974.4]
  input  [63:0] io_ins_330, // @[:@122974.4]
  input  [63:0] io_ins_331, // @[:@122974.4]
  input  [63:0] io_ins_332, // @[:@122974.4]
  input  [63:0] io_ins_333, // @[:@122974.4]
  input  [63:0] io_ins_334, // @[:@122974.4]
  input  [63:0] io_ins_335, // @[:@122974.4]
  input  [63:0] io_ins_336, // @[:@122974.4]
  input  [63:0] io_ins_337, // @[:@122974.4]
  input  [63:0] io_ins_338, // @[:@122974.4]
  input  [63:0] io_ins_339, // @[:@122974.4]
  input  [63:0] io_ins_340, // @[:@122974.4]
  input  [63:0] io_ins_341, // @[:@122974.4]
  input  [63:0] io_ins_342, // @[:@122974.4]
  input  [63:0] io_ins_343, // @[:@122974.4]
  input  [63:0] io_ins_344, // @[:@122974.4]
  input  [63:0] io_ins_345, // @[:@122974.4]
  input  [63:0] io_ins_346, // @[:@122974.4]
  input  [63:0] io_ins_347, // @[:@122974.4]
  input  [63:0] io_ins_348, // @[:@122974.4]
  input  [63:0] io_ins_349, // @[:@122974.4]
  input  [63:0] io_ins_350, // @[:@122974.4]
  input  [63:0] io_ins_351, // @[:@122974.4]
  input  [63:0] io_ins_352, // @[:@122974.4]
  input  [63:0] io_ins_353, // @[:@122974.4]
  input  [63:0] io_ins_354, // @[:@122974.4]
  input  [63:0] io_ins_355, // @[:@122974.4]
  input  [63:0] io_ins_356, // @[:@122974.4]
  input  [63:0] io_ins_357, // @[:@122974.4]
  input  [63:0] io_ins_358, // @[:@122974.4]
  input  [63:0] io_ins_359, // @[:@122974.4]
  input  [63:0] io_ins_360, // @[:@122974.4]
  input  [63:0] io_ins_361, // @[:@122974.4]
  input  [63:0] io_ins_362, // @[:@122974.4]
  input  [63:0] io_ins_363, // @[:@122974.4]
  input  [63:0] io_ins_364, // @[:@122974.4]
  input  [63:0] io_ins_365, // @[:@122974.4]
  input  [63:0] io_ins_366, // @[:@122974.4]
  input  [63:0] io_ins_367, // @[:@122974.4]
  input  [63:0] io_ins_368, // @[:@122974.4]
  input  [63:0] io_ins_369, // @[:@122974.4]
  input  [63:0] io_ins_370, // @[:@122974.4]
  input  [63:0] io_ins_371, // @[:@122974.4]
  input  [63:0] io_ins_372, // @[:@122974.4]
  input  [63:0] io_ins_373, // @[:@122974.4]
  input  [63:0] io_ins_374, // @[:@122974.4]
  input  [63:0] io_ins_375, // @[:@122974.4]
  input  [63:0] io_ins_376, // @[:@122974.4]
  input  [63:0] io_ins_377, // @[:@122974.4]
  input  [63:0] io_ins_378, // @[:@122974.4]
  input  [63:0] io_ins_379, // @[:@122974.4]
  input  [63:0] io_ins_380, // @[:@122974.4]
  input  [63:0] io_ins_381, // @[:@122974.4]
  input  [63:0] io_ins_382, // @[:@122974.4]
  input  [63:0] io_ins_383, // @[:@122974.4]
  input  [63:0] io_ins_384, // @[:@122974.4]
  input  [63:0] io_ins_385, // @[:@122974.4]
  input  [63:0] io_ins_386, // @[:@122974.4]
  input  [63:0] io_ins_387, // @[:@122974.4]
  input  [63:0] io_ins_388, // @[:@122974.4]
  input  [63:0] io_ins_389, // @[:@122974.4]
  input  [63:0] io_ins_390, // @[:@122974.4]
  input  [63:0] io_ins_391, // @[:@122974.4]
  input  [63:0] io_ins_392, // @[:@122974.4]
  input  [63:0] io_ins_393, // @[:@122974.4]
  input  [63:0] io_ins_394, // @[:@122974.4]
  input  [63:0] io_ins_395, // @[:@122974.4]
  input  [63:0] io_ins_396, // @[:@122974.4]
  input  [63:0] io_ins_397, // @[:@122974.4]
  input  [63:0] io_ins_398, // @[:@122974.4]
  input  [63:0] io_ins_399, // @[:@122974.4]
  input  [63:0] io_ins_400, // @[:@122974.4]
  input  [63:0] io_ins_401, // @[:@122974.4]
  input  [63:0] io_ins_402, // @[:@122974.4]
  input  [63:0] io_ins_403, // @[:@122974.4]
  input  [63:0] io_ins_404, // @[:@122974.4]
  input  [63:0] io_ins_405, // @[:@122974.4]
  input  [63:0] io_ins_406, // @[:@122974.4]
  input  [63:0] io_ins_407, // @[:@122974.4]
  input  [63:0] io_ins_408, // @[:@122974.4]
  input  [63:0] io_ins_409, // @[:@122974.4]
  input  [63:0] io_ins_410, // @[:@122974.4]
  input  [63:0] io_ins_411, // @[:@122974.4]
  input  [63:0] io_ins_412, // @[:@122974.4]
  input  [63:0] io_ins_413, // @[:@122974.4]
  input  [63:0] io_ins_414, // @[:@122974.4]
  input  [63:0] io_ins_415, // @[:@122974.4]
  input  [63:0] io_ins_416, // @[:@122974.4]
  input  [63:0] io_ins_417, // @[:@122974.4]
  input  [63:0] io_ins_418, // @[:@122974.4]
  input  [63:0] io_ins_419, // @[:@122974.4]
  input  [63:0] io_ins_420, // @[:@122974.4]
  input  [63:0] io_ins_421, // @[:@122974.4]
  input  [63:0] io_ins_422, // @[:@122974.4]
  input  [63:0] io_ins_423, // @[:@122974.4]
  input  [63:0] io_ins_424, // @[:@122974.4]
  input  [63:0] io_ins_425, // @[:@122974.4]
  input  [63:0] io_ins_426, // @[:@122974.4]
  input  [63:0] io_ins_427, // @[:@122974.4]
  input  [63:0] io_ins_428, // @[:@122974.4]
  input  [63:0] io_ins_429, // @[:@122974.4]
  input  [63:0] io_ins_430, // @[:@122974.4]
  input  [63:0] io_ins_431, // @[:@122974.4]
  input  [63:0] io_ins_432, // @[:@122974.4]
  input  [63:0] io_ins_433, // @[:@122974.4]
  input  [63:0] io_ins_434, // @[:@122974.4]
  input  [63:0] io_ins_435, // @[:@122974.4]
  input  [63:0] io_ins_436, // @[:@122974.4]
  input  [63:0] io_ins_437, // @[:@122974.4]
  input  [63:0] io_ins_438, // @[:@122974.4]
  input  [63:0] io_ins_439, // @[:@122974.4]
  input  [63:0] io_ins_440, // @[:@122974.4]
  input  [63:0] io_ins_441, // @[:@122974.4]
  input  [63:0] io_ins_442, // @[:@122974.4]
  input  [63:0] io_ins_443, // @[:@122974.4]
  input  [63:0] io_ins_444, // @[:@122974.4]
  input  [63:0] io_ins_445, // @[:@122974.4]
  input  [63:0] io_ins_446, // @[:@122974.4]
  input  [63:0] io_ins_447, // @[:@122974.4]
  input  [63:0] io_ins_448, // @[:@122974.4]
  input  [63:0] io_ins_449, // @[:@122974.4]
  input  [63:0] io_ins_450, // @[:@122974.4]
  input  [63:0] io_ins_451, // @[:@122974.4]
  input  [63:0] io_ins_452, // @[:@122974.4]
  input  [63:0] io_ins_453, // @[:@122974.4]
  input  [63:0] io_ins_454, // @[:@122974.4]
  input  [63:0] io_ins_455, // @[:@122974.4]
  input  [63:0] io_ins_456, // @[:@122974.4]
  input  [63:0] io_ins_457, // @[:@122974.4]
  input  [63:0] io_ins_458, // @[:@122974.4]
  input  [63:0] io_ins_459, // @[:@122974.4]
  input  [63:0] io_ins_460, // @[:@122974.4]
  input  [63:0] io_ins_461, // @[:@122974.4]
  input  [63:0] io_ins_462, // @[:@122974.4]
  input  [63:0] io_ins_463, // @[:@122974.4]
  input  [63:0] io_ins_464, // @[:@122974.4]
  input  [63:0] io_ins_465, // @[:@122974.4]
  input  [63:0] io_ins_466, // @[:@122974.4]
  input  [63:0] io_ins_467, // @[:@122974.4]
  input  [63:0] io_ins_468, // @[:@122974.4]
  input  [63:0] io_ins_469, // @[:@122974.4]
  input  [63:0] io_ins_470, // @[:@122974.4]
  input  [63:0] io_ins_471, // @[:@122974.4]
  input  [63:0] io_ins_472, // @[:@122974.4]
  input  [63:0] io_ins_473, // @[:@122974.4]
  input  [63:0] io_ins_474, // @[:@122974.4]
  input  [63:0] io_ins_475, // @[:@122974.4]
  input  [63:0] io_ins_476, // @[:@122974.4]
  input  [63:0] io_ins_477, // @[:@122974.4]
  input  [63:0] io_ins_478, // @[:@122974.4]
  input  [63:0] io_ins_479, // @[:@122974.4]
  input  [63:0] io_ins_480, // @[:@122974.4]
  input  [63:0] io_ins_481, // @[:@122974.4]
  input  [63:0] io_ins_482, // @[:@122974.4]
  input  [63:0] io_ins_483, // @[:@122974.4]
  input  [63:0] io_ins_484, // @[:@122974.4]
  input  [63:0] io_ins_485, // @[:@122974.4]
  input  [63:0] io_ins_486, // @[:@122974.4]
  input  [63:0] io_ins_487, // @[:@122974.4]
  input  [63:0] io_ins_488, // @[:@122974.4]
  input  [63:0] io_ins_489, // @[:@122974.4]
  input  [63:0] io_ins_490, // @[:@122974.4]
  input  [63:0] io_ins_491, // @[:@122974.4]
  input  [63:0] io_ins_492, // @[:@122974.4]
  input  [63:0] io_ins_493, // @[:@122974.4]
  input  [63:0] io_ins_494, // @[:@122974.4]
  input  [63:0] io_ins_495, // @[:@122974.4]
  input  [63:0] io_ins_496, // @[:@122974.4]
  input  [63:0] io_ins_497, // @[:@122974.4]
  input  [63:0] io_ins_498, // @[:@122974.4]
  input  [63:0] io_ins_499, // @[:@122974.4]
  input  [63:0] io_ins_500, // @[:@122974.4]
  input  [63:0] io_ins_501, // @[:@122974.4]
  input  [63:0] io_ins_502, // @[:@122974.4]
  input  [8:0]  io_sel, // @[:@122974.4]
  output [63:0] io_out // @[:@122974.4]
);
  wire [63:0] _GEN_1; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_2; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_3; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_4; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_5; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_6; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_7; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_8; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_9; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_10; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_11; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_12; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_13; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_14; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_15; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_16; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_17; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_18; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_19; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_20; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_21; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_22; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_23; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_24; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_25; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_26; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_27; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_28; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_29; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_30; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_31; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_32; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_33; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_34; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_35; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_36; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_37; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_38; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_39; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_40; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_41; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_42; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_43; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_44; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_45; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_46; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_47; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_48; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_49; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_50; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_51; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_52; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_53; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_54; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_55; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_56; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_57; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_58; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_59; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_60; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_61; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_62; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_63; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_64; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_65; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_66; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_67; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_68; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_69; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_70; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_71; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_72; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_73; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_74; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_75; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_76; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_77; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_78; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_79; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_80; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_81; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_82; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_83; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_84; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_85; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_86; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_87; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_88; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_89; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_90; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_91; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_92; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_93; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_94; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_95; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_96; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_97; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_98; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_99; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_100; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_101; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_102; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_103; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_104; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_105; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_106; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_107; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_108; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_109; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_110; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_111; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_112; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_113; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_114; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_115; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_116; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_117; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_118; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_119; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_120; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_121; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_122; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_123; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_124; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_125; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_126; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_127; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_128; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_129; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_130; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_131; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_132; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_133; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_134; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_135; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_136; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_137; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_138; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_139; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_140; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_141; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_142; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_143; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_144; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_145; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_146; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_147; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_148; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_149; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_150; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_151; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_152; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_153; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_154; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_155; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_156; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_157; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_158; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_159; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_160; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_161; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_162; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_163; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_164; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_165; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_166; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_167; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_168; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_169; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_170; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_171; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_172; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_173; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_174; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_175; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_176; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_177; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_178; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_179; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_180; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_181; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_182; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_183; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_184; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_185; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_186; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_187; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_188; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_189; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_190; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_191; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_192; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_193; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_194; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_195; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_196; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_197; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_198; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_199; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_200; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_201; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_202; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_203; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_204; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_205; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_206; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_207; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_208; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_209; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_210; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_211; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_212; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_213; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_214; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_215; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_216; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_217; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_218; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_219; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_220; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_221; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_222; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_223; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_224; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_225; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_226; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_227; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_228; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_229; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_230; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_231; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_232; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_233; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_234; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_235; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_236; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_237; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_238; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_239; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_240; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_241; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_242; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_243; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_244; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_245; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_246; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_247; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_248; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_249; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_250; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_251; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_252; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_253; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_254; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_255; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_256; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_257; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_258; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_259; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_260; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_261; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_262; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_263; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_264; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_265; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_266; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_267; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_268; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_269; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_270; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_271; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_272; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_273; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_274; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_275; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_276; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_277; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_278; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_279; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_280; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_281; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_282; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_283; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_284; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_285; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_286; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_287; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_288; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_289; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_290; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_291; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_292; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_293; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_294; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_295; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_296; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_297; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_298; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_299; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_300; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_301; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_302; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_303; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_304; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_305; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_306; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_307; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_308; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_309; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_310; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_311; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_312; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_313; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_314; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_315; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_316; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_317; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_318; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_319; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_320; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_321; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_322; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_323; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_324; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_325; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_326; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_327; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_328; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_329; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_330; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_331; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_332; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_333; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_334; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_335; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_336; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_337; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_338; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_339; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_340; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_341; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_342; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_343; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_344; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_345; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_346; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_347; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_348; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_349; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_350; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_351; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_352; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_353; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_354; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_355; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_356; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_357; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_358; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_359; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_360; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_361; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_362; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_363; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_364; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_365; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_366; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_367; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_368; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_369; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_370; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_371; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_372; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_373; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_374; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_375; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_376; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_377; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_378; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_379; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_380; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_381; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_382; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_383; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_384; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_385; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_386; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_387; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_388; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_389; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_390; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_391; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_392; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_393; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_394; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_395; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_396; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_397; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_398; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_399; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_400; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_401; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_402; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_403; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_404; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_405; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_406; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_407; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_408; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_409; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_410; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_411; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_412; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_413; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_414; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_415; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_416; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_417; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_418; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_419; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_420; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_421; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_422; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_423; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_424; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_425; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_426; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_427; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_428; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_429; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_430; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_431; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_432; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_433; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_434; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_435; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_436; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_437; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_438; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_439; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_440; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_441; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_442; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_443; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_444; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_445; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_446; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_447; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_448; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_449; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_450; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_451; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_452; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_453; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_454; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_455; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_456; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_457; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_458; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_459; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_460; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_461; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_462; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_463; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_464; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_465; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_466; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_467; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_468; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_469; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_470; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_471; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_472; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_473; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_474; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_475; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_476; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_477; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_478; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_479; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_480; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_481; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_482; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_483; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_484; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_485; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_486; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_487; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_488; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_489; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_490; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_491; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_492; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_493; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_494; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_495; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_496; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_497; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_498; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_499; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_500; // @[MuxN.scala 16:10:@122976.4]
  wire [63:0] _GEN_501; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_1 = 9'h1 == io_sel ? io_ins_1 : io_ins_0; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_2 = 9'h2 == io_sel ? io_ins_2 : _GEN_1; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_3 = 9'h3 == io_sel ? io_ins_3 : _GEN_2; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_4 = 9'h4 == io_sel ? io_ins_4 : _GEN_3; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_5 = 9'h5 == io_sel ? io_ins_5 : _GEN_4; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_6 = 9'h6 == io_sel ? io_ins_6 : _GEN_5; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_7 = 9'h7 == io_sel ? io_ins_7 : _GEN_6; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_8 = 9'h8 == io_sel ? io_ins_8 : _GEN_7; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_9 = 9'h9 == io_sel ? io_ins_9 : _GEN_8; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_10 = 9'ha == io_sel ? io_ins_10 : _GEN_9; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_11 = 9'hb == io_sel ? io_ins_11 : _GEN_10; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_12 = 9'hc == io_sel ? io_ins_12 : _GEN_11; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_13 = 9'hd == io_sel ? io_ins_13 : _GEN_12; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_14 = 9'he == io_sel ? io_ins_14 : _GEN_13; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_15 = 9'hf == io_sel ? io_ins_15 : _GEN_14; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_16 = 9'h10 == io_sel ? io_ins_16 : _GEN_15; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_17 = 9'h11 == io_sel ? io_ins_17 : _GEN_16; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_18 = 9'h12 == io_sel ? io_ins_18 : _GEN_17; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_19 = 9'h13 == io_sel ? io_ins_19 : _GEN_18; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_20 = 9'h14 == io_sel ? io_ins_20 : _GEN_19; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_21 = 9'h15 == io_sel ? io_ins_21 : _GEN_20; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_22 = 9'h16 == io_sel ? io_ins_22 : _GEN_21; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_23 = 9'h17 == io_sel ? io_ins_23 : _GEN_22; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_24 = 9'h18 == io_sel ? io_ins_24 : _GEN_23; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_25 = 9'h19 == io_sel ? io_ins_25 : _GEN_24; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_26 = 9'h1a == io_sel ? io_ins_26 : _GEN_25; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_27 = 9'h1b == io_sel ? io_ins_27 : _GEN_26; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_28 = 9'h1c == io_sel ? io_ins_28 : _GEN_27; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_29 = 9'h1d == io_sel ? io_ins_29 : _GEN_28; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_30 = 9'h1e == io_sel ? io_ins_30 : _GEN_29; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_31 = 9'h1f == io_sel ? io_ins_31 : _GEN_30; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_32 = 9'h20 == io_sel ? io_ins_32 : _GEN_31; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_33 = 9'h21 == io_sel ? io_ins_33 : _GEN_32; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_34 = 9'h22 == io_sel ? io_ins_34 : _GEN_33; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_35 = 9'h23 == io_sel ? io_ins_35 : _GEN_34; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_36 = 9'h24 == io_sel ? io_ins_36 : _GEN_35; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_37 = 9'h25 == io_sel ? io_ins_37 : _GEN_36; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_38 = 9'h26 == io_sel ? io_ins_38 : _GEN_37; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_39 = 9'h27 == io_sel ? io_ins_39 : _GEN_38; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_40 = 9'h28 == io_sel ? io_ins_40 : _GEN_39; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_41 = 9'h29 == io_sel ? io_ins_41 : _GEN_40; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_42 = 9'h2a == io_sel ? io_ins_42 : _GEN_41; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_43 = 9'h2b == io_sel ? io_ins_43 : _GEN_42; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_44 = 9'h2c == io_sel ? io_ins_44 : _GEN_43; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_45 = 9'h2d == io_sel ? io_ins_45 : _GEN_44; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_46 = 9'h2e == io_sel ? io_ins_46 : _GEN_45; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_47 = 9'h2f == io_sel ? io_ins_47 : _GEN_46; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_48 = 9'h30 == io_sel ? io_ins_48 : _GEN_47; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_49 = 9'h31 == io_sel ? io_ins_49 : _GEN_48; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_50 = 9'h32 == io_sel ? io_ins_50 : _GEN_49; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_51 = 9'h33 == io_sel ? io_ins_51 : _GEN_50; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_52 = 9'h34 == io_sel ? io_ins_52 : _GEN_51; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_53 = 9'h35 == io_sel ? io_ins_53 : _GEN_52; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_54 = 9'h36 == io_sel ? io_ins_54 : _GEN_53; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_55 = 9'h37 == io_sel ? io_ins_55 : _GEN_54; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_56 = 9'h38 == io_sel ? io_ins_56 : _GEN_55; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_57 = 9'h39 == io_sel ? io_ins_57 : _GEN_56; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_58 = 9'h3a == io_sel ? io_ins_58 : _GEN_57; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_59 = 9'h3b == io_sel ? io_ins_59 : _GEN_58; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_60 = 9'h3c == io_sel ? io_ins_60 : _GEN_59; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_61 = 9'h3d == io_sel ? io_ins_61 : _GEN_60; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_62 = 9'h3e == io_sel ? io_ins_62 : _GEN_61; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_63 = 9'h3f == io_sel ? io_ins_63 : _GEN_62; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_64 = 9'h40 == io_sel ? io_ins_64 : _GEN_63; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_65 = 9'h41 == io_sel ? io_ins_65 : _GEN_64; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_66 = 9'h42 == io_sel ? io_ins_66 : _GEN_65; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_67 = 9'h43 == io_sel ? io_ins_67 : _GEN_66; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_68 = 9'h44 == io_sel ? io_ins_68 : _GEN_67; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_69 = 9'h45 == io_sel ? io_ins_69 : _GEN_68; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_70 = 9'h46 == io_sel ? io_ins_70 : _GEN_69; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_71 = 9'h47 == io_sel ? io_ins_71 : _GEN_70; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_72 = 9'h48 == io_sel ? io_ins_72 : _GEN_71; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_73 = 9'h49 == io_sel ? io_ins_73 : _GEN_72; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_74 = 9'h4a == io_sel ? io_ins_74 : _GEN_73; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_75 = 9'h4b == io_sel ? io_ins_75 : _GEN_74; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_76 = 9'h4c == io_sel ? io_ins_76 : _GEN_75; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_77 = 9'h4d == io_sel ? io_ins_77 : _GEN_76; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_78 = 9'h4e == io_sel ? io_ins_78 : _GEN_77; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_79 = 9'h4f == io_sel ? io_ins_79 : _GEN_78; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_80 = 9'h50 == io_sel ? io_ins_80 : _GEN_79; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_81 = 9'h51 == io_sel ? io_ins_81 : _GEN_80; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_82 = 9'h52 == io_sel ? io_ins_82 : _GEN_81; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_83 = 9'h53 == io_sel ? io_ins_83 : _GEN_82; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_84 = 9'h54 == io_sel ? io_ins_84 : _GEN_83; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_85 = 9'h55 == io_sel ? io_ins_85 : _GEN_84; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_86 = 9'h56 == io_sel ? io_ins_86 : _GEN_85; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_87 = 9'h57 == io_sel ? io_ins_87 : _GEN_86; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_88 = 9'h58 == io_sel ? io_ins_88 : _GEN_87; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_89 = 9'h59 == io_sel ? io_ins_89 : _GEN_88; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_90 = 9'h5a == io_sel ? io_ins_90 : _GEN_89; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_91 = 9'h5b == io_sel ? io_ins_91 : _GEN_90; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_92 = 9'h5c == io_sel ? io_ins_92 : _GEN_91; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_93 = 9'h5d == io_sel ? io_ins_93 : _GEN_92; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_94 = 9'h5e == io_sel ? io_ins_94 : _GEN_93; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_95 = 9'h5f == io_sel ? io_ins_95 : _GEN_94; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_96 = 9'h60 == io_sel ? io_ins_96 : _GEN_95; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_97 = 9'h61 == io_sel ? io_ins_97 : _GEN_96; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_98 = 9'h62 == io_sel ? io_ins_98 : _GEN_97; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_99 = 9'h63 == io_sel ? io_ins_99 : _GEN_98; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_100 = 9'h64 == io_sel ? io_ins_100 : _GEN_99; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_101 = 9'h65 == io_sel ? io_ins_101 : _GEN_100; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_102 = 9'h66 == io_sel ? io_ins_102 : _GEN_101; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_103 = 9'h67 == io_sel ? io_ins_103 : _GEN_102; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_104 = 9'h68 == io_sel ? io_ins_104 : _GEN_103; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_105 = 9'h69 == io_sel ? io_ins_105 : _GEN_104; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_106 = 9'h6a == io_sel ? io_ins_106 : _GEN_105; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_107 = 9'h6b == io_sel ? io_ins_107 : _GEN_106; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_108 = 9'h6c == io_sel ? io_ins_108 : _GEN_107; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_109 = 9'h6d == io_sel ? io_ins_109 : _GEN_108; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_110 = 9'h6e == io_sel ? io_ins_110 : _GEN_109; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_111 = 9'h6f == io_sel ? io_ins_111 : _GEN_110; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_112 = 9'h70 == io_sel ? io_ins_112 : _GEN_111; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_113 = 9'h71 == io_sel ? io_ins_113 : _GEN_112; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_114 = 9'h72 == io_sel ? io_ins_114 : _GEN_113; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_115 = 9'h73 == io_sel ? io_ins_115 : _GEN_114; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_116 = 9'h74 == io_sel ? io_ins_116 : _GEN_115; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_117 = 9'h75 == io_sel ? io_ins_117 : _GEN_116; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_118 = 9'h76 == io_sel ? io_ins_118 : _GEN_117; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_119 = 9'h77 == io_sel ? io_ins_119 : _GEN_118; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_120 = 9'h78 == io_sel ? io_ins_120 : _GEN_119; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_121 = 9'h79 == io_sel ? io_ins_121 : _GEN_120; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_122 = 9'h7a == io_sel ? io_ins_122 : _GEN_121; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_123 = 9'h7b == io_sel ? io_ins_123 : _GEN_122; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_124 = 9'h7c == io_sel ? io_ins_124 : _GEN_123; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_125 = 9'h7d == io_sel ? io_ins_125 : _GEN_124; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_126 = 9'h7e == io_sel ? io_ins_126 : _GEN_125; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_127 = 9'h7f == io_sel ? io_ins_127 : _GEN_126; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_128 = 9'h80 == io_sel ? io_ins_128 : _GEN_127; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_129 = 9'h81 == io_sel ? io_ins_129 : _GEN_128; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_130 = 9'h82 == io_sel ? io_ins_130 : _GEN_129; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_131 = 9'h83 == io_sel ? io_ins_131 : _GEN_130; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_132 = 9'h84 == io_sel ? io_ins_132 : _GEN_131; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_133 = 9'h85 == io_sel ? io_ins_133 : _GEN_132; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_134 = 9'h86 == io_sel ? io_ins_134 : _GEN_133; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_135 = 9'h87 == io_sel ? io_ins_135 : _GEN_134; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_136 = 9'h88 == io_sel ? io_ins_136 : _GEN_135; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_137 = 9'h89 == io_sel ? io_ins_137 : _GEN_136; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_138 = 9'h8a == io_sel ? io_ins_138 : _GEN_137; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_139 = 9'h8b == io_sel ? io_ins_139 : _GEN_138; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_140 = 9'h8c == io_sel ? io_ins_140 : _GEN_139; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_141 = 9'h8d == io_sel ? io_ins_141 : _GEN_140; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_142 = 9'h8e == io_sel ? io_ins_142 : _GEN_141; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_143 = 9'h8f == io_sel ? io_ins_143 : _GEN_142; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_144 = 9'h90 == io_sel ? io_ins_144 : _GEN_143; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_145 = 9'h91 == io_sel ? io_ins_145 : _GEN_144; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_146 = 9'h92 == io_sel ? io_ins_146 : _GEN_145; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_147 = 9'h93 == io_sel ? io_ins_147 : _GEN_146; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_148 = 9'h94 == io_sel ? io_ins_148 : _GEN_147; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_149 = 9'h95 == io_sel ? io_ins_149 : _GEN_148; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_150 = 9'h96 == io_sel ? io_ins_150 : _GEN_149; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_151 = 9'h97 == io_sel ? io_ins_151 : _GEN_150; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_152 = 9'h98 == io_sel ? io_ins_152 : _GEN_151; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_153 = 9'h99 == io_sel ? io_ins_153 : _GEN_152; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_154 = 9'h9a == io_sel ? io_ins_154 : _GEN_153; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_155 = 9'h9b == io_sel ? io_ins_155 : _GEN_154; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_156 = 9'h9c == io_sel ? io_ins_156 : _GEN_155; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_157 = 9'h9d == io_sel ? io_ins_157 : _GEN_156; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_158 = 9'h9e == io_sel ? io_ins_158 : _GEN_157; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_159 = 9'h9f == io_sel ? io_ins_159 : _GEN_158; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_160 = 9'ha0 == io_sel ? io_ins_160 : _GEN_159; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_161 = 9'ha1 == io_sel ? io_ins_161 : _GEN_160; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_162 = 9'ha2 == io_sel ? io_ins_162 : _GEN_161; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_163 = 9'ha3 == io_sel ? io_ins_163 : _GEN_162; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_164 = 9'ha4 == io_sel ? io_ins_164 : _GEN_163; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_165 = 9'ha5 == io_sel ? io_ins_165 : _GEN_164; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_166 = 9'ha6 == io_sel ? io_ins_166 : _GEN_165; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_167 = 9'ha7 == io_sel ? io_ins_167 : _GEN_166; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_168 = 9'ha8 == io_sel ? io_ins_168 : _GEN_167; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_169 = 9'ha9 == io_sel ? io_ins_169 : _GEN_168; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_170 = 9'haa == io_sel ? io_ins_170 : _GEN_169; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_171 = 9'hab == io_sel ? io_ins_171 : _GEN_170; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_172 = 9'hac == io_sel ? io_ins_172 : _GEN_171; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_173 = 9'had == io_sel ? io_ins_173 : _GEN_172; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_174 = 9'hae == io_sel ? io_ins_174 : _GEN_173; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_175 = 9'haf == io_sel ? io_ins_175 : _GEN_174; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_176 = 9'hb0 == io_sel ? io_ins_176 : _GEN_175; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_177 = 9'hb1 == io_sel ? io_ins_177 : _GEN_176; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_178 = 9'hb2 == io_sel ? io_ins_178 : _GEN_177; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_179 = 9'hb3 == io_sel ? io_ins_179 : _GEN_178; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_180 = 9'hb4 == io_sel ? io_ins_180 : _GEN_179; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_181 = 9'hb5 == io_sel ? io_ins_181 : _GEN_180; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_182 = 9'hb6 == io_sel ? io_ins_182 : _GEN_181; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_183 = 9'hb7 == io_sel ? io_ins_183 : _GEN_182; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_184 = 9'hb8 == io_sel ? io_ins_184 : _GEN_183; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_185 = 9'hb9 == io_sel ? io_ins_185 : _GEN_184; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_186 = 9'hba == io_sel ? io_ins_186 : _GEN_185; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_187 = 9'hbb == io_sel ? io_ins_187 : _GEN_186; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_188 = 9'hbc == io_sel ? io_ins_188 : _GEN_187; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_189 = 9'hbd == io_sel ? io_ins_189 : _GEN_188; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_190 = 9'hbe == io_sel ? io_ins_190 : _GEN_189; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_191 = 9'hbf == io_sel ? io_ins_191 : _GEN_190; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_192 = 9'hc0 == io_sel ? io_ins_192 : _GEN_191; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_193 = 9'hc1 == io_sel ? io_ins_193 : _GEN_192; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_194 = 9'hc2 == io_sel ? io_ins_194 : _GEN_193; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_195 = 9'hc3 == io_sel ? io_ins_195 : _GEN_194; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_196 = 9'hc4 == io_sel ? io_ins_196 : _GEN_195; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_197 = 9'hc5 == io_sel ? io_ins_197 : _GEN_196; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_198 = 9'hc6 == io_sel ? io_ins_198 : _GEN_197; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_199 = 9'hc7 == io_sel ? io_ins_199 : _GEN_198; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_200 = 9'hc8 == io_sel ? io_ins_200 : _GEN_199; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_201 = 9'hc9 == io_sel ? io_ins_201 : _GEN_200; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_202 = 9'hca == io_sel ? io_ins_202 : _GEN_201; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_203 = 9'hcb == io_sel ? io_ins_203 : _GEN_202; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_204 = 9'hcc == io_sel ? io_ins_204 : _GEN_203; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_205 = 9'hcd == io_sel ? io_ins_205 : _GEN_204; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_206 = 9'hce == io_sel ? io_ins_206 : _GEN_205; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_207 = 9'hcf == io_sel ? io_ins_207 : _GEN_206; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_208 = 9'hd0 == io_sel ? io_ins_208 : _GEN_207; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_209 = 9'hd1 == io_sel ? io_ins_209 : _GEN_208; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_210 = 9'hd2 == io_sel ? io_ins_210 : _GEN_209; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_211 = 9'hd3 == io_sel ? io_ins_211 : _GEN_210; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_212 = 9'hd4 == io_sel ? io_ins_212 : _GEN_211; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_213 = 9'hd5 == io_sel ? io_ins_213 : _GEN_212; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_214 = 9'hd6 == io_sel ? io_ins_214 : _GEN_213; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_215 = 9'hd7 == io_sel ? io_ins_215 : _GEN_214; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_216 = 9'hd8 == io_sel ? io_ins_216 : _GEN_215; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_217 = 9'hd9 == io_sel ? io_ins_217 : _GEN_216; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_218 = 9'hda == io_sel ? io_ins_218 : _GEN_217; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_219 = 9'hdb == io_sel ? io_ins_219 : _GEN_218; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_220 = 9'hdc == io_sel ? io_ins_220 : _GEN_219; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_221 = 9'hdd == io_sel ? io_ins_221 : _GEN_220; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_222 = 9'hde == io_sel ? io_ins_222 : _GEN_221; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_223 = 9'hdf == io_sel ? io_ins_223 : _GEN_222; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_224 = 9'he0 == io_sel ? io_ins_224 : _GEN_223; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_225 = 9'he1 == io_sel ? io_ins_225 : _GEN_224; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_226 = 9'he2 == io_sel ? io_ins_226 : _GEN_225; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_227 = 9'he3 == io_sel ? io_ins_227 : _GEN_226; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_228 = 9'he4 == io_sel ? io_ins_228 : _GEN_227; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_229 = 9'he5 == io_sel ? io_ins_229 : _GEN_228; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_230 = 9'he6 == io_sel ? io_ins_230 : _GEN_229; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_231 = 9'he7 == io_sel ? io_ins_231 : _GEN_230; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_232 = 9'he8 == io_sel ? io_ins_232 : _GEN_231; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_233 = 9'he9 == io_sel ? io_ins_233 : _GEN_232; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_234 = 9'hea == io_sel ? io_ins_234 : _GEN_233; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_235 = 9'heb == io_sel ? io_ins_235 : _GEN_234; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_236 = 9'hec == io_sel ? io_ins_236 : _GEN_235; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_237 = 9'hed == io_sel ? io_ins_237 : _GEN_236; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_238 = 9'hee == io_sel ? io_ins_238 : _GEN_237; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_239 = 9'hef == io_sel ? io_ins_239 : _GEN_238; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_240 = 9'hf0 == io_sel ? io_ins_240 : _GEN_239; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_241 = 9'hf1 == io_sel ? io_ins_241 : _GEN_240; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_242 = 9'hf2 == io_sel ? io_ins_242 : _GEN_241; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_243 = 9'hf3 == io_sel ? io_ins_243 : _GEN_242; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_244 = 9'hf4 == io_sel ? io_ins_244 : _GEN_243; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_245 = 9'hf5 == io_sel ? io_ins_245 : _GEN_244; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_246 = 9'hf6 == io_sel ? io_ins_246 : _GEN_245; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_247 = 9'hf7 == io_sel ? io_ins_247 : _GEN_246; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_248 = 9'hf8 == io_sel ? io_ins_248 : _GEN_247; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_249 = 9'hf9 == io_sel ? io_ins_249 : _GEN_248; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_250 = 9'hfa == io_sel ? io_ins_250 : _GEN_249; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_251 = 9'hfb == io_sel ? io_ins_251 : _GEN_250; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_252 = 9'hfc == io_sel ? io_ins_252 : _GEN_251; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_253 = 9'hfd == io_sel ? io_ins_253 : _GEN_252; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_254 = 9'hfe == io_sel ? io_ins_254 : _GEN_253; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_255 = 9'hff == io_sel ? io_ins_255 : _GEN_254; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_256 = 9'h100 == io_sel ? io_ins_256 : _GEN_255; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_257 = 9'h101 == io_sel ? io_ins_257 : _GEN_256; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_258 = 9'h102 == io_sel ? io_ins_258 : _GEN_257; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_259 = 9'h103 == io_sel ? io_ins_259 : _GEN_258; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_260 = 9'h104 == io_sel ? io_ins_260 : _GEN_259; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_261 = 9'h105 == io_sel ? io_ins_261 : _GEN_260; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_262 = 9'h106 == io_sel ? io_ins_262 : _GEN_261; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_263 = 9'h107 == io_sel ? io_ins_263 : _GEN_262; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_264 = 9'h108 == io_sel ? io_ins_264 : _GEN_263; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_265 = 9'h109 == io_sel ? io_ins_265 : _GEN_264; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_266 = 9'h10a == io_sel ? io_ins_266 : _GEN_265; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_267 = 9'h10b == io_sel ? io_ins_267 : _GEN_266; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_268 = 9'h10c == io_sel ? io_ins_268 : _GEN_267; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_269 = 9'h10d == io_sel ? io_ins_269 : _GEN_268; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_270 = 9'h10e == io_sel ? io_ins_270 : _GEN_269; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_271 = 9'h10f == io_sel ? io_ins_271 : _GEN_270; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_272 = 9'h110 == io_sel ? io_ins_272 : _GEN_271; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_273 = 9'h111 == io_sel ? io_ins_273 : _GEN_272; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_274 = 9'h112 == io_sel ? io_ins_274 : _GEN_273; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_275 = 9'h113 == io_sel ? io_ins_275 : _GEN_274; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_276 = 9'h114 == io_sel ? io_ins_276 : _GEN_275; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_277 = 9'h115 == io_sel ? io_ins_277 : _GEN_276; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_278 = 9'h116 == io_sel ? io_ins_278 : _GEN_277; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_279 = 9'h117 == io_sel ? io_ins_279 : _GEN_278; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_280 = 9'h118 == io_sel ? io_ins_280 : _GEN_279; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_281 = 9'h119 == io_sel ? io_ins_281 : _GEN_280; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_282 = 9'h11a == io_sel ? io_ins_282 : _GEN_281; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_283 = 9'h11b == io_sel ? io_ins_283 : _GEN_282; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_284 = 9'h11c == io_sel ? io_ins_284 : _GEN_283; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_285 = 9'h11d == io_sel ? io_ins_285 : _GEN_284; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_286 = 9'h11e == io_sel ? io_ins_286 : _GEN_285; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_287 = 9'h11f == io_sel ? io_ins_287 : _GEN_286; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_288 = 9'h120 == io_sel ? io_ins_288 : _GEN_287; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_289 = 9'h121 == io_sel ? io_ins_289 : _GEN_288; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_290 = 9'h122 == io_sel ? io_ins_290 : _GEN_289; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_291 = 9'h123 == io_sel ? io_ins_291 : _GEN_290; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_292 = 9'h124 == io_sel ? io_ins_292 : _GEN_291; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_293 = 9'h125 == io_sel ? io_ins_293 : _GEN_292; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_294 = 9'h126 == io_sel ? io_ins_294 : _GEN_293; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_295 = 9'h127 == io_sel ? io_ins_295 : _GEN_294; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_296 = 9'h128 == io_sel ? io_ins_296 : _GEN_295; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_297 = 9'h129 == io_sel ? io_ins_297 : _GEN_296; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_298 = 9'h12a == io_sel ? io_ins_298 : _GEN_297; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_299 = 9'h12b == io_sel ? io_ins_299 : _GEN_298; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_300 = 9'h12c == io_sel ? io_ins_300 : _GEN_299; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_301 = 9'h12d == io_sel ? io_ins_301 : _GEN_300; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_302 = 9'h12e == io_sel ? io_ins_302 : _GEN_301; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_303 = 9'h12f == io_sel ? io_ins_303 : _GEN_302; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_304 = 9'h130 == io_sel ? io_ins_304 : _GEN_303; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_305 = 9'h131 == io_sel ? io_ins_305 : _GEN_304; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_306 = 9'h132 == io_sel ? io_ins_306 : _GEN_305; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_307 = 9'h133 == io_sel ? io_ins_307 : _GEN_306; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_308 = 9'h134 == io_sel ? io_ins_308 : _GEN_307; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_309 = 9'h135 == io_sel ? io_ins_309 : _GEN_308; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_310 = 9'h136 == io_sel ? io_ins_310 : _GEN_309; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_311 = 9'h137 == io_sel ? io_ins_311 : _GEN_310; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_312 = 9'h138 == io_sel ? io_ins_312 : _GEN_311; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_313 = 9'h139 == io_sel ? io_ins_313 : _GEN_312; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_314 = 9'h13a == io_sel ? io_ins_314 : _GEN_313; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_315 = 9'h13b == io_sel ? io_ins_315 : _GEN_314; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_316 = 9'h13c == io_sel ? io_ins_316 : _GEN_315; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_317 = 9'h13d == io_sel ? io_ins_317 : _GEN_316; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_318 = 9'h13e == io_sel ? io_ins_318 : _GEN_317; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_319 = 9'h13f == io_sel ? io_ins_319 : _GEN_318; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_320 = 9'h140 == io_sel ? io_ins_320 : _GEN_319; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_321 = 9'h141 == io_sel ? io_ins_321 : _GEN_320; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_322 = 9'h142 == io_sel ? io_ins_322 : _GEN_321; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_323 = 9'h143 == io_sel ? io_ins_323 : _GEN_322; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_324 = 9'h144 == io_sel ? io_ins_324 : _GEN_323; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_325 = 9'h145 == io_sel ? io_ins_325 : _GEN_324; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_326 = 9'h146 == io_sel ? io_ins_326 : _GEN_325; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_327 = 9'h147 == io_sel ? io_ins_327 : _GEN_326; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_328 = 9'h148 == io_sel ? io_ins_328 : _GEN_327; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_329 = 9'h149 == io_sel ? io_ins_329 : _GEN_328; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_330 = 9'h14a == io_sel ? io_ins_330 : _GEN_329; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_331 = 9'h14b == io_sel ? io_ins_331 : _GEN_330; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_332 = 9'h14c == io_sel ? io_ins_332 : _GEN_331; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_333 = 9'h14d == io_sel ? io_ins_333 : _GEN_332; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_334 = 9'h14e == io_sel ? io_ins_334 : _GEN_333; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_335 = 9'h14f == io_sel ? io_ins_335 : _GEN_334; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_336 = 9'h150 == io_sel ? io_ins_336 : _GEN_335; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_337 = 9'h151 == io_sel ? io_ins_337 : _GEN_336; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_338 = 9'h152 == io_sel ? io_ins_338 : _GEN_337; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_339 = 9'h153 == io_sel ? io_ins_339 : _GEN_338; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_340 = 9'h154 == io_sel ? io_ins_340 : _GEN_339; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_341 = 9'h155 == io_sel ? io_ins_341 : _GEN_340; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_342 = 9'h156 == io_sel ? io_ins_342 : _GEN_341; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_343 = 9'h157 == io_sel ? io_ins_343 : _GEN_342; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_344 = 9'h158 == io_sel ? io_ins_344 : _GEN_343; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_345 = 9'h159 == io_sel ? io_ins_345 : _GEN_344; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_346 = 9'h15a == io_sel ? io_ins_346 : _GEN_345; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_347 = 9'h15b == io_sel ? io_ins_347 : _GEN_346; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_348 = 9'h15c == io_sel ? io_ins_348 : _GEN_347; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_349 = 9'h15d == io_sel ? io_ins_349 : _GEN_348; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_350 = 9'h15e == io_sel ? io_ins_350 : _GEN_349; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_351 = 9'h15f == io_sel ? io_ins_351 : _GEN_350; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_352 = 9'h160 == io_sel ? io_ins_352 : _GEN_351; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_353 = 9'h161 == io_sel ? io_ins_353 : _GEN_352; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_354 = 9'h162 == io_sel ? io_ins_354 : _GEN_353; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_355 = 9'h163 == io_sel ? io_ins_355 : _GEN_354; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_356 = 9'h164 == io_sel ? io_ins_356 : _GEN_355; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_357 = 9'h165 == io_sel ? io_ins_357 : _GEN_356; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_358 = 9'h166 == io_sel ? io_ins_358 : _GEN_357; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_359 = 9'h167 == io_sel ? io_ins_359 : _GEN_358; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_360 = 9'h168 == io_sel ? io_ins_360 : _GEN_359; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_361 = 9'h169 == io_sel ? io_ins_361 : _GEN_360; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_362 = 9'h16a == io_sel ? io_ins_362 : _GEN_361; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_363 = 9'h16b == io_sel ? io_ins_363 : _GEN_362; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_364 = 9'h16c == io_sel ? io_ins_364 : _GEN_363; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_365 = 9'h16d == io_sel ? io_ins_365 : _GEN_364; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_366 = 9'h16e == io_sel ? io_ins_366 : _GEN_365; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_367 = 9'h16f == io_sel ? io_ins_367 : _GEN_366; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_368 = 9'h170 == io_sel ? io_ins_368 : _GEN_367; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_369 = 9'h171 == io_sel ? io_ins_369 : _GEN_368; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_370 = 9'h172 == io_sel ? io_ins_370 : _GEN_369; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_371 = 9'h173 == io_sel ? io_ins_371 : _GEN_370; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_372 = 9'h174 == io_sel ? io_ins_372 : _GEN_371; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_373 = 9'h175 == io_sel ? io_ins_373 : _GEN_372; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_374 = 9'h176 == io_sel ? io_ins_374 : _GEN_373; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_375 = 9'h177 == io_sel ? io_ins_375 : _GEN_374; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_376 = 9'h178 == io_sel ? io_ins_376 : _GEN_375; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_377 = 9'h179 == io_sel ? io_ins_377 : _GEN_376; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_378 = 9'h17a == io_sel ? io_ins_378 : _GEN_377; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_379 = 9'h17b == io_sel ? io_ins_379 : _GEN_378; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_380 = 9'h17c == io_sel ? io_ins_380 : _GEN_379; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_381 = 9'h17d == io_sel ? io_ins_381 : _GEN_380; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_382 = 9'h17e == io_sel ? io_ins_382 : _GEN_381; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_383 = 9'h17f == io_sel ? io_ins_383 : _GEN_382; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_384 = 9'h180 == io_sel ? io_ins_384 : _GEN_383; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_385 = 9'h181 == io_sel ? io_ins_385 : _GEN_384; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_386 = 9'h182 == io_sel ? io_ins_386 : _GEN_385; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_387 = 9'h183 == io_sel ? io_ins_387 : _GEN_386; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_388 = 9'h184 == io_sel ? io_ins_388 : _GEN_387; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_389 = 9'h185 == io_sel ? io_ins_389 : _GEN_388; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_390 = 9'h186 == io_sel ? io_ins_390 : _GEN_389; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_391 = 9'h187 == io_sel ? io_ins_391 : _GEN_390; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_392 = 9'h188 == io_sel ? io_ins_392 : _GEN_391; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_393 = 9'h189 == io_sel ? io_ins_393 : _GEN_392; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_394 = 9'h18a == io_sel ? io_ins_394 : _GEN_393; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_395 = 9'h18b == io_sel ? io_ins_395 : _GEN_394; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_396 = 9'h18c == io_sel ? io_ins_396 : _GEN_395; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_397 = 9'h18d == io_sel ? io_ins_397 : _GEN_396; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_398 = 9'h18e == io_sel ? io_ins_398 : _GEN_397; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_399 = 9'h18f == io_sel ? io_ins_399 : _GEN_398; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_400 = 9'h190 == io_sel ? io_ins_400 : _GEN_399; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_401 = 9'h191 == io_sel ? io_ins_401 : _GEN_400; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_402 = 9'h192 == io_sel ? io_ins_402 : _GEN_401; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_403 = 9'h193 == io_sel ? io_ins_403 : _GEN_402; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_404 = 9'h194 == io_sel ? io_ins_404 : _GEN_403; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_405 = 9'h195 == io_sel ? io_ins_405 : _GEN_404; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_406 = 9'h196 == io_sel ? io_ins_406 : _GEN_405; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_407 = 9'h197 == io_sel ? io_ins_407 : _GEN_406; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_408 = 9'h198 == io_sel ? io_ins_408 : _GEN_407; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_409 = 9'h199 == io_sel ? io_ins_409 : _GEN_408; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_410 = 9'h19a == io_sel ? io_ins_410 : _GEN_409; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_411 = 9'h19b == io_sel ? io_ins_411 : _GEN_410; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_412 = 9'h19c == io_sel ? io_ins_412 : _GEN_411; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_413 = 9'h19d == io_sel ? io_ins_413 : _GEN_412; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_414 = 9'h19e == io_sel ? io_ins_414 : _GEN_413; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_415 = 9'h19f == io_sel ? io_ins_415 : _GEN_414; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_416 = 9'h1a0 == io_sel ? io_ins_416 : _GEN_415; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_417 = 9'h1a1 == io_sel ? io_ins_417 : _GEN_416; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_418 = 9'h1a2 == io_sel ? io_ins_418 : _GEN_417; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_419 = 9'h1a3 == io_sel ? io_ins_419 : _GEN_418; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_420 = 9'h1a4 == io_sel ? io_ins_420 : _GEN_419; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_421 = 9'h1a5 == io_sel ? io_ins_421 : _GEN_420; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_422 = 9'h1a6 == io_sel ? io_ins_422 : _GEN_421; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_423 = 9'h1a7 == io_sel ? io_ins_423 : _GEN_422; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_424 = 9'h1a8 == io_sel ? io_ins_424 : _GEN_423; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_425 = 9'h1a9 == io_sel ? io_ins_425 : _GEN_424; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_426 = 9'h1aa == io_sel ? io_ins_426 : _GEN_425; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_427 = 9'h1ab == io_sel ? io_ins_427 : _GEN_426; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_428 = 9'h1ac == io_sel ? io_ins_428 : _GEN_427; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_429 = 9'h1ad == io_sel ? io_ins_429 : _GEN_428; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_430 = 9'h1ae == io_sel ? io_ins_430 : _GEN_429; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_431 = 9'h1af == io_sel ? io_ins_431 : _GEN_430; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_432 = 9'h1b0 == io_sel ? io_ins_432 : _GEN_431; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_433 = 9'h1b1 == io_sel ? io_ins_433 : _GEN_432; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_434 = 9'h1b2 == io_sel ? io_ins_434 : _GEN_433; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_435 = 9'h1b3 == io_sel ? io_ins_435 : _GEN_434; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_436 = 9'h1b4 == io_sel ? io_ins_436 : _GEN_435; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_437 = 9'h1b5 == io_sel ? io_ins_437 : _GEN_436; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_438 = 9'h1b6 == io_sel ? io_ins_438 : _GEN_437; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_439 = 9'h1b7 == io_sel ? io_ins_439 : _GEN_438; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_440 = 9'h1b8 == io_sel ? io_ins_440 : _GEN_439; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_441 = 9'h1b9 == io_sel ? io_ins_441 : _GEN_440; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_442 = 9'h1ba == io_sel ? io_ins_442 : _GEN_441; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_443 = 9'h1bb == io_sel ? io_ins_443 : _GEN_442; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_444 = 9'h1bc == io_sel ? io_ins_444 : _GEN_443; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_445 = 9'h1bd == io_sel ? io_ins_445 : _GEN_444; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_446 = 9'h1be == io_sel ? io_ins_446 : _GEN_445; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_447 = 9'h1bf == io_sel ? io_ins_447 : _GEN_446; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_448 = 9'h1c0 == io_sel ? io_ins_448 : _GEN_447; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_449 = 9'h1c1 == io_sel ? io_ins_449 : _GEN_448; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_450 = 9'h1c2 == io_sel ? io_ins_450 : _GEN_449; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_451 = 9'h1c3 == io_sel ? io_ins_451 : _GEN_450; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_452 = 9'h1c4 == io_sel ? io_ins_452 : _GEN_451; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_453 = 9'h1c5 == io_sel ? io_ins_453 : _GEN_452; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_454 = 9'h1c6 == io_sel ? io_ins_454 : _GEN_453; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_455 = 9'h1c7 == io_sel ? io_ins_455 : _GEN_454; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_456 = 9'h1c8 == io_sel ? io_ins_456 : _GEN_455; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_457 = 9'h1c9 == io_sel ? io_ins_457 : _GEN_456; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_458 = 9'h1ca == io_sel ? io_ins_458 : _GEN_457; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_459 = 9'h1cb == io_sel ? io_ins_459 : _GEN_458; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_460 = 9'h1cc == io_sel ? io_ins_460 : _GEN_459; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_461 = 9'h1cd == io_sel ? io_ins_461 : _GEN_460; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_462 = 9'h1ce == io_sel ? io_ins_462 : _GEN_461; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_463 = 9'h1cf == io_sel ? io_ins_463 : _GEN_462; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_464 = 9'h1d0 == io_sel ? io_ins_464 : _GEN_463; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_465 = 9'h1d1 == io_sel ? io_ins_465 : _GEN_464; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_466 = 9'h1d2 == io_sel ? io_ins_466 : _GEN_465; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_467 = 9'h1d3 == io_sel ? io_ins_467 : _GEN_466; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_468 = 9'h1d4 == io_sel ? io_ins_468 : _GEN_467; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_469 = 9'h1d5 == io_sel ? io_ins_469 : _GEN_468; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_470 = 9'h1d6 == io_sel ? io_ins_470 : _GEN_469; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_471 = 9'h1d7 == io_sel ? io_ins_471 : _GEN_470; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_472 = 9'h1d8 == io_sel ? io_ins_472 : _GEN_471; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_473 = 9'h1d9 == io_sel ? io_ins_473 : _GEN_472; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_474 = 9'h1da == io_sel ? io_ins_474 : _GEN_473; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_475 = 9'h1db == io_sel ? io_ins_475 : _GEN_474; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_476 = 9'h1dc == io_sel ? io_ins_476 : _GEN_475; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_477 = 9'h1dd == io_sel ? io_ins_477 : _GEN_476; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_478 = 9'h1de == io_sel ? io_ins_478 : _GEN_477; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_479 = 9'h1df == io_sel ? io_ins_479 : _GEN_478; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_480 = 9'h1e0 == io_sel ? io_ins_480 : _GEN_479; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_481 = 9'h1e1 == io_sel ? io_ins_481 : _GEN_480; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_482 = 9'h1e2 == io_sel ? io_ins_482 : _GEN_481; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_483 = 9'h1e3 == io_sel ? io_ins_483 : _GEN_482; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_484 = 9'h1e4 == io_sel ? io_ins_484 : _GEN_483; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_485 = 9'h1e5 == io_sel ? io_ins_485 : _GEN_484; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_486 = 9'h1e6 == io_sel ? io_ins_486 : _GEN_485; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_487 = 9'h1e7 == io_sel ? io_ins_487 : _GEN_486; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_488 = 9'h1e8 == io_sel ? io_ins_488 : _GEN_487; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_489 = 9'h1e9 == io_sel ? io_ins_489 : _GEN_488; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_490 = 9'h1ea == io_sel ? io_ins_490 : _GEN_489; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_491 = 9'h1eb == io_sel ? io_ins_491 : _GEN_490; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_492 = 9'h1ec == io_sel ? io_ins_492 : _GEN_491; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_493 = 9'h1ed == io_sel ? io_ins_493 : _GEN_492; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_494 = 9'h1ee == io_sel ? io_ins_494 : _GEN_493; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_495 = 9'h1ef == io_sel ? io_ins_495 : _GEN_494; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_496 = 9'h1f0 == io_sel ? io_ins_496 : _GEN_495; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_497 = 9'h1f1 == io_sel ? io_ins_497 : _GEN_496; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_498 = 9'h1f2 == io_sel ? io_ins_498 : _GEN_497; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_499 = 9'h1f3 == io_sel ? io_ins_499 : _GEN_498; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_500 = 9'h1f4 == io_sel ? io_ins_500 : _GEN_499; // @[MuxN.scala 16:10:@122976.4]
  assign _GEN_501 = 9'h1f5 == io_sel ? io_ins_501 : _GEN_500; // @[MuxN.scala 16:10:@122976.4]
  assign io_out = 9'h1f6 == io_sel ? io_ins_502 : _GEN_501; // @[MuxN.scala 16:10:@122976.4]
endmodule
module RegFile( // @[:@122978.2]
  input         clock, // @[:@122979.4]
  input         reset, // @[:@122980.4]
  input  [31:0] io_raddr, // @[:@122981.4]
  input         io_wen, // @[:@122981.4]
  input  [31:0] io_waddr, // @[:@122981.4]
  input  [63:0] io_wdata, // @[:@122981.4]
  output [63:0] io_rdata, // @[:@122981.4]
  input         io_reset, // @[:@122981.4]
  output [63:0] io_argIns_0, // @[:@122981.4]
  output [63:0] io_argIns_1, // @[:@122981.4]
  output [63:0] io_argIns_2, // @[:@122981.4]
  output [63:0] io_argIns_3, // @[:@122981.4]
  input         io_argOuts_0_valid, // @[:@122981.4]
  input  [63:0] io_argOuts_0_bits, // @[:@122981.4]
  input         io_argOuts_1_valid, // @[:@122981.4]
  input  [63:0] io_argOuts_1_bits // @[:@122981.4]
);
  wire  regs_0_clock; // @[RegFile.scala 66:20:@124991.4]
  wire  regs_0_reset; // @[RegFile.scala 66:20:@124991.4]
  wire [63:0] regs_0_io_in; // @[RegFile.scala 66:20:@124991.4]
  wire  regs_0_io_reset; // @[RegFile.scala 66:20:@124991.4]
  wire [63:0] regs_0_io_out; // @[RegFile.scala 66:20:@124991.4]
  wire  regs_0_io_enable; // @[RegFile.scala 66:20:@124991.4]
  wire  regs_1_clock; // @[RegFile.scala 66:20:@125003.4]
  wire  regs_1_reset; // @[RegFile.scala 66:20:@125003.4]
  wire [63:0] regs_1_io_in; // @[RegFile.scala 66:20:@125003.4]
  wire  regs_1_io_reset; // @[RegFile.scala 66:20:@125003.4]
  wire [63:0] regs_1_io_out; // @[RegFile.scala 66:20:@125003.4]
  wire  regs_1_io_enable; // @[RegFile.scala 66:20:@125003.4]
  wire  regs_2_clock; // @[RegFile.scala 66:20:@125022.4]
  wire  regs_2_reset; // @[RegFile.scala 66:20:@125022.4]
  wire [63:0] regs_2_io_in; // @[RegFile.scala 66:20:@125022.4]
  wire  regs_2_io_reset; // @[RegFile.scala 66:20:@125022.4]
  wire [63:0] regs_2_io_out; // @[RegFile.scala 66:20:@125022.4]
  wire  regs_2_io_enable; // @[RegFile.scala 66:20:@125022.4]
  wire  regs_3_clock; // @[RegFile.scala 66:20:@125034.4]
  wire  regs_3_reset; // @[RegFile.scala 66:20:@125034.4]
  wire [63:0] regs_3_io_in; // @[RegFile.scala 66:20:@125034.4]
  wire  regs_3_io_reset; // @[RegFile.scala 66:20:@125034.4]
  wire [63:0] regs_3_io_out; // @[RegFile.scala 66:20:@125034.4]
  wire  regs_3_io_enable; // @[RegFile.scala 66:20:@125034.4]
  wire  regs_4_clock; // @[RegFile.scala 66:20:@125046.4]
  wire  regs_4_reset; // @[RegFile.scala 66:20:@125046.4]
  wire [63:0] regs_4_io_in; // @[RegFile.scala 66:20:@125046.4]
  wire  regs_4_io_reset; // @[RegFile.scala 66:20:@125046.4]
  wire [63:0] regs_4_io_out; // @[RegFile.scala 66:20:@125046.4]
  wire  regs_4_io_enable; // @[RegFile.scala 66:20:@125046.4]
  wire  regs_5_clock; // @[RegFile.scala 66:20:@125060.4]
  wire  regs_5_reset; // @[RegFile.scala 66:20:@125060.4]
  wire [63:0] regs_5_io_in; // @[RegFile.scala 66:20:@125060.4]
  wire  regs_5_io_reset; // @[RegFile.scala 66:20:@125060.4]
  wire [63:0] regs_5_io_out; // @[RegFile.scala 66:20:@125060.4]
  wire  regs_5_io_enable; // @[RegFile.scala 66:20:@125060.4]
  wire  regs_6_clock; // @[RegFile.scala 66:20:@125074.4]
  wire  regs_6_reset; // @[RegFile.scala 66:20:@125074.4]
  wire [63:0] regs_6_io_in; // @[RegFile.scala 66:20:@125074.4]
  wire  regs_6_io_reset; // @[RegFile.scala 66:20:@125074.4]
  wire [63:0] regs_6_io_out; // @[RegFile.scala 66:20:@125074.4]
  wire  regs_6_io_enable; // @[RegFile.scala 66:20:@125074.4]
  wire  regs_7_clock; // @[RegFile.scala 66:20:@125088.4]
  wire  regs_7_reset; // @[RegFile.scala 66:20:@125088.4]
  wire [63:0] regs_7_io_in; // @[RegFile.scala 66:20:@125088.4]
  wire  regs_7_io_reset; // @[RegFile.scala 66:20:@125088.4]
  wire [63:0] regs_7_io_out; // @[RegFile.scala 66:20:@125088.4]
  wire  regs_7_io_enable; // @[RegFile.scala 66:20:@125088.4]
  wire  regs_8_clock; // @[RegFile.scala 66:20:@125102.4]
  wire  regs_8_reset; // @[RegFile.scala 66:20:@125102.4]
  wire [63:0] regs_8_io_in; // @[RegFile.scala 66:20:@125102.4]
  wire  regs_8_io_reset; // @[RegFile.scala 66:20:@125102.4]
  wire [63:0] regs_8_io_out; // @[RegFile.scala 66:20:@125102.4]
  wire  regs_8_io_enable; // @[RegFile.scala 66:20:@125102.4]
  wire  regs_9_clock; // @[RegFile.scala 66:20:@125116.4]
  wire  regs_9_reset; // @[RegFile.scala 66:20:@125116.4]
  wire [63:0] regs_9_io_in; // @[RegFile.scala 66:20:@125116.4]
  wire  regs_9_io_reset; // @[RegFile.scala 66:20:@125116.4]
  wire [63:0] regs_9_io_out; // @[RegFile.scala 66:20:@125116.4]
  wire  regs_9_io_enable; // @[RegFile.scala 66:20:@125116.4]
  wire  regs_10_clock; // @[RegFile.scala 66:20:@125130.4]
  wire  regs_10_reset; // @[RegFile.scala 66:20:@125130.4]
  wire [63:0] regs_10_io_in; // @[RegFile.scala 66:20:@125130.4]
  wire  regs_10_io_reset; // @[RegFile.scala 66:20:@125130.4]
  wire [63:0] regs_10_io_out; // @[RegFile.scala 66:20:@125130.4]
  wire  regs_10_io_enable; // @[RegFile.scala 66:20:@125130.4]
  wire  regs_11_clock; // @[RegFile.scala 66:20:@125144.4]
  wire  regs_11_reset; // @[RegFile.scala 66:20:@125144.4]
  wire [63:0] regs_11_io_in; // @[RegFile.scala 66:20:@125144.4]
  wire  regs_11_io_reset; // @[RegFile.scala 66:20:@125144.4]
  wire [63:0] regs_11_io_out; // @[RegFile.scala 66:20:@125144.4]
  wire  regs_11_io_enable; // @[RegFile.scala 66:20:@125144.4]
  wire  regs_12_clock; // @[RegFile.scala 66:20:@125158.4]
  wire  regs_12_reset; // @[RegFile.scala 66:20:@125158.4]
  wire [63:0] regs_12_io_in; // @[RegFile.scala 66:20:@125158.4]
  wire  regs_12_io_reset; // @[RegFile.scala 66:20:@125158.4]
  wire [63:0] regs_12_io_out; // @[RegFile.scala 66:20:@125158.4]
  wire  regs_12_io_enable; // @[RegFile.scala 66:20:@125158.4]
  wire  regs_13_clock; // @[RegFile.scala 66:20:@125172.4]
  wire  regs_13_reset; // @[RegFile.scala 66:20:@125172.4]
  wire [63:0] regs_13_io_in; // @[RegFile.scala 66:20:@125172.4]
  wire  regs_13_io_reset; // @[RegFile.scala 66:20:@125172.4]
  wire [63:0] regs_13_io_out; // @[RegFile.scala 66:20:@125172.4]
  wire  regs_13_io_enable; // @[RegFile.scala 66:20:@125172.4]
  wire  regs_14_clock; // @[RegFile.scala 66:20:@125186.4]
  wire  regs_14_reset; // @[RegFile.scala 66:20:@125186.4]
  wire [63:0] regs_14_io_in; // @[RegFile.scala 66:20:@125186.4]
  wire  regs_14_io_reset; // @[RegFile.scala 66:20:@125186.4]
  wire [63:0] regs_14_io_out; // @[RegFile.scala 66:20:@125186.4]
  wire  regs_14_io_enable; // @[RegFile.scala 66:20:@125186.4]
  wire  regs_15_clock; // @[RegFile.scala 66:20:@125200.4]
  wire  regs_15_reset; // @[RegFile.scala 66:20:@125200.4]
  wire [63:0] regs_15_io_in; // @[RegFile.scala 66:20:@125200.4]
  wire  regs_15_io_reset; // @[RegFile.scala 66:20:@125200.4]
  wire [63:0] regs_15_io_out; // @[RegFile.scala 66:20:@125200.4]
  wire  regs_15_io_enable; // @[RegFile.scala 66:20:@125200.4]
  wire  regs_16_clock; // @[RegFile.scala 66:20:@125214.4]
  wire  regs_16_reset; // @[RegFile.scala 66:20:@125214.4]
  wire [63:0] regs_16_io_in; // @[RegFile.scala 66:20:@125214.4]
  wire  regs_16_io_reset; // @[RegFile.scala 66:20:@125214.4]
  wire [63:0] regs_16_io_out; // @[RegFile.scala 66:20:@125214.4]
  wire  regs_16_io_enable; // @[RegFile.scala 66:20:@125214.4]
  wire  regs_17_clock; // @[RegFile.scala 66:20:@125228.4]
  wire  regs_17_reset; // @[RegFile.scala 66:20:@125228.4]
  wire [63:0] regs_17_io_in; // @[RegFile.scala 66:20:@125228.4]
  wire  regs_17_io_reset; // @[RegFile.scala 66:20:@125228.4]
  wire [63:0] regs_17_io_out; // @[RegFile.scala 66:20:@125228.4]
  wire  regs_17_io_enable; // @[RegFile.scala 66:20:@125228.4]
  wire  regs_18_clock; // @[RegFile.scala 66:20:@125242.4]
  wire  regs_18_reset; // @[RegFile.scala 66:20:@125242.4]
  wire [63:0] regs_18_io_in; // @[RegFile.scala 66:20:@125242.4]
  wire  regs_18_io_reset; // @[RegFile.scala 66:20:@125242.4]
  wire [63:0] regs_18_io_out; // @[RegFile.scala 66:20:@125242.4]
  wire  regs_18_io_enable; // @[RegFile.scala 66:20:@125242.4]
  wire  regs_19_clock; // @[RegFile.scala 66:20:@125256.4]
  wire  regs_19_reset; // @[RegFile.scala 66:20:@125256.4]
  wire [63:0] regs_19_io_in; // @[RegFile.scala 66:20:@125256.4]
  wire  regs_19_io_reset; // @[RegFile.scala 66:20:@125256.4]
  wire [63:0] regs_19_io_out; // @[RegFile.scala 66:20:@125256.4]
  wire  regs_19_io_enable; // @[RegFile.scala 66:20:@125256.4]
  wire  regs_20_clock; // @[RegFile.scala 66:20:@125270.4]
  wire  regs_20_reset; // @[RegFile.scala 66:20:@125270.4]
  wire [63:0] regs_20_io_in; // @[RegFile.scala 66:20:@125270.4]
  wire  regs_20_io_reset; // @[RegFile.scala 66:20:@125270.4]
  wire [63:0] regs_20_io_out; // @[RegFile.scala 66:20:@125270.4]
  wire  regs_20_io_enable; // @[RegFile.scala 66:20:@125270.4]
  wire  regs_21_clock; // @[RegFile.scala 66:20:@125284.4]
  wire  regs_21_reset; // @[RegFile.scala 66:20:@125284.4]
  wire [63:0] regs_21_io_in; // @[RegFile.scala 66:20:@125284.4]
  wire  regs_21_io_reset; // @[RegFile.scala 66:20:@125284.4]
  wire [63:0] regs_21_io_out; // @[RegFile.scala 66:20:@125284.4]
  wire  regs_21_io_enable; // @[RegFile.scala 66:20:@125284.4]
  wire  regs_22_clock; // @[RegFile.scala 66:20:@125298.4]
  wire  regs_22_reset; // @[RegFile.scala 66:20:@125298.4]
  wire [63:0] regs_22_io_in; // @[RegFile.scala 66:20:@125298.4]
  wire  regs_22_io_reset; // @[RegFile.scala 66:20:@125298.4]
  wire [63:0] regs_22_io_out; // @[RegFile.scala 66:20:@125298.4]
  wire  regs_22_io_enable; // @[RegFile.scala 66:20:@125298.4]
  wire  regs_23_clock; // @[RegFile.scala 66:20:@125312.4]
  wire  regs_23_reset; // @[RegFile.scala 66:20:@125312.4]
  wire [63:0] regs_23_io_in; // @[RegFile.scala 66:20:@125312.4]
  wire  regs_23_io_reset; // @[RegFile.scala 66:20:@125312.4]
  wire [63:0] regs_23_io_out; // @[RegFile.scala 66:20:@125312.4]
  wire  regs_23_io_enable; // @[RegFile.scala 66:20:@125312.4]
  wire  regs_24_clock; // @[RegFile.scala 66:20:@125326.4]
  wire  regs_24_reset; // @[RegFile.scala 66:20:@125326.4]
  wire [63:0] regs_24_io_in; // @[RegFile.scala 66:20:@125326.4]
  wire  regs_24_io_reset; // @[RegFile.scala 66:20:@125326.4]
  wire [63:0] regs_24_io_out; // @[RegFile.scala 66:20:@125326.4]
  wire  regs_24_io_enable; // @[RegFile.scala 66:20:@125326.4]
  wire  regs_25_clock; // @[RegFile.scala 66:20:@125340.4]
  wire  regs_25_reset; // @[RegFile.scala 66:20:@125340.4]
  wire [63:0] regs_25_io_in; // @[RegFile.scala 66:20:@125340.4]
  wire  regs_25_io_reset; // @[RegFile.scala 66:20:@125340.4]
  wire [63:0] regs_25_io_out; // @[RegFile.scala 66:20:@125340.4]
  wire  regs_25_io_enable; // @[RegFile.scala 66:20:@125340.4]
  wire  regs_26_clock; // @[RegFile.scala 66:20:@125354.4]
  wire  regs_26_reset; // @[RegFile.scala 66:20:@125354.4]
  wire [63:0] regs_26_io_in; // @[RegFile.scala 66:20:@125354.4]
  wire  regs_26_io_reset; // @[RegFile.scala 66:20:@125354.4]
  wire [63:0] regs_26_io_out; // @[RegFile.scala 66:20:@125354.4]
  wire  regs_26_io_enable; // @[RegFile.scala 66:20:@125354.4]
  wire  regs_27_clock; // @[RegFile.scala 66:20:@125368.4]
  wire  regs_27_reset; // @[RegFile.scala 66:20:@125368.4]
  wire [63:0] regs_27_io_in; // @[RegFile.scala 66:20:@125368.4]
  wire  regs_27_io_reset; // @[RegFile.scala 66:20:@125368.4]
  wire [63:0] regs_27_io_out; // @[RegFile.scala 66:20:@125368.4]
  wire  regs_27_io_enable; // @[RegFile.scala 66:20:@125368.4]
  wire  regs_28_clock; // @[RegFile.scala 66:20:@125382.4]
  wire  regs_28_reset; // @[RegFile.scala 66:20:@125382.4]
  wire [63:0] regs_28_io_in; // @[RegFile.scala 66:20:@125382.4]
  wire  regs_28_io_reset; // @[RegFile.scala 66:20:@125382.4]
  wire [63:0] regs_28_io_out; // @[RegFile.scala 66:20:@125382.4]
  wire  regs_28_io_enable; // @[RegFile.scala 66:20:@125382.4]
  wire  regs_29_clock; // @[RegFile.scala 66:20:@125396.4]
  wire  regs_29_reset; // @[RegFile.scala 66:20:@125396.4]
  wire [63:0] regs_29_io_in; // @[RegFile.scala 66:20:@125396.4]
  wire  regs_29_io_reset; // @[RegFile.scala 66:20:@125396.4]
  wire [63:0] regs_29_io_out; // @[RegFile.scala 66:20:@125396.4]
  wire  regs_29_io_enable; // @[RegFile.scala 66:20:@125396.4]
  wire  regs_30_clock; // @[RegFile.scala 66:20:@125410.4]
  wire  regs_30_reset; // @[RegFile.scala 66:20:@125410.4]
  wire [63:0] regs_30_io_in; // @[RegFile.scala 66:20:@125410.4]
  wire  regs_30_io_reset; // @[RegFile.scala 66:20:@125410.4]
  wire [63:0] regs_30_io_out; // @[RegFile.scala 66:20:@125410.4]
  wire  regs_30_io_enable; // @[RegFile.scala 66:20:@125410.4]
  wire  regs_31_clock; // @[RegFile.scala 66:20:@125424.4]
  wire  regs_31_reset; // @[RegFile.scala 66:20:@125424.4]
  wire [63:0] regs_31_io_in; // @[RegFile.scala 66:20:@125424.4]
  wire  regs_31_io_reset; // @[RegFile.scala 66:20:@125424.4]
  wire [63:0] regs_31_io_out; // @[RegFile.scala 66:20:@125424.4]
  wire  regs_31_io_enable; // @[RegFile.scala 66:20:@125424.4]
  wire  regs_32_clock; // @[RegFile.scala 66:20:@125438.4]
  wire  regs_32_reset; // @[RegFile.scala 66:20:@125438.4]
  wire [63:0] regs_32_io_in; // @[RegFile.scala 66:20:@125438.4]
  wire  regs_32_io_reset; // @[RegFile.scala 66:20:@125438.4]
  wire [63:0] regs_32_io_out; // @[RegFile.scala 66:20:@125438.4]
  wire  regs_32_io_enable; // @[RegFile.scala 66:20:@125438.4]
  wire  regs_33_clock; // @[RegFile.scala 66:20:@125452.4]
  wire  regs_33_reset; // @[RegFile.scala 66:20:@125452.4]
  wire [63:0] regs_33_io_in; // @[RegFile.scala 66:20:@125452.4]
  wire  regs_33_io_reset; // @[RegFile.scala 66:20:@125452.4]
  wire [63:0] regs_33_io_out; // @[RegFile.scala 66:20:@125452.4]
  wire  regs_33_io_enable; // @[RegFile.scala 66:20:@125452.4]
  wire  regs_34_clock; // @[RegFile.scala 66:20:@125466.4]
  wire  regs_34_reset; // @[RegFile.scala 66:20:@125466.4]
  wire [63:0] regs_34_io_in; // @[RegFile.scala 66:20:@125466.4]
  wire  regs_34_io_reset; // @[RegFile.scala 66:20:@125466.4]
  wire [63:0] regs_34_io_out; // @[RegFile.scala 66:20:@125466.4]
  wire  regs_34_io_enable; // @[RegFile.scala 66:20:@125466.4]
  wire  regs_35_clock; // @[RegFile.scala 66:20:@125480.4]
  wire  regs_35_reset; // @[RegFile.scala 66:20:@125480.4]
  wire [63:0] regs_35_io_in; // @[RegFile.scala 66:20:@125480.4]
  wire  regs_35_io_reset; // @[RegFile.scala 66:20:@125480.4]
  wire [63:0] regs_35_io_out; // @[RegFile.scala 66:20:@125480.4]
  wire  regs_35_io_enable; // @[RegFile.scala 66:20:@125480.4]
  wire  regs_36_clock; // @[RegFile.scala 66:20:@125494.4]
  wire  regs_36_reset; // @[RegFile.scala 66:20:@125494.4]
  wire [63:0] regs_36_io_in; // @[RegFile.scala 66:20:@125494.4]
  wire  regs_36_io_reset; // @[RegFile.scala 66:20:@125494.4]
  wire [63:0] regs_36_io_out; // @[RegFile.scala 66:20:@125494.4]
  wire  regs_36_io_enable; // @[RegFile.scala 66:20:@125494.4]
  wire  regs_37_clock; // @[RegFile.scala 66:20:@125508.4]
  wire  regs_37_reset; // @[RegFile.scala 66:20:@125508.4]
  wire [63:0] regs_37_io_in; // @[RegFile.scala 66:20:@125508.4]
  wire  regs_37_io_reset; // @[RegFile.scala 66:20:@125508.4]
  wire [63:0] regs_37_io_out; // @[RegFile.scala 66:20:@125508.4]
  wire  regs_37_io_enable; // @[RegFile.scala 66:20:@125508.4]
  wire  regs_38_clock; // @[RegFile.scala 66:20:@125522.4]
  wire  regs_38_reset; // @[RegFile.scala 66:20:@125522.4]
  wire [63:0] regs_38_io_in; // @[RegFile.scala 66:20:@125522.4]
  wire  regs_38_io_reset; // @[RegFile.scala 66:20:@125522.4]
  wire [63:0] regs_38_io_out; // @[RegFile.scala 66:20:@125522.4]
  wire  regs_38_io_enable; // @[RegFile.scala 66:20:@125522.4]
  wire  regs_39_clock; // @[RegFile.scala 66:20:@125536.4]
  wire  regs_39_reset; // @[RegFile.scala 66:20:@125536.4]
  wire [63:0] regs_39_io_in; // @[RegFile.scala 66:20:@125536.4]
  wire  regs_39_io_reset; // @[RegFile.scala 66:20:@125536.4]
  wire [63:0] regs_39_io_out; // @[RegFile.scala 66:20:@125536.4]
  wire  regs_39_io_enable; // @[RegFile.scala 66:20:@125536.4]
  wire  regs_40_clock; // @[RegFile.scala 66:20:@125550.4]
  wire  regs_40_reset; // @[RegFile.scala 66:20:@125550.4]
  wire [63:0] regs_40_io_in; // @[RegFile.scala 66:20:@125550.4]
  wire  regs_40_io_reset; // @[RegFile.scala 66:20:@125550.4]
  wire [63:0] regs_40_io_out; // @[RegFile.scala 66:20:@125550.4]
  wire  regs_40_io_enable; // @[RegFile.scala 66:20:@125550.4]
  wire  regs_41_clock; // @[RegFile.scala 66:20:@125564.4]
  wire  regs_41_reset; // @[RegFile.scala 66:20:@125564.4]
  wire [63:0] regs_41_io_in; // @[RegFile.scala 66:20:@125564.4]
  wire  regs_41_io_reset; // @[RegFile.scala 66:20:@125564.4]
  wire [63:0] regs_41_io_out; // @[RegFile.scala 66:20:@125564.4]
  wire  regs_41_io_enable; // @[RegFile.scala 66:20:@125564.4]
  wire  regs_42_clock; // @[RegFile.scala 66:20:@125578.4]
  wire  regs_42_reset; // @[RegFile.scala 66:20:@125578.4]
  wire [63:0] regs_42_io_in; // @[RegFile.scala 66:20:@125578.4]
  wire  regs_42_io_reset; // @[RegFile.scala 66:20:@125578.4]
  wire [63:0] regs_42_io_out; // @[RegFile.scala 66:20:@125578.4]
  wire  regs_42_io_enable; // @[RegFile.scala 66:20:@125578.4]
  wire  regs_43_clock; // @[RegFile.scala 66:20:@125592.4]
  wire  regs_43_reset; // @[RegFile.scala 66:20:@125592.4]
  wire [63:0] regs_43_io_in; // @[RegFile.scala 66:20:@125592.4]
  wire  regs_43_io_reset; // @[RegFile.scala 66:20:@125592.4]
  wire [63:0] regs_43_io_out; // @[RegFile.scala 66:20:@125592.4]
  wire  regs_43_io_enable; // @[RegFile.scala 66:20:@125592.4]
  wire  regs_44_clock; // @[RegFile.scala 66:20:@125606.4]
  wire  regs_44_reset; // @[RegFile.scala 66:20:@125606.4]
  wire [63:0] regs_44_io_in; // @[RegFile.scala 66:20:@125606.4]
  wire  regs_44_io_reset; // @[RegFile.scala 66:20:@125606.4]
  wire [63:0] regs_44_io_out; // @[RegFile.scala 66:20:@125606.4]
  wire  regs_44_io_enable; // @[RegFile.scala 66:20:@125606.4]
  wire  regs_45_clock; // @[RegFile.scala 66:20:@125620.4]
  wire  regs_45_reset; // @[RegFile.scala 66:20:@125620.4]
  wire [63:0] regs_45_io_in; // @[RegFile.scala 66:20:@125620.4]
  wire  regs_45_io_reset; // @[RegFile.scala 66:20:@125620.4]
  wire [63:0] regs_45_io_out; // @[RegFile.scala 66:20:@125620.4]
  wire  regs_45_io_enable; // @[RegFile.scala 66:20:@125620.4]
  wire  regs_46_clock; // @[RegFile.scala 66:20:@125634.4]
  wire  regs_46_reset; // @[RegFile.scala 66:20:@125634.4]
  wire [63:0] regs_46_io_in; // @[RegFile.scala 66:20:@125634.4]
  wire  regs_46_io_reset; // @[RegFile.scala 66:20:@125634.4]
  wire [63:0] regs_46_io_out; // @[RegFile.scala 66:20:@125634.4]
  wire  regs_46_io_enable; // @[RegFile.scala 66:20:@125634.4]
  wire  regs_47_clock; // @[RegFile.scala 66:20:@125648.4]
  wire  regs_47_reset; // @[RegFile.scala 66:20:@125648.4]
  wire [63:0] regs_47_io_in; // @[RegFile.scala 66:20:@125648.4]
  wire  regs_47_io_reset; // @[RegFile.scala 66:20:@125648.4]
  wire [63:0] regs_47_io_out; // @[RegFile.scala 66:20:@125648.4]
  wire  regs_47_io_enable; // @[RegFile.scala 66:20:@125648.4]
  wire  regs_48_clock; // @[RegFile.scala 66:20:@125662.4]
  wire  regs_48_reset; // @[RegFile.scala 66:20:@125662.4]
  wire [63:0] regs_48_io_in; // @[RegFile.scala 66:20:@125662.4]
  wire  regs_48_io_reset; // @[RegFile.scala 66:20:@125662.4]
  wire [63:0] regs_48_io_out; // @[RegFile.scala 66:20:@125662.4]
  wire  regs_48_io_enable; // @[RegFile.scala 66:20:@125662.4]
  wire  regs_49_clock; // @[RegFile.scala 66:20:@125676.4]
  wire  regs_49_reset; // @[RegFile.scala 66:20:@125676.4]
  wire [63:0] regs_49_io_in; // @[RegFile.scala 66:20:@125676.4]
  wire  regs_49_io_reset; // @[RegFile.scala 66:20:@125676.4]
  wire [63:0] regs_49_io_out; // @[RegFile.scala 66:20:@125676.4]
  wire  regs_49_io_enable; // @[RegFile.scala 66:20:@125676.4]
  wire  regs_50_clock; // @[RegFile.scala 66:20:@125690.4]
  wire  regs_50_reset; // @[RegFile.scala 66:20:@125690.4]
  wire [63:0] regs_50_io_in; // @[RegFile.scala 66:20:@125690.4]
  wire  regs_50_io_reset; // @[RegFile.scala 66:20:@125690.4]
  wire [63:0] regs_50_io_out; // @[RegFile.scala 66:20:@125690.4]
  wire  regs_50_io_enable; // @[RegFile.scala 66:20:@125690.4]
  wire  regs_51_clock; // @[RegFile.scala 66:20:@125704.4]
  wire  regs_51_reset; // @[RegFile.scala 66:20:@125704.4]
  wire [63:0] regs_51_io_in; // @[RegFile.scala 66:20:@125704.4]
  wire  regs_51_io_reset; // @[RegFile.scala 66:20:@125704.4]
  wire [63:0] regs_51_io_out; // @[RegFile.scala 66:20:@125704.4]
  wire  regs_51_io_enable; // @[RegFile.scala 66:20:@125704.4]
  wire  regs_52_clock; // @[RegFile.scala 66:20:@125718.4]
  wire  regs_52_reset; // @[RegFile.scala 66:20:@125718.4]
  wire [63:0] regs_52_io_in; // @[RegFile.scala 66:20:@125718.4]
  wire  regs_52_io_reset; // @[RegFile.scala 66:20:@125718.4]
  wire [63:0] regs_52_io_out; // @[RegFile.scala 66:20:@125718.4]
  wire  regs_52_io_enable; // @[RegFile.scala 66:20:@125718.4]
  wire  regs_53_clock; // @[RegFile.scala 66:20:@125732.4]
  wire  regs_53_reset; // @[RegFile.scala 66:20:@125732.4]
  wire [63:0] regs_53_io_in; // @[RegFile.scala 66:20:@125732.4]
  wire  regs_53_io_reset; // @[RegFile.scala 66:20:@125732.4]
  wire [63:0] regs_53_io_out; // @[RegFile.scala 66:20:@125732.4]
  wire  regs_53_io_enable; // @[RegFile.scala 66:20:@125732.4]
  wire  regs_54_clock; // @[RegFile.scala 66:20:@125746.4]
  wire  regs_54_reset; // @[RegFile.scala 66:20:@125746.4]
  wire [63:0] regs_54_io_in; // @[RegFile.scala 66:20:@125746.4]
  wire  regs_54_io_reset; // @[RegFile.scala 66:20:@125746.4]
  wire [63:0] regs_54_io_out; // @[RegFile.scala 66:20:@125746.4]
  wire  regs_54_io_enable; // @[RegFile.scala 66:20:@125746.4]
  wire  regs_55_clock; // @[RegFile.scala 66:20:@125760.4]
  wire  regs_55_reset; // @[RegFile.scala 66:20:@125760.4]
  wire [63:0] regs_55_io_in; // @[RegFile.scala 66:20:@125760.4]
  wire  regs_55_io_reset; // @[RegFile.scala 66:20:@125760.4]
  wire [63:0] regs_55_io_out; // @[RegFile.scala 66:20:@125760.4]
  wire  regs_55_io_enable; // @[RegFile.scala 66:20:@125760.4]
  wire  regs_56_clock; // @[RegFile.scala 66:20:@125774.4]
  wire  regs_56_reset; // @[RegFile.scala 66:20:@125774.4]
  wire [63:0] regs_56_io_in; // @[RegFile.scala 66:20:@125774.4]
  wire  regs_56_io_reset; // @[RegFile.scala 66:20:@125774.4]
  wire [63:0] regs_56_io_out; // @[RegFile.scala 66:20:@125774.4]
  wire  regs_56_io_enable; // @[RegFile.scala 66:20:@125774.4]
  wire  regs_57_clock; // @[RegFile.scala 66:20:@125788.4]
  wire  regs_57_reset; // @[RegFile.scala 66:20:@125788.4]
  wire [63:0] regs_57_io_in; // @[RegFile.scala 66:20:@125788.4]
  wire  regs_57_io_reset; // @[RegFile.scala 66:20:@125788.4]
  wire [63:0] regs_57_io_out; // @[RegFile.scala 66:20:@125788.4]
  wire  regs_57_io_enable; // @[RegFile.scala 66:20:@125788.4]
  wire  regs_58_clock; // @[RegFile.scala 66:20:@125802.4]
  wire  regs_58_reset; // @[RegFile.scala 66:20:@125802.4]
  wire [63:0] regs_58_io_in; // @[RegFile.scala 66:20:@125802.4]
  wire  regs_58_io_reset; // @[RegFile.scala 66:20:@125802.4]
  wire [63:0] regs_58_io_out; // @[RegFile.scala 66:20:@125802.4]
  wire  regs_58_io_enable; // @[RegFile.scala 66:20:@125802.4]
  wire  regs_59_clock; // @[RegFile.scala 66:20:@125816.4]
  wire  regs_59_reset; // @[RegFile.scala 66:20:@125816.4]
  wire [63:0] regs_59_io_in; // @[RegFile.scala 66:20:@125816.4]
  wire  regs_59_io_reset; // @[RegFile.scala 66:20:@125816.4]
  wire [63:0] regs_59_io_out; // @[RegFile.scala 66:20:@125816.4]
  wire  regs_59_io_enable; // @[RegFile.scala 66:20:@125816.4]
  wire  regs_60_clock; // @[RegFile.scala 66:20:@125830.4]
  wire  regs_60_reset; // @[RegFile.scala 66:20:@125830.4]
  wire [63:0] regs_60_io_in; // @[RegFile.scala 66:20:@125830.4]
  wire  regs_60_io_reset; // @[RegFile.scala 66:20:@125830.4]
  wire [63:0] regs_60_io_out; // @[RegFile.scala 66:20:@125830.4]
  wire  regs_60_io_enable; // @[RegFile.scala 66:20:@125830.4]
  wire  regs_61_clock; // @[RegFile.scala 66:20:@125844.4]
  wire  regs_61_reset; // @[RegFile.scala 66:20:@125844.4]
  wire [63:0] regs_61_io_in; // @[RegFile.scala 66:20:@125844.4]
  wire  regs_61_io_reset; // @[RegFile.scala 66:20:@125844.4]
  wire [63:0] regs_61_io_out; // @[RegFile.scala 66:20:@125844.4]
  wire  regs_61_io_enable; // @[RegFile.scala 66:20:@125844.4]
  wire  regs_62_clock; // @[RegFile.scala 66:20:@125858.4]
  wire  regs_62_reset; // @[RegFile.scala 66:20:@125858.4]
  wire [63:0] regs_62_io_in; // @[RegFile.scala 66:20:@125858.4]
  wire  regs_62_io_reset; // @[RegFile.scala 66:20:@125858.4]
  wire [63:0] regs_62_io_out; // @[RegFile.scala 66:20:@125858.4]
  wire  regs_62_io_enable; // @[RegFile.scala 66:20:@125858.4]
  wire  regs_63_clock; // @[RegFile.scala 66:20:@125872.4]
  wire  regs_63_reset; // @[RegFile.scala 66:20:@125872.4]
  wire [63:0] regs_63_io_in; // @[RegFile.scala 66:20:@125872.4]
  wire  regs_63_io_reset; // @[RegFile.scala 66:20:@125872.4]
  wire [63:0] regs_63_io_out; // @[RegFile.scala 66:20:@125872.4]
  wire  regs_63_io_enable; // @[RegFile.scala 66:20:@125872.4]
  wire  regs_64_clock; // @[RegFile.scala 66:20:@125886.4]
  wire  regs_64_reset; // @[RegFile.scala 66:20:@125886.4]
  wire [63:0] regs_64_io_in; // @[RegFile.scala 66:20:@125886.4]
  wire  regs_64_io_reset; // @[RegFile.scala 66:20:@125886.4]
  wire [63:0] regs_64_io_out; // @[RegFile.scala 66:20:@125886.4]
  wire  regs_64_io_enable; // @[RegFile.scala 66:20:@125886.4]
  wire  regs_65_clock; // @[RegFile.scala 66:20:@125900.4]
  wire  regs_65_reset; // @[RegFile.scala 66:20:@125900.4]
  wire [63:0] regs_65_io_in; // @[RegFile.scala 66:20:@125900.4]
  wire  regs_65_io_reset; // @[RegFile.scala 66:20:@125900.4]
  wire [63:0] regs_65_io_out; // @[RegFile.scala 66:20:@125900.4]
  wire  regs_65_io_enable; // @[RegFile.scala 66:20:@125900.4]
  wire  regs_66_clock; // @[RegFile.scala 66:20:@125914.4]
  wire  regs_66_reset; // @[RegFile.scala 66:20:@125914.4]
  wire [63:0] regs_66_io_in; // @[RegFile.scala 66:20:@125914.4]
  wire  regs_66_io_reset; // @[RegFile.scala 66:20:@125914.4]
  wire [63:0] regs_66_io_out; // @[RegFile.scala 66:20:@125914.4]
  wire  regs_66_io_enable; // @[RegFile.scala 66:20:@125914.4]
  wire  regs_67_clock; // @[RegFile.scala 66:20:@125928.4]
  wire  regs_67_reset; // @[RegFile.scala 66:20:@125928.4]
  wire [63:0] regs_67_io_in; // @[RegFile.scala 66:20:@125928.4]
  wire  regs_67_io_reset; // @[RegFile.scala 66:20:@125928.4]
  wire [63:0] regs_67_io_out; // @[RegFile.scala 66:20:@125928.4]
  wire  regs_67_io_enable; // @[RegFile.scala 66:20:@125928.4]
  wire  regs_68_clock; // @[RegFile.scala 66:20:@125942.4]
  wire  regs_68_reset; // @[RegFile.scala 66:20:@125942.4]
  wire [63:0] regs_68_io_in; // @[RegFile.scala 66:20:@125942.4]
  wire  regs_68_io_reset; // @[RegFile.scala 66:20:@125942.4]
  wire [63:0] regs_68_io_out; // @[RegFile.scala 66:20:@125942.4]
  wire  regs_68_io_enable; // @[RegFile.scala 66:20:@125942.4]
  wire  regs_69_clock; // @[RegFile.scala 66:20:@125956.4]
  wire  regs_69_reset; // @[RegFile.scala 66:20:@125956.4]
  wire [63:0] regs_69_io_in; // @[RegFile.scala 66:20:@125956.4]
  wire  regs_69_io_reset; // @[RegFile.scala 66:20:@125956.4]
  wire [63:0] regs_69_io_out; // @[RegFile.scala 66:20:@125956.4]
  wire  regs_69_io_enable; // @[RegFile.scala 66:20:@125956.4]
  wire  regs_70_clock; // @[RegFile.scala 66:20:@125970.4]
  wire  regs_70_reset; // @[RegFile.scala 66:20:@125970.4]
  wire [63:0] regs_70_io_in; // @[RegFile.scala 66:20:@125970.4]
  wire  regs_70_io_reset; // @[RegFile.scala 66:20:@125970.4]
  wire [63:0] regs_70_io_out; // @[RegFile.scala 66:20:@125970.4]
  wire  regs_70_io_enable; // @[RegFile.scala 66:20:@125970.4]
  wire  regs_71_clock; // @[RegFile.scala 66:20:@125984.4]
  wire  regs_71_reset; // @[RegFile.scala 66:20:@125984.4]
  wire [63:0] regs_71_io_in; // @[RegFile.scala 66:20:@125984.4]
  wire  regs_71_io_reset; // @[RegFile.scala 66:20:@125984.4]
  wire [63:0] regs_71_io_out; // @[RegFile.scala 66:20:@125984.4]
  wire  regs_71_io_enable; // @[RegFile.scala 66:20:@125984.4]
  wire  regs_72_clock; // @[RegFile.scala 66:20:@125998.4]
  wire  regs_72_reset; // @[RegFile.scala 66:20:@125998.4]
  wire [63:0] regs_72_io_in; // @[RegFile.scala 66:20:@125998.4]
  wire  regs_72_io_reset; // @[RegFile.scala 66:20:@125998.4]
  wire [63:0] regs_72_io_out; // @[RegFile.scala 66:20:@125998.4]
  wire  regs_72_io_enable; // @[RegFile.scala 66:20:@125998.4]
  wire  regs_73_clock; // @[RegFile.scala 66:20:@126012.4]
  wire  regs_73_reset; // @[RegFile.scala 66:20:@126012.4]
  wire [63:0] regs_73_io_in; // @[RegFile.scala 66:20:@126012.4]
  wire  regs_73_io_reset; // @[RegFile.scala 66:20:@126012.4]
  wire [63:0] regs_73_io_out; // @[RegFile.scala 66:20:@126012.4]
  wire  regs_73_io_enable; // @[RegFile.scala 66:20:@126012.4]
  wire  regs_74_clock; // @[RegFile.scala 66:20:@126026.4]
  wire  regs_74_reset; // @[RegFile.scala 66:20:@126026.4]
  wire [63:0] regs_74_io_in; // @[RegFile.scala 66:20:@126026.4]
  wire  regs_74_io_reset; // @[RegFile.scala 66:20:@126026.4]
  wire [63:0] regs_74_io_out; // @[RegFile.scala 66:20:@126026.4]
  wire  regs_74_io_enable; // @[RegFile.scala 66:20:@126026.4]
  wire  regs_75_clock; // @[RegFile.scala 66:20:@126040.4]
  wire  regs_75_reset; // @[RegFile.scala 66:20:@126040.4]
  wire [63:0] regs_75_io_in; // @[RegFile.scala 66:20:@126040.4]
  wire  regs_75_io_reset; // @[RegFile.scala 66:20:@126040.4]
  wire [63:0] regs_75_io_out; // @[RegFile.scala 66:20:@126040.4]
  wire  regs_75_io_enable; // @[RegFile.scala 66:20:@126040.4]
  wire  regs_76_clock; // @[RegFile.scala 66:20:@126054.4]
  wire  regs_76_reset; // @[RegFile.scala 66:20:@126054.4]
  wire [63:0] regs_76_io_in; // @[RegFile.scala 66:20:@126054.4]
  wire  regs_76_io_reset; // @[RegFile.scala 66:20:@126054.4]
  wire [63:0] regs_76_io_out; // @[RegFile.scala 66:20:@126054.4]
  wire  regs_76_io_enable; // @[RegFile.scala 66:20:@126054.4]
  wire  regs_77_clock; // @[RegFile.scala 66:20:@126068.4]
  wire  regs_77_reset; // @[RegFile.scala 66:20:@126068.4]
  wire [63:0] regs_77_io_in; // @[RegFile.scala 66:20:@126068.4]
  wire  regs_77_io_reset; // @[RegFile.scala 66:20:@126068.4]
  wire [63:0] regs_77_io_out; // @[RegFile.scala 66:20:@126068.4]
  wire  regs_77_io_enable; // @[RegFile.scala 66:20:@126068.4]
  wire  regs_78_clock; // @[RegFile.scala 66:20:@126082.4]
  wire  regs_78_reset; // @[RegFile.scala 66:20:@126082.4]
  wire [63:0] regs_78_io_in; // @[RegFile.scala 66:20:@126082.4]
  wire  regs_78_io_reset; // @[RegFile.scala 66:20:@126082.4]
  wire [63:0] regs_78_io_out; // @[RegFile.scala 66:20:@126082.4]
  wire  regs_78_io_enable; // @[RegFile.scala 66:20:@126082.4]
  wire  regs_79_clock; // @[RegFile.scala 66:20:@126096.4]
  wire  regs_79_reset; // @[RegFile.scala 66:20:@126096.4]
  wire [63:0] regs_79_io_in; // @[RegFile.scala 66:20:@126096.4]
  wire  regs_79_io_reset; // @[RegFile.scala 66:20:@126096.4]
  wire [63:0] regs_79_io_out; // @[RegFile.scala 66:20:@126096.4]
  wire  regs_79_io_enable; // @[RegFile.scala 66:20:@126096.4]
  wire  regs_80_clock; // @[RegFile.scala 66:20:@126110.4]
  wire  regs_80_reset; // @[RegFile.scala 66:20:@126110.4]
  wire [63:0] regs_80_io_in; // @[RegFile.scala 66:20:@126110.4]
  wire  regs_80_io_reset; // @[RegFile.scala 66:20:@126110.4]
  wire [63:0] regs_80_io_out; // @[RegFile.scala 66:20:@126110.4]
  wire  regs_80_io_enable; // @[RegFile.scala 66:20:@126110.4]
  wire  regs_81_clock; // @[RegFile.scala 66:20:@126124.4]
  wire  regs_81_reset; // @[RegFile.scala 66:20:@126124.4]
  wire [63:0] regs_81_io_in; // @[RegFile.scala 66:20:@126124.4]
  wire  regs_81_io_reset; // @[RegFile.scala 66:20:@126124.4]
  wire [63:0] regs_81_io_out; // @[RegFile.scala 66:20:@126124.4]
  wire  regs_81_io_enable; // @[RegFile.scala 66:20:@126124.4]
  wire  regs_82_clock; // @[RegFile.scala 66:20:@126138.4]
  wire  regs_82_reset; // @[RegFile.scala 66:20:@126138.4]
  wire [63:0] regs_82_io_in; // @[RegFile.scala 66:20:@126138.4]
  wire  regs_82_io_reset; // @[RegFile.scala 66:20:@126138.4]
  wire [63:0] regs_82_io_out; // @[RegFile.scala 66:20:@126138.4]
  wire  regs_82_io_enable; // @[RegFile.scala 66:20:@126138.4]
  wire  regs_83_clock; // @[RegFile.scala 66:20:@126152.4]
  wire  regs_83_reset; // @[RegFile.scala 66:20:@126152.4]
  wire [63:0] regs_83_io_in; // @[RegFile.scala 66:20:@126152.4]
  wire  regs_83_io_reset; // @[RegFile.scala 66:20:@126152.4]
  wire [63:0] regs_83_io_out; // @[RegFile.scala 66:20:@126152.4]
  wire  regs_83_io_enable; // @[RegFile.scala 66:20:@126152.4]
  wire  regs_84_clock; // @[RegFile.scala 66:20:@126166.4]
  wire  regs_84_reset; // @[RegFile.scala 66:20:@126166.4]
  wire [63:0] regs_84_io_in; // @[RegFile.scala 66:20:@126166.4]
  wire  regs_84_io_reset; // @[RegFile.scala 66:20:@126166.4]
  wire [63:0] regs_84_io_out; // @[RegFile.scala 66:20:@126166.4]
  wire  regs_84_io_enable; // @[RegFile.scala 66:20:@126166.4]
  wire  regs_85_clock; // @[RegFile.scala 66:20:@126180.4]
  wire  regs_85_reset; // @[RegFile.scala 66:20:@126180.4]
  wire [63:0] regs_85_io_in; // @[RegFile.scala 66:20:@126180.4]
  wire  regs_85_io_reset; // @[RegFile.scala 66:20:@126180.4]
  wire [63:0] regs_85_io_out; // @[RegFile.scala 66:20:@126180.4]
  wire  regs_85_io_enable; // @[RegFile.scala 66:20:@126180.4]
  wire  regs_86_clock; // @[RegFile.scala 66:20:@126194.4]
  wire  regs_86_reset; // @[RegFile.scala 66:20:@126194.4]
  wire [63:0] regs_86_io_in; // @[RegFile.scala 66:20:@126194.4]
  wire  regs_86_io_reset; // @[RegFile.scala 66:20:@126194.4]
  wire [63:0] regs_86_io_out; // @[RegFile.scala 66:20:@126194.4]
  wire  regs_86_io_enable; // @[RegFile.scala 66:20:@126194.4]
  wire  regs_87_clock; // @[RegFile.scala 66:20:@126208.4]
  wire  regs_87_reset; // @[RegFile.scala 66:20:@126208.4]
  wire [63:0] regs_87_io_in; // @[RegFile.scala 66:20:@126208.4]
  wire  regs_87_io_reset; // @[RegFile.scala 66:20:@126208.4]
  wire [63:0] regs_87_io_out; // @[RegFile.scala 66:20:@126208.4]
  wire  regs_87_io_enable; // @[RegFile.scala 66:20:@126208.4]
  wire  regs_88_clock; // @[RegFile.scala 66:20:@126222.4]
  wire  regs_88_reset; // @[RegFile.scala 66:20:@126222.4]
  wire [63:0] regs_88_io_in; // @[RegFile.scala 66:20:@126222.4]
  wire  regs_88_io_reset; // @[RegFile.scala 66:20:@126222.4]
  wire [63:0] regs_88_io_out; // @[RegFile.scala 66:20:@126222.4]
  wire  regs_88_io_enable; // @[RegFile.scala 66:20:@126222.4]
  wire  regs_89_clock; // @[RegFile.scala 66:20:@126236.4]
  wire  regs_89_reset; // @[RegFile.scala 66:20:@126236.4]
  wire [63:0] regs_89_io_in; // @[RegFile.scala 66:20:@126236.4]
  wire  regs_89_io_reset; // @[RegFile.scala 66:20:@126236.4]
  wire [63:0] regs_89_io_out; // @[RegFile.scala 66:20:@126236.4]
  wire  regs_89_io_enable; // @[RegFile.scala 66:20:@126236.4]
  wire  regs_90_clock; // @[RegFile.scala 66:20:@126250.4]
  wire  regs_90_reset; // @[RegFile.scala 66:20:@126250.4]
  wire [63:0] regs_90_io_in; // @[RegFile.scala 66:20:@126250.4]
  wire  regs_90_io_reset; // @[RegFile.scala 66:20:@126250.4]
  wire [63:0] regs_90_io_out; // @[RegFile.scala 66:20:@126250.4]
  wire  regs_90_io_enable; // @[RegFile.scala 66:20:@126250.4]
  wire  regs_91_clock; // @[RegFile.scala 66:20:@126264.4]
  wire  regs_91_reset; // @[RegFile.scala 66:20:@126264.4]
  wire [63:0] regs_91_io_in; // @[RegFile.scala 66:20:@126264.4]
  wire  regs_91_io_reset; // @[RegFile.scala 66:20:@126264.4]
  wire [63:0] regs_91_io_out; // @[RegFile.scala 66:20:@126264.4]
  wire  regs_91_io_enable; // @[RegFile.scala 66:20:@126264.4]
  wire  regs_92_clock; // @[RegFile.scala 66:20:@126278.4]
  wire  regs_92_reset; // @[RegFile.scala 66:20:@126278.4]
  wire [63:0] regs_92_io_in; // @[RegFile.scala 66:20:@126278.4]
  wire  regs_92_io_reset; // @[RegFile.scala 66:20:@126278.4]
  wire [63:0] regs_92_io_out; // @[RegFile.scala 66:20:@126278.4]
  wire  regs_92_io_enable; // @[RegFile.scala 66:20:@126278.4]
  wire  regs_93_clock; // @[RegFile.scala 66:20:@126292.4]
  wire  regs_93_reset; // @[RegFile.scala 66:20:@126292.4]
  wire [63:0] regs_93_io_in; // @[RegFile.scala 66:20:@126292.4]
  wire  regs_93_io_reset; // @[RegFile.scala 66:20:@126292.4]
  wire [63:0] regs_93_io_out; // @[RegFile.scala 66:20:@126292.4]
  wire  regs_93_io_enable; // @[RegFile.scala 66:20:@126292.4]
  wire  regs_94_clock; // @[RegFile.scala 66:20:@126306.4]
  wire  regs_94_reset; // @[RegFile.scala 66:20:@126306.4]
  wire [63:0] regs_94_io_in; // @[RegFile.scala 66:20:@126306.4]
  wire  regs_94_io_reset; // @[RegFile.scala 66:20:@126306.4]
  wire [63:0] regs_94_io_out; // @[RegFile.scala 66:20:@126306.4]
  wire  regs_94_io_enable; // @[RegFile.scala 66:20:@126306.4]
  wire  regs_95_clock; // @[RegFile.scala 66:20:@126320.4]
  wire  regs_95_reset; // @[RegFile.scala 66:20:@126320.4]
  wire [63:0] regs_95_io_in; // @[RegFile.scala 66:20:@126320.4]
  wire  regs_95_io_reset; // @[RegFile.scala 66:20:@126320.4]
  wire [63:0] regs_95_io_out; // @[RegFile.scala 66:20:@126320.4]
  wire  regs_95_io_enable; // @[RegFile.scala 66:20:@126320.4]
  wire  regs_96_clock; // @[RegFile.scala 66:20:@126334.4]
  wire  regs_96_reset; // @[RegFile.scala 66:20:@126334.4]
  wire [63:0] regs_96_io_in; // @[RegFile.scala 66:20:@126334.4]
  wire  regs_96_io_reset; // @[RegFile.scala 66:20:@126334.4]
  wire [63:0] regs_96_io_out; // @[RegFile.scala 66:20:@126334.4]
  wire  regs_96_io_enable; // @[RegFile.scala 66:20:@126334.4]
  wire  regs_97_clock; // @[RegFile.scala 66:20:@126348.4]
  wire  regs_97_reset; // @[RegFile.scala 66:20:@126348.4]
  wire [63:0] regs_97_io_in; // @[RegFile.scala 66:20:@126348.4]
  wire  regs_97_io_reset; // @[RegFile.scala 66:20:@126348.4]
  wire [63:0] regs_97_io_out; // @[RegFile.scala 66:20:@126348.4]
  wire  regs_97_io_enable; // @[RegFile.scala 66:20:@126348.4]
  wire  regs_98_clock; // @[RegFile.scala 66:20:@126362.4]
  wire  regs_98_reset; // @[RegFile.scala 66:20:@126362.4]
  wire [63:0] regs_98_io_in; // @[RegFile.scala 66:20:@126362.4]
  wire  regs_98_io_reset; // @[RegFile.scala 66:20:@126362.4]
  wire [63:0] regs_98_io_out; // @[RegFile.scala 66:20:@126362.4]
  wire  regs_98_io_enable; // @[RegFile.scala 66:20:@126362.4]
  wire  regs_99_clock; // @[RegFile.scala 66:20:@126376.4]
  wire  regs_99_reset; // @[RegFile.scala 66:20:@126376.4]
  wire [63:0] regs_99_io_in; // @[RegFile.scala 66:20:@126376.4]
  wire  regs_99_io_reset; // @[RegFile.scala 66:20:@126376.4]
  wire [63:0] regs_99_io_out; // @[RegFile.scala 66:20:@126376.4]
  wire  regs_99_io_enable; // @[RegFile.scala 66:20:@126376.4]
  wire  regs_100_clock; // @[RegFile.scala 66:20:@126390.4]
  wire  regs_100_reset; // @[RegFile.scala 66:20:@126390.4]
  wire [63:0] regs_100_io_in; // @[RegFile.scala 66:20:@126390.4]
  wire  regs_100_io_reset; // @[RegFile.scala 66:20:@126390.4]
  wire [63:0] regs_100_io_out; // @[RegFile.scala 66:20:@126390.4]
  wire  regs_100_io_enable; // @[RegFile.scala 66:20:@126390.4]
  wire  regs_101_clock; // @[RegFile.scala 66:20:@126404.4]
  wire  regs_101_reset; // @[RegFile.scala 66:20:@126404.4]
  wire [63:0] regs_101_io_in; // @[RegFile.scala 66:20:@126404.4]
  wire  regs_101_io_reset; // @[RegFile.scala 66:20:@126404.4]
  wire [63:0] regs_101_io_out; // @[RegFile.scala 66:20:@126404.4]
  wire  regs_101_io_enable; // @[RegFile.scala 66:20:@126404.4]
  wire  regs_102_clock; // @[RegFile.scala 66:20:@126418.4]
  wire  regs_102_reset; // @[RegFile.scala 66:20:@126418.4]
  wire [63:0] regs_102_io_in; // @[RegFile.scala 66:20:@126418.4]
  wire  regs_102_io_reset; // @[RegFile.scala 66:20:@126418.4]
  wire [63:0] regs_102_io_out; // @[RegFile.scala 66:20:@126418.4]
  wire  regs_102_io_enable; // @[RegFile.scala 66:20:@126418.4]
  wire  regs_103_clock; // @[RegFile.scala 66:20:@126432.4]
  wire  regs_103_reset; // @[RegFile.scala 66:20:@126432.4]
  wire [63:0] regs_103_io_in; // @[RegFile.scala 66:20:@126432.4]
  wire  regs_103_io_reset; // @[RegFile.scala 66:20:@126432.4]
  wire [63:0] regs_103_io_out; // @[RegFile.scala 66:20:@126432.4]
  wire  regs_103_io_enable; // @[RegFile.scala 66:20:@126432.4]
  wire  regs_104_clock; // @[RegFile.scala 66:20:@126446.4]
  wire  regs_104_reset; // @[RegFile.scala 66:20:@126446.4]
  wire [63:0] regs_104_io_in; // @[RegFile.scala 66:20:@126446.4]
  wire  regs_104_io_reset; // @[RegFile.scala 66:20:@126446.4]
  wire [63:0] regs_104_io_out; // @[RegFile.scala 66:20:@126446.4]
  wire  regs_104_io_enable; // @[RegFile.scala 66:20:@126446.4]
  wire  regs_105_clock; // @[RegFile.scala 66:20:@126460.4]
  wire  regs_105_reset; // @[RegFile.scala 66:20:@126460.4]
  wire [63:0] regs_105_io_in; // @[RegFile.scala 66:20:@126460.4]
  wire  regs_105_io_reset; // @[RegFile.scala 66:20:@126460.4]
  wire [63:0] regs_105_io_out; // @[RegFile.scala 66:20:@126460.4]
  wire  regs_105_io_enable; // @[RegFile.scala 66:20:@126460.4]
  wire  regs_106_clock; // @[RegFile.scala 66:20:@126474.4]
  wire  regs_106_reset; // @[RegFile.scala 66:20:@126474.4]
  wire [63:0] regs_106_io_in; // @[RegFile.scala 66:20:@126474.4]
  wire  regs_106_io_reset; // @[RegFile.scala 66:20:@126474.4]
  wire [63:0] regs_106_io_out; // @[RegFile.scala 66:20:@126474.4]
  wire  regs_106_io_enable; // @[RegFile.scala 66:20:@126474.4]
  wire  regs_107_clock; // @[RegFile.scala 66:20:@126488.4]
  wire  regs_107_reset; // @[RegFile.scala 66:20:@126488.4]
  wire [63:0] regs_107_io_in; // @[RegFile.scala 66:20:@126488.4]
  wire  regs_107_io_reset; // @[RegFile.scala 66:20:@126488.4]
  wire [63:0] regs_107_io_out; // @[RegFile.scala 66:20:@126488.4]
  wire  regs_107_io_enable; // @[RegFile.scala 66:20:@126488.4]
  wire  regs_108_clock; // @[RegFile.scala 66:20:@126502.4]
  wire  regs_108_reset; // @[RegFile.scala 66:20:@126502.4]
  wire [63:0] regs_108_io_in; // @[RegFile.scala 66:20:@126502.4]
  wire  regs_108_io_reset; // @[RegFile.scala 66:20:@126502.4]
  wire [63:0] regs_108_io_out; // @[RegFile.scala 66:20:@126502.4]
  wire  regs_108_io_enable; // @[RegFile.scala 66:20:@126502.4]
  wire  regs_109_clock; // @[RegFile.scala 66:20:@126516.4]
  wire  regs_109_reset; // @[RegFile.scala 66:20:@126516.4]
  wire [63:0] regs_109_io_in; // @[RegFile.scala 66:20:@126516.4]
  wire  regs_109_io_reset; // @[RegFile.scala 66:20:@126516.4]
  wire [63:0] regs_109_io_out; // @[RegFile.scala 66:20:@126516.4]
  wire  regs_109_io_enable; // @[RegFile.scala 66:20:@126516.4]
  wire  regs_110_clock; // @[RegFile.scala 66:20:@126530.4]
  wire  regs_110_reset; // @[RegFile.scala 66:20:@126530.4]
  wire [63:0] regs_110_io_in; // @[RegFile.scala 66:20:@126530.4]
  wire  regs_110_io_reset; // @[RegFile.scala 66:20:@126530.4]
  wire [63:0] regs_110_io_out; // @[RegFile.scala 66:20:@126530.4]
  wire  regs_110_io_enable; // @[RegFile.scala 66:20:@126530.4]
  wire  regs_111_clock; // @[RegFile.scala 66:20:@126544.4]
  wire  regs_111_reset; // @[RegFile.scala 66:20:@126544.4]
  wire [63:0] regs_111_io_in; // @[RegFile.scala 66:20:@126544.4]
  wire  regs_111_io_reset; // @[RegFile.scala 66:20:@126544.4]
  wire [63:0] regs_111_io_out; // @[RegFile.scala 66:20:@126544.4]
  wire  regs_111_io_enable; // @[RegFile.scala 66:20:@126544.4]
  wire  regs_112_clock; // @[RegFile.scala 66:20:@126558.4]
  wire  regs_112_reset; // @[RegFile.scala 66:20:@126558.4]
  wire [63:0] regs_112_io_in; // @[RegFile.scala 66:20:@126558.4]
  wire  regs_112_io_reset; // @[RegFile.scala 66:20:@126558.4]
  wire [63:0] regs_112_io_out; // @[RegFile.scala 66:20:@126558.4]
  wire  regs_112_io_enable; // @[RegFile.scala 66:20:@126558.4]
  wire  regs_113_clock; // @[RegFile.scala 66:20:@126572.4]
  wire  regs_113_reset; // @[RegFile.scala 66:20:@126572.4]
  wire [63:0] regs_113_io_in; // @[RegFile.scala 66:20:@126572.4]
  wire  regs_113_io_reset; // @[RegFile.scala 66:20:@126572.4]
  wire [63:0] regs_113_io_out; // @[RegFile.scala 66:20:@126572.4]
  wire  regs_113_io_enable; // @[RegFile.scala 66:20:@126572.4]
  wire  regs_114_clock; // @[RegFile.scala 66:20:@126586.4]
  wire  regs_114_reset; // @[RegFile.scala 66:20:@126586.4]
  wire [63:0] regs_114_io_in; // @[RegFile.scala 66:20:@126586.4]
  wire  regs_114_io_reset; // @[RegFile.scala 66:20:@126586.4]
  wire [63:0] regs_114_io_out; // @[RegFile.scala 66:20:@126586.4]
  wire  regs_114_io_enable; // @[RegFile.scala 66:20:@126586.4]
  wire  regs_115_clock; // @[RegFile.scala 66:20:@126600.4]
  wire  regs_115_reset; // @[RegFile.scala 66:20:@126600.4]
  wire [63:0] regs_115_io_in; // @[RegFile.scala 66:20:@126600.4]
  wire  regs_115_io_reset; // @[RegFile.scala 66:20:@126600.4]
  wire [63:0] regs_115_io_out; // @[RegFile.scala 66:20:@126600.4]
  wire  regs_115_io_enable; // @[RegFile.scala 66:20:@126600.4]
  wire  regs_116_clock; // @[RegFile.scala 66:20:@126614.4]
  wire  regs_116_reset; // @[RegFile.scala 66:20:@126614.4]
  wire [63:0] regs_116_io_in; // @[RegFile.scala 66:20:@126614.4]
  wire  regs_116_io_reset; // @[RegFile.scala 66:20:@126614.4]
  wire [63:0] regs_116_io_out; // @[RegFile.scala 66:20:@126614.4]
  wire  regs_116_io_enable; // @[RegFile.scala 66:20:@126614.4]
  wire  regs_117_clock; // @[RegFile.scala 66:20:@126628.4]
  wire  regs_117_reset; // @[RegFile.scala 66:20:@126628.4]
  wire [63:0] regs_117_io_in; // @[RegFile.scala 66:20:@126628.4]
  wire  regs_117_io_reset; // @[RegFile.scala 66:20:@126628.4]
  wire [63:0] regs_117_io_out; // @[RegFile.scala 66:20:@126628.4]
  wire  regs_117_io_enable; // @[RegFile.scala 66:20:@126628.4]
  wire  regs_118_clock; // @[RegFile.scala 66:20:@126642.4]
  wire  regs_118_reset; // @[RegFile.scala 66:20:@126642.4]
  wire [63:0] regs_118_io_in; // @[RegFile.scala 66:20:@126642.4]
  wire  regs_118_io_reset; // @[RegFile.scala 66:20:@126642.4]
  wire [63:0] regs_118_io_out; // @[RegFile.scala 66:20:@126642.4]
  wire  regs_118_io_enable; // @[RegFile.scala 66:20:@126642.4]
  wire  regs_119_clock; // @[RegFile.scala 66:20:@126656.4]
  wire  regs_119_reset; // @[RegFile.scala 66:20:@126656.4]
  wire [63:0] regs_119_io_in; // @[RegFile.scala 66:20:@126656.4]
  wire  regs_119_io_reset; // @[RegFile.scala 66:20:@126656.4]
  wire [63:0] regs_119_io_out; // @[RegFile.scala 66:20:@126656.4]
  wire  regs_119_io_enable; // @[RegFile.scala 66:20:@126656.4]
  wire  regs_120_clock; // @[RegFile.scala 66:20:@126670.4]
  wire  regs_120_reset; // @[RegFile.scala 66:20:@126670.4]
  wire [63:0] regs_120_io_in; // @[RegFile.scala 66:20:@126670.4]
  wire  regs_120_io_reset; // @[RegFile.scala 66:20:@126670.4]
  wire [63:0] regs_120_io_out; // @[RegFile.scala 66:20:@126670.4]
  wire  regs_120_io_enable; // @[RegFile.scala 66:20:@126670.4]
  wire  regs_121_clock; // @[RegFile.scala 66:20:@126684.4]
  wire  regs_121_reset; // @[RegFile.scala 66:20:@126684.4]
  wire [63:0] regs_121_io_in; // @[RegFile.scala 66:20:@126684.4]
  wire  regs_121_io_reset; // @[RegFile.scala 66:20:@126684.4]
  wire [63:0] regs_121_io_out; // @[RegFile.scala 66:20:@126684.4]
  wire  regs_121_io_enable; // @[RegFile.scala 66:20:@126684.4]
  wire  regs_122_clock; // @[RegFile.scala 66:20:@126698.4]
  wire  regs_122_reset; // @[RegFile.scala 66:20:@126698.4]
  wire [63:0] regs_122_io_in; // @[RegFile.scala 66:20:@126698.4]
  wire  regs_122_io_reset; // @[RegFile.scala 66:20:@126698.4]
  wire [63:0] regs_122_io_out; // @[RegFile.scala 66:20:@126698.4]
  wire  regs_122_io_enable; // @[RegFile.scala 66:20:@126698.4]
  wire  regs_123_clock; // @[RegFile.scala 66:20:@126712.4]
  wire  regs_123_reset; // @[RegFile.scala 66:20:@126712.4]
  wire [63:0] regs_123_io_in; // @[RegFile.scala 66:20:@126712.4]
  wire  regs_123_io_reset; // @[RegFile.scala 66:20:@126712.4]
  wire [63:0] regs_123_io_out; // @[RegFile.scala 66:20:@126712.4]
  wire  regs_123_io_enable; // @[RegFile.scala 66:20:@126712.4]
  wire  regs_124_clock; // @[RegFile.scala 66:20:@126726.4]
  wire  regs_124_reset; // @[RegFile.scala 66:20:@126726.4]
  wire [63:0] regs_124_io_in; // @[RegFile.scala 66:20:@126726.4]
  wire  regs_124_io_reset; // @[RegFile.scala 66:20:@126726.4]
  wire [63:0] regs_124_io_out; // @[RegFile.scala 66:20:@126726.4]
  wire  regs_124_io_enable; // @[RegFile.scala 66:20:@126726.4]
  wire  regs_125_clock; // @[RegFile.scala 66:20:@126740.4]
  wire  regs_125_reset; // @[RegFile.scala 66:20:@126740.4]
  wire [63:0] regs_125_io_in; // @[RegFile.scala 66:20:@126740.4]
  wire  regs_125_io_reset; // @[RegFile.scala 66:20:@126740.4]
  wire [63:0] regs_125_io_out; // @[RegFile.scala 66:20:@126740.4]
  wire  regs_125_io_enable; // @[RegFile.scala 66:20:@126740.4]
  wire  regs_126_clock; // @[RegFile.scala 66:20:@126754.4]
  wire  regs_126_reset; // @[RegFile.scala 66:20:@126754.4]
  wire [63:0] regs_126_io_in; // @[RegFile.scala 66:20:@126754.4]
  wire  regs_126_io_reset; // @[RegFile.scala 66:20:@126754.4]
  wire [63:0] regs_126_io_out; // @[RegFile.scala 66:20:@126754.4]
  wire  regs_126_io_enable; // @[RegFile.scala 66:20:@126754.4]
  wire  regs_127_clock; // @[RegFile.scala 66:20:@126768.4]
  wire  regs_127_reset; // @[RegFile.scala 66:20:@126768.4]
  wire [63:0] regs_127_io_in; // @[RegFile.scala 66:20:@126768.4]
  wire  regs_127_io_reset; // @[RegFile.scala 66:20:@126768.4]
  wire [63:0] regs_127_io_out; // @[RegFile.scala 66:20:@126768.4]
  wire  regs_127_io_enable; // @[RegFile.scala 66:20:@126768.4]
  wire  regs_128_clock; // @[RegFile.scala 66:20:@126782.4]
  wire  regs_128_reset; // @[RegFile.scala 66:20:@126782.4]
  wire [63:0] regs_128_io_in; // @[RegFile.scala 66:20:@126782.4]
  wire  regs_128_io_reset; // @[RegFile.scala 66:20:@126782.4]
  wire [63:0] regs_128_io_out; // @[RegFile.scala 66:20:@126782.4]
  wire  regs_128_io_enable; // @[RegFile.scala 66:20:@126782.4]
  wire  regs_129_clock; // @[RegFile.scala 66:20:@126796.4]
  wire  regs_129_reset; // @[RegFile.scala 66:20:@126796.4]
  wire [63:0] regs_129_io_in; // @[RegFile.scala 66:20:@126796.4]
  wire  regs_129_io_reset; // @[RegFile.scala 66:20:@126796.4]
  wire [63:0] regs_129_io_out; // @[RegFile.scala 66:20:@126796.4]
  wire  regs_129_io_enable; // @[RegFile.scala 66:20:@126796.4]
  wire  regs_130_clock; // @[RegFile.scala 66:20:@126810.4]
  wire  regs_130_reset; // @[RegFile.scala 66:20:@126810.4]
  wire [63:0] regs_130_io_in; // @[RegFile.scala 66:20:@126810.4]
  wire  regs_130_io_reset; // @[RegFile.scala 66:20:@126810.4]
  wire [63:0] regs_130_io_out; // @[RegFile.scala 66:20:@126810.4]
  wire  regs_130_io_enable; // @[RegFile.scala 66:20:@126810.4]
  wire  regs_131_clock; // @[RegFile.scala 66:20:@126824.4]
  wire  regs_131_reset; // @[RegFile.scala 66:20:@126824.4]
  wire [63:0] regs_131_io_in; // @[RegFile.scala 66:20:@126824.4]
  wire  regs_131_io_reset; // @[RegFile.scala 66:20:@126824.4]
  wire [63:0] regs_131_io_out; // @[RegFile.scala 66:20:@126824.4]
  wire  regs_131_io_enable; // @[RegFile.scala 66:20:@126824.4]
  wire  regs_132_clock; // @[RegFile.scala 66:20:@126838.4]
  wire  regs_132_reset; // @[RegFile.scala 66:20:@126838.4]
  wire [63:0] regs_132_io_in; // @[RegFile.scala 66:20:@126838.4]
  wire  regs_132_io_reset; // @[RegFile.scala 66:20:@126838.4]
  wire [63:0] regs_132_io_out; // @[RegFile.scala 66:20:@126838.4]
  wire  regs_132_io_enable; // @[RegFile.scala 66:20:@126838.4]
  wire  regs_133_clock; // @[RegFile.scala 66:20:@126852.4]
  wire  regs_133_reset; // @[RegFile.scala 66:20:@126852.4]
  wire [63:0] regs_133_io_in; // @[RegFile.scala 66:20:@126852.4]
  wire  regs_133_io_reset; // @[RegFile.scala 66:20:@126852.4]
  wire [63:0] regs_133_io_out; // @[RegFile.scala 66:20:@126852.4]
  wire  regs_133_io_enable; // @[RegFile.scala 66:20:@126852.4]
  wire  regs_134_clock; // @[RegFile.scala 66:20:@126866.4]
  wire  regs_134_reset; // @[RegFile.scala 66:20:@126866.4]
  wire [63:0] regs_134_io_in; // @[RegFile.scala 66:20:@126866.4]
  wire  regs_134_io_reset; // @[RegFile.scala 66:20:@126866.4]
  wire [63:0] regs_134_io_out; // @[RegFile.scala 66:20:@126866.4]
  wire  regs_134_io_enable; // @[RegFile.scala 66:20:@126866.4]
  wire  regs_135_clock; // @[RegFile.scala 66:20:@126880.4]
  wire  regs_135_reset; // @[RegFile.scala 66:20:@126880.4]
  wire [63:0] regs_135_io_in; // @[RegFile.scala 66:20:@126880.4]
  wire  regs_135_io_reset; // @[RegFile.scala 66:20:@126880.4]
  wire [63:0] regs_135_io_out; // @[RegFile.scala 66:20:@126880.4]
  wire  regs_135_io_enable; // @[RegFile.scala 66:20:@126880.4]
  wire  regs_136_clock; // @[RegFile.scala 66:20:@126894.4]
  wire  regs_136_reset; // @[RegFile.scala 66:20:@126894.4]
  wire [63:0] regs_136_io_in; // @[RegFile.scala 66:20:@126894.4]
  wire  regs_136_io_reset; // @[RegFile.scala 66:20:@126894.4]
  wire [63:0] regs_136_io_out; // @[RegFile.scala 66:20:@126894.4]
  wire  regs_136_io_enable; // @[RegFile.scala 66:20:@126894.4]
  wire  regs_137_clock; // @[RegFile.scala 66:20:@126908.4]
  wire  regs_137_reset; // @[RegFile.scala 66:20:@126908.4]
  wire [63:0] regs_137_io_in; // @[RegFile.scala 66:20:@126908.4]
  wire  regs_137_io_reset; // @[RegFile.scala 66:20:@126908.4]
  wire [63:0] regs_137_io_out; // @[RegFile.scala 66:20:@126908.4]
  wire  regs_137_io_enable; // @[RegFile.scala 66:20:@126908.4]
  wire  regs_138_clock; // @[RegFile.scala 66:20:@126922.4]
  wire  regs_138_reset; // @[RegFile.scala 66:20:@126922.4]
  wire [63:0] regs_138_io_in; // @[RegFile.scala 66:20:@126922.4]
  wire  regs_138_io_reset; // @[RegFile.scala 66:20:@126922.4]
  wire [63:0] regs_138_io_out; // @[RegFile.scala 66:20:@126922.4]
  wire  regs_138_io_enable; // @[RegFile.scala 66:20:@126922.4]
  wire  regs_139_clock; // @[RegFile.scala 66:20:@126936.4]
  wire  regs_139_reset; // @[RegFile.scala 66:20:@126936.4]
  wire [63:0] regs_139_io_in; // @[RegFile.scala 66:20:@126936.4]
  wire  regs_139_io_reset; // @[RegFile.scala 66:20:@126936.4]
  wire [63:0] regs_139_io_out; // @[RegFile.scala 66:20:@126936.4]
  wire  regs_139_io_enable; // @[RegFile.scala 66:20:@126936.4]
  wire  regs_140_clock; // @[RegFile.scala 66:20:@126950.4]
  wire  regs_140_reset; // @[RegFile.scala 66:20:@126950.4]
  wire [63:0] regs_140_io_in; // @[RegFile.scala 66:20:@126950.4]
  wire  regs_140_io_reset; // @[RegFile.scala 66:20:@126950.4]
  wire [63:0] regs_140_io_out; // @[RegFile.scala 66:20:@126950.4]
  wire  regs_140_io_enable; // @[RegFile.scala 66:20:@126950.4]
  wire  regs_141_clock; // @[RegFile.scala 66:20:@126964.4]
  wire  regs_141_reset; // @[RegFile.scala 66:20:@126964.4]
  wire [63:0] regs_141_io_in; // @[RegFile.scala 66:20:@126964.4]
  wire  regs_141_io_reset; // @[RegFile.scala 66:20:@126964.4]
  wire [63:0] regs_141_io_out; // @[RegFile.scala 66:20:@126964.4]
  wire  regs_141_io_enable; // @[RegFile.scala 66:20:@126964.4]
  wire  regs_142_clock; // @[RegFile.scala 66:20:@126978.4]
  wire  regs_142_reset; // @[RegFile.scala 66:20:@126978.4]
  wire [63:0] regs_142_io_in; // @[RegFile.scala 66:20:@126978.4]
  wire  regs_142_io_reset; // @[RegFile.scala 66:20:@126978.4]
  wire [63:0] regs_142_io_out; // @[RegFile.scala 66:20:@126978.4]
  wire  regs_142_io_enable; // @[RegFile.scala 66:20:@126978.4]
  wire  regs_143_clock; // @[RegFile.scala 66:20:@126992.4]
  wire  regs_143_reset; // @[RegFile.scala 66:20:@126992.4]
  wire [63:0] regs_143_io_in; // @[RegFile.scala 66:20:@126992.4]
  wire  regs_143_io_reset; // @[RegFile.scala 66:20:@126992.4]
  wire [63:0] regs_143_io_out; // @[RegFile.scala 66:20:@126992.4]
  wire  regs_143_io_enable; // @[RegFile.scala 66:20:@126992.4]
  wire  regs_144_clock; // @[RegFile.scala 66:20:@127006.4]
  wire  regs_144_reset; // @[RegFile.scala 66:20:@127006.4]
  wire [63:0] regs_144_io_in; // @[RegFile.scala 66:20:@127006.4]
  wire  regs_144_io_reset; // @[RegFile.scala 66:20:@127006.4]
  wire [63:0] regs_144_io_out; // @[RegFile.scala 66:20:@127006.4]
  wire  regs_144_io_enable; // @[RegFile.scala 66:20:@127006.4]
  wire  regs_145_clock; // @[RegFile.scala 66:20:@127020.4]
  wire  regs_145_reset; // @[RegFile.scala 66:20:@127020.4]
  wire [63:0] regs_145_io_in; // @[RegFile.scala 66:20:@127020.4]
  wire  regs_145_io_reset; // @[RegFile.scala 66:20:@127020.4]
  wire [63:0] regs_145_io_out; // @[RegFile.scala 66:20:@127020.4]
  wire  regs_145_io_enable; // @[RegFile.scala 66:20:@127020.4]
  wire  regs_146_clock; // @[RegFile.scala 66:20:@127034.4]
  wire  regs_146_reset; // @[RegFile.scala 66:20:@127034.4]
  wire [63:0] regs_146_io_in; // @[RegFile.scala 66:20:@127034.4]
  wire  regs_146_io_reset; // @[RegFile.scala 66:20:@127034.4]
  wire [63:0] regs_146_io_out; // @[RegFile.scala 66:20:@127034.4]
  wire  regs_146_io_enable; // @[RegFile.scala 66:20:@127034.4]
  wire  regs_147_clock; // @[RegFile.scala 66:20:@127048.4]
  wire  regs_147_reset; // @[RegFile.scala 66:20:@127048.4]
  wire [63:0] regs_147_io_in; // @[RegFile.scala 66:20:@127048.4]
  wire  regs_147_io_reset; // @[RegFile.scala 66:20:@127048.4]
  wire [63:0] regs_147_io_out; // @[RegFile.scala 66:20:@127048.4]
  wire  regs_147_io_enable; // @[RegFile.scala 66:20:@127048.4]
  wire  regs_148_clock; // @[RegFile.scala 66:20:@127062.4]
  wire  regs_148_reset; // @[RegFile.scala 66:20:@127062.4]
  wire [63:0] regs_148_io_in; // @[RegFile.scala 66:20:@127062.4]
  wire  regs_148_io_reset; // @[RegFile.scala 66:20:@127062.4]
  wire [63:0] regs_148_io_out; // @[RegFile.scala 66:20:@127062.4]
  wire  regs_148_io_enable; // @[RegFile.scala 66:20:@127062.4]
  wire  regs_149_clock; // @[RegFile.scala 66:20:@127076.4]
  wire  regs_149_reset; // @[RegFile.scala 66:20:@127076.4]
  wire [63:0] regs_149_io_in; // @[RegFile.scala 66:20:@127076.4]
  wire  regs_149_io_reset; // @[RegFile.scala 66:20:@127076.4]
  wire [63:0] regs_149_io_out; // @[RegFile.scala 66:20:@127076.4]
  wire  regs_149_io_enable; // @[RegFile.scala 66:20:@127076.4]
  wire  regs_150_clock; // @[RegFile.scala 66:20:@127090.4]
  wire  regs_150_reset; // @[RegFile.scala 66:20:@127090.4]
  wire [63:0] regs_150_io_in; // @[RegFile.scala 66:20:@127090.4]
  wire  regs_150_io_reset; // @[RegFile.scala 66:20:@127090.4]
  wire [63:0] regs_150_io_out; // @[RegFile.scala 66:20:@127090.4]
  wire  regs_150_io_enable; // @[RegFile.scala 66:20:@127090.4]
  wire  regs_151_clock; // @[RegFile.scala 66:20:@127104.4]
  wire  regs_151_reset; // @[RegFile.scala 66:20:@127104.4]
  wire [63:0] regs_151_io_in; // @[RegFile.scala 66:20:@127104.4]
  wire  regs_151_io_reset; // @[RegFile.scala 66:20:@127104.4]
  wire [63:0] regs_151_io_out; // @[RegFile.scala 66:20:@127104.4]
  wire  regs_151_io_enable; // @[RegFile.scala 66:20:@127104.4]
  wire  regs_152_clock; // @[RegFile.scala 66:20:@127118.4]
  wire  regs_152_reset; // @[RegFile.scala 66:20:@127118.4]
  wire [63:0] regs_152_io_in; // @[RegFile.scala 66:20:@127118.4]
  wire  regs_152_io_reset; // @[RegFile.scala 66:20:@127118.4]
  wire [63:0] regs_152_io_out; // @[RegFile.scala 66:20:@127118.4]
  wire  regs_152_io_enable; // @[RegFile.scala 66:20:@127118.4]
  wire  regs_153_clock; // @[RegFile.scala 66:20:@127132.4]
  wire  regs_153_reset; // @[RegFile.scala 66:20:@127132.4]
  wire [63:0] regs_153_io_in; // @[RegFile.scala 66:20:@127132.4]
  wire  regs_153_io_reset; // @[RegFile.scala 66:20:@127132.4]
  wire [63:0] regs_153_io_out; // @[RegFile.scala 66:20:@127132.4]
  wire  regs_153_io_enable; // @[RegFile.scala 66:20:@127132.4]
  wire  regs_154_clock; // @[RegFile.scala 66:20:@127146.4]
  wire  regs_154_reset; // @[RegFile.scala 66:20:@127146.4]
  wire [63:0] regs_154_io_in; // @[RegFile.scala 66:20:@127146.4]
  wire  regs_154_io_reset; // @[RegFile.scala 66:20:@127146.4]
  wire [63:0] regs_154_io_out; // @[RegFile.scala 66:20:@127146.4]
  wire  regs_154_io_enable; // @[RegFile.scala 66:20:@127146.4]
  wire  regs_155_clock; // @[RegFile.scala 66:20:@127160.4]
  wire  regs_155_reset; // @[RegFile.scala 66:20:@127160.4]
  wire [63:0] regs_155_io_in; // @[RegFile.scala 66:20:@127160.4]
  wire  regs_155_io_reset; // @[RegFile.scala 66:20:@127160.4]
  wire [63:0] regs_155_io_out; // @[RegFile.scala 66:20:@127160.4]
  wire  regs_155_io_enable; // @[RegFile.scala 66:20:@127160.4]
  wire  regs_156_clock; // @[RegFile.scala 66:20:@127174.4]
  wire  regs_156_reset; // @[RegFile.scala 66:20:@127174.4]
  wire [63:0] regs_156_io_in; // @[RegFile.scala 66:20:@127174.4]
  wire  regs_156_io_reset; // @[RegFile.scala 66:20:@127174.4]
  wire [63:0] regs_156_io_out; // @[RegFile.scala 66:20:@127174.4]
  wire  regs_156_io_enable; // @[RegFile.scala 66:20:@127174.4]
  wire  regs_157_clock; // @[RegFile.scala 66:20:@127188.4]
  wire  regs_157_reset; // @[RegFile.scala 66:20:@127188.4]
  wire [63:0] regs_157_io_in; // @[RegFile.scala 66:20:@127188.4]
  wire  regs_157_io_reset; // @[RegFile.scala 66:20:@127188.4]
  wire [63:0] regs_157_io_out; // @[RegFile.scala 66:20:@127188.4]
  wire  regs_157_io_enable; // @[RegFile.scala 66:20:@127188.4]
  wire  regs_158_clock; // @[RegFile.scala 66:20:@127202.4]
  wire  regs_158_reset; // @[RegFile.scala 66:20:@127202.4]
  wire [63:0] regs_158_io_in; // @[RegFile.scala 66:20:@127202.4]
  wire  regs_158_io_reset; // @[RegFile.scala 66:20:@127202.4]
  wire [63:0] regs_158_io_out; // @[RegFile.scala 66:20:@127202.4]
  wire  regs_158_io_enable; // @[RegFile.scala 66:20:@127202.4]
  wire  regs_159_clock; // @[RegFile.scala 66:20:@127216.4]
  wire  regs_159_reset; // @[RegFile.scala 66:20:@127216.4]
  wire [63:0] regs_159_io_in; // @[RegFile.scala 66:20:@127216.4]
  wire  regs_159_io_reset; // @[RegFile.scala 66:20:@127216.4]
  wire [63:0] regs_159_io_out; // @[RegFile.scala 66:20:@127216.4]
  wire  regs_159_io_enable; // @[RegFile.scala 66:20:@127216.4]
  wire  regs_160_clock; // @[RegFile.scala 66:20:@127230.4]
  wire  regs_160_reset; // @[RegFile.scala 66:20:@127230.4]
  wire [63:0] regs_160_io_in; // @[RegFile.scala 66:20:@127230.4]
  wire  regs_160_io_reset; // @[RegFile.scala 66:20:@127230.4]
  wire [63:0] regs_160_io_out; // @[RegFile.scala 66:20:@127230.4]
  wire  regs_160_io_enable; // @[RegFile.scala 66:20:@127230.4]
  wire  regs_161_clock; // @[RegFile.scala 66:20:@127244.4]
  wire  regs_161_reset; // @[RegFile.scala 66:20:@127244.4]
  wire [63:0] regs_161_io_in; // @[RegFile.scala 66:20:@127244.4]
  wire  regs_161_io_reset; // @[RegFile.scala 66:20:@127244.4]
  wire [63:0] regs_161_io_out; // @[RegFile.scala 66:20:@127244.4]
  wire  regs_161_io_enable; // @[RegFile.scala 66:20:@127244.4]
  wire  regs_162_clock; // @[RegFile.scala 66:20:@127258.4]
  wire  regs_162_reset; // @[RegFile.scala 66:20:@127258.4]
  wire [63:0] regs_162_io_in; // @[RegFile.scala 66:20:@127258.4]
  wire  regs_162_io_reset; // @[RegFile.scala 66:20:@127258.4]
  wire [63:0] regs_162_io_out; // @[RegFile.scala 66:20:@127258.4]
  wire  regs_162_io_enable; // @[RegFile.scala 66:20:@127258.4]
  wire  regs_163_clock; // @[RegFile.scala 66:20:@127272.4]
  wire  regs_163_reset; // @[RegFile.scala 66:20:@127272.4]
  wire [63:0] regs_163_io_in; // @[RegFile.scala 66:20:@127272.4]
  wire  regs_163_io_reset; // @[RegFile.scala 66:20:@127272.4]
  wire [63:0] regs_163_io_out; // @[RegFile.scala 66:20:@127272.4]
  wire  regs_163_io_enable; // @[RegFile.scala 66:20:@127272.4]
  wire  regs_164_clock; // @[RegFile.scala 66:20:@127286.4]
  wire  regs_164_reset; // @[RegFile.scala 66:20:@127286.4]
  wire [63:0] regs_164_io_in; // @[RegFile.scala 66:20:@127286.4]
  wire  regs_164_io_reset; // @[RegFile.scala 66:20:@127286.4]
  wire [63:0] regs_164_io_out; // @[RegFile.scala 66:20:@127286.4]
  wire  regs_164_io_enable; // @[RegFile.scala 66:20:@127286.4]
  wire  regs_165_clock; // @[RegFile.scala 66:20:@127300.4]
  wire  regs_165_reset; // @[RegFile.scala 66:20:@127300.4]
  wire [63:0] regs_165_io_in; // @[RegFile.scala 66:20:@127300.4]
  wire  regs_165_io_reset; // @[RegFile.scala 66:20:@127300.4]
  wire [63:0] regs_165_io_out; // @[RegFile.scala 66:20:@127300.4]
  wire  regs_165_io_enable; // @[RegFile.scala 66:20:@127300.4]
  wire  regs_166_clock; // @[RegFile.scala 66:20:@127314.4]
  wire  regs_166_reset; // @[RegFile.scala 66:20:@127314.4]
  wire [63:0] regs_166_io_in; // @[RegFile.scala 66:20:@127314.4]
  wire  regs_166_io_reset; // @[RegFile.scala 66:20:@127314.4]
  wire [63:0] regs_166_io_out; // @[RegFile.scala 66:20:@127314.4]
  wire  regs_166_io_enable; // @[RegFile.scala 66:20:@127314.4]
  wire  regs_167_clock; // @[RegFile.scala 66:20:@127328.4]
  wire  regs_167_reset; // @[RegFile.scala 66:20:@127328.4]
  wire [63:0] regs_167_io_in; // @[RegFile.scala 66:20:@127328.4]
  wire  regs_167_io_reset; // @[RegFile.scala 66:20:@127328.4]
  wire [63:0] regs_167_io_out; // @[RegFile.scala 66:20:@127328.4]
  wire  regs_167_io_enable; // @[RegFile.scala 66:20:@127328.4]
  wire  regs_168_clock; // @[RegFile.scala 66:20:@127342.4]
  wire  regs_168_reset; // @[RegFile.scala 66:20:@127342.4]
  wire [63:0] regs_168_io_in; // @[RegFile.scala 66:20:@127342.4]
  wire  regs_168_io_reset; // @[RegFile.scala 66:20:@127342.4]
  wire [63:0] regs_168_io_out; // @[RegFile.scala 66:20:@127342.4]
  wire  regs_168_io_enable; // @[RegFile.scala 66:20:@127342.4]
  wire  regs_169_clock; // @[RegFile.scala 66:20:@127356.4]
  wire  regs_169_reset; // @[RegFile.scala 66:20:@127356.4]
  wire [63:0] regs_169_io_in; // @[RegFile.scala 66:20:@127356.4]
  wire  regs_169_io_reset; // @[RegFile.scala 66:20:@127356.4]
  wire [63:0] regs_169_io_out; // @[RegFile.scala 66:20:@127356.4]
  wire  regs_169_io_enable; // @[RegFile.scala 66:20:@127356.4]
  wire  regs_170_clock; // @[RegFile.scala 66:20:@127370.4]
  wire  regs_170_reset; // @[RegFile.scala 66:20:@127370.4]
  wire [63:0] regs_170_io_in; // @[RegFile.scala 66:20:@127370.4]
  wire  regs_170_io_reset; // @[RegFile.scala 66:20:@127370.4]
  wire [63:0] regs_170_io_out; // @[RegFile.scala 66:20:@127370.4]
  wire  regs_170_io_enable; // @[RegFile.scala 66:20:@127370.4]
  wire  regs_171_clock; // @[RegFile.scala 66:20:@127384.4]
  wire  regs_171_reset; // @[RegFile.scala 66:20:@127384.4]
  wire [63:0] regs_171_io_in; // @[RegFile.scala 66:20:@127384.4]
  wire  regs_171_io_reset; // @[RegFile.scala 66:20:@127384.4]
  wire [63:0] regs_171_io_out; // @[RegFile.scala 66:20:@127384.4]
  wire  regs_171_io_enable; // @[RegFile.scala 66:20:@127384.4]
  wire  regs_172_clock; // @[RegFile.scala 66:20:@127398.4]
  wire  regs_172_reset; // @[RegFile.scala 66:20:@127398.4]
  wire [63:0] regs_172_io_in; // @[RegFile.scala 66:20:@127398.4]
  wire  regs_172_io_reset; // @[RegFile.scala 66:20:@127398.4]
  wire [63:0] regs_172_io_out; // @[RegFile.scala 66:20:@127398.4]
  wire  regs_172_io_enable; // @[RegFile.scala 66:20:@127398.4]
  wire  regs_173_clock; // @[RegFile.scala 66:20:@127412.4]
  wire  regs_173_reset; // @[RegFile.scala 66:20:@127412.4]
  wire [63:0] regs_173_io_in; // @[RegFile.scala 66:20:@127412.4]
  wire  regs_173_io_reset; // @[RegFile.scala 66:20:@127412.4]
  wire [63:0] regs_173_io_out; // @[RegFile.scala 66:20:@127412.4]
  wire  regs_173_io_enable; // @[RegFile.scala 66:20:@127412.4]
  wire  regs_174_clock; // @[RegFile.scala 66:20:@127426.4]
  wire  regs_174_reset; // @[RegFile.scala 66:20:@127426.4]
  wire [63:0] regs_174_io_in; // @[RegFile.scala 66:20:@127426.4]
  wire  regs_174_io_reset; // @[RegFile.scala 66:20:@127426.4]
  wire [63:0] regs_174_io_out; // @[RegFile.scala 66:20:@127426.4]
  wire  regs_174_io_enable; // @[RegFile.scala 66:20:@127426.4]
  wire  regs_175_clock; // @[RegFile.scala 66:20:@127440.4]
  wire  regs_175_reset; // @[RegFile.scala 66:20:@127440.4]
  wire [63:0] regs_175_io_in; // @[RegFile.scala 66:20:@127440.4]
  wire  regs_175_io_reset; // @[RegFile.scala 66:20:@127440.4]
  wire [63:0] regs_175_io_out; // @[RegFile.scala 66:20:@127440.4]
  wire  regs_175_io_enable; // @[RegFile.scala 66:20:@127440.4]
  wire  regs_176_clock; // @[RegFile.scala 66:20:@127454.4]
  wire  regs_176_reset; // @[RegFile.scala 66:20:@127454.4]
  wire [63:0] regs_176_io_in; // @[RegFile.scala 66:20:@127454.4]
  wire  regs_176_io_reset; // @[RegFile.scala 66:20:@127454.4]
  wire [63:0] regs_176_io_out; // @[RegFile.scala 66:20:@127454.4]
  wire  regs_176_io_enable; // @[RegFile.scala 66:20:@127454.4]
  wire  regs_177_clock; // @[RegFile.scala 66:20:@127468.4]
  wire  regs_177_reset; // @[RegFile.scala 66:20:@127468.4]
  wire [63:0] regs_177_io_in; // @[RegFile.scala 66:20:@127468.4]
  wire  regs_177_io_reset; // @[RegFile.scala 66:20:@127468.4]
  wire [63:0] regs_177_io_out; // @[RegFile.scala 66:20:@127468.4]
  wire  regs_177_io_enable; // @[RegFile.scala 66:20:@127468.4]
  wire  regs_178_clock; // @[RegFile.scala 66:20:@127482.4]
  wire  regs_178_reset; // @[RegFile.scala 66:20:@127482.4]
  wire [63:0] regs_178_io_in; // @[RegFile.scala 66:20:@127482.4]
  wire  regs_178_io_reset; // @[RegFile.scala 66:20:@127482.4]
  wire [63:0] regs_178_io_out; // @[RegFile.scala 66:20:@127482.4]
  wire  regs_178_io_enable; // @[RegFile.scala 66:20:@127482.4]
  wire  regs_179_clock; // @[RegFile.scala 66:20:@127496.4]
  wire  regs_179_reset; // @[RegFile.scala 66:20:@127496.4]
  wire [63:0] regs_179_io_in; // @[RegFile.scala 66:20:@127496.4]
  wire  regs_179_io_reset; // @[RegFile.scala 66:20:@127496.4]
  wire [63:0] regs_179_io_out; // @[RegFile.scala 66:20:@127496.4]
  wire  regs_179_io_enable; // @[RegFile.scala 66:20:@127496.4]
  wire  regs_180_clock; // @[RegFile.scala 66:20:@127510.4]
  wire  regs_180_reset; // @[RegFile.scala 66:20:@127510.4]
  wire [63:0] regs_180_io_in; // @[RegFile.scala 66:20:@127510.4]
  wire  regs_180_io_reset; // @[RegFile.scala 66:20:@127510.4]
  wire [63:0] regs_180_io_out; // @[RegFile.scala 66:20:@127510.4]
  wire  regs_180_io_enable; // @[RegFile.scala 66:20:@127510.4]
  wire  regs_181_clock; // @[RegFile.scala 66:20:@127524.4]
  wire  regs_181_reset; // @[RegFile.scala 66:20:@127524.4]
  wire [63:0] regs_181_io_in; // @[RegFile.scala 66:20:@127524.4]
  wire  regs_181_io_reset; // @[RegFile.scala 66:20:@127524.4]
  wire [63:0] regs_181_io_out; // @[RegFile.scala 66:20:@127524.4]
  wire  regs_181_io_enable; // @[RegFile.scala 66:20:@127524.4]
  wire  regs_182_clock; // @[RegFile.scala 66:20:@127538.4]
  wire  regs_182_reset; // @[RegFile.scala 66:20:@127538.4]
  wire [63:0] regs_182_io_in; // @[RegFile.scala 66:20:@127538.4]
  wire  regs_182_io_reset; // @[RegFile.scala 66:20:@127538.4]
  wire [63:0] regs_182_io_out; // @[RegFile.scala 66:20:@127538.4]
  wire  regs_182_io_enable; // @[RegFile.scala 66:20:@127538.4]
  wire  regs_183_clock; // @[RegFile.scala 66:20:@127552.4]
  wire  regs_183_reset; // @[RegFile.scala 66:20:@127552.4]
  wire [63:0] regs_183_io_in; // @[RegFile.scala 66:20:@127552.4]
  wire  regs_183_io_reset; // @[RegFile.scala 66:20:@127552.4]
  wire [63:0] regs_183_io_out; // @[RegFile.scala 66:20:@127552.4]
  wire  regs_183_io_enable; // @[RegFile.scala 66:20:@127552.4]
  wire  regs_184_clock; // @[RegFile.scala 66:20:@127566.4]
  wire  regs_184_reset; // @[RegFile.scala 66:20:@127566.4]
  wire [63:0] regs_184_io_in; // @[RegFile.scala 66:20:@127566.4]
  wire  regs_184_io_reset; // @[RegFile.scala 66:20:@127566.4]
  wire [63:0] regs_184_io_out; // @[RegFile.scala 66:20:@127566.4]
  wire  regs_184_io_enable; // @[RegFile.scala 66:20:@127566.4]
  wire  regs_185_clock; // @[RegFile.scala 66:20:@127580.4]
  wire  regs_185_reset; // @[RegFile.scala 66:20:@127580.4]
  wire [63:0] regs_185_io_in; // @[RegFile.scala 66:20:@127580.4]
  wire  regs_185_io_reset; // @[RegFile.scala 66:20:@127580.4]
  wire [63:0] regs_185_io_out; // @[RegFile.scala 66:20:@127580.4]
  wire  regs_185_io_enable; // @[RegFile.scala 66:20:@127580.4]
  wire  regs_186_clock; // @[RegFile.scala 66:20:@127594.4]
  wire  regs_186_reset; // @[RegFile.scala 66:20:@127594.4]
  wire [63:0] regs_186_io_in; // @[RegFile.scala 66:20:@127594.4]
  wire  regs_186_io_reset; // @[RegFile.scala 66:20:@127594.4]
  wire [63:0] regs_186_io_out; // @[RegFile.scala 66:20:@127594.4]
  wire  regs_186_io_enable; // @[RegFile.scala 66:20:@127594.4]
  wire  regs_187_clock; // @[RegFile.scala 66:20:@127608.4]
  wire  regs_187_reset; // @[RegFile.scala 66:20:@127608.4]
  wire [63:0] regs_187_io_in; // @[RegFile.scala 66:20:@127608.4]
  wire  regs_187_io_reset; // @[RegFile.scala 66:20:@127608.4]
  wire [63:0] regs_187_io_out; // @[RegFile.scala 66:20:@127608.4]
  wire  regs_187_io_enable; // @[RegFile.scala 66:20:@127608.4]
  wire  regs_188_clock; // @[RegFile.scala 66:20:@127622.4]
  wire  regs_188_reset; // @[RegFile.scala 66:20:@127622.4]
  wire [63:0] regs_188_io_in; // @[RegFile.scala 66:20:@127622.4]
  wire  regs_188_io_reset; // @[RegFile.scala 66:20:@127622.4]
  wire [63:0] regs_188_io_out; // @[RegFile.scala 66:20:@127622.4]
  wire  regs_188_io_enable; // @[RegFile.scala 66:20:@127622.4]
  wire  regs_189_clock; // @[RegFile.scala 66:20:@127636.4]
  wire  regs_189_reset; // @[RegFile.scala 66:20:@127636.4]
  wire [63:0] regs_189_io_in; // @[RegFile.scala 66:20:@127636.4]
  wire  regs_189_io_reset; // @[RegFile.scala 66:20:@127636.4]
  wire [63:0] regs_189_io_out; // @[RegFile.scala 66:20:@127636.4]
  wire  regs_189_io_enable; // @[RegFile.scala 66:20:@127636.4]
  wire  regs_190_clock; // @[RegFile.scala 66:20:@127650.4]
  wire  regs_190_reset; // @[RegFile.scala 66:20:@127650.4]
  wire [63:0] regs_190_io_in; // @[RegFile.scala 66:20:@127650.4]
  wire  regs_190_io_reset; // @[RegFile.scala 66:20:@127650.4]
  wire [63:0] regs_190_io_out; // @[RegFile.scala 66:20:@127650.4]
  wire  regs_190_io_enable; // @[RegFile.scala 66:20:@127650.4]
  wire  regs_191_clock; // @[RegFile.scala 66:20:@127664.4]
  wire  regs_191_reset; // @[RegFile.scala 66:20:@127664.4]
  wire [63:0] regs_191_io_in; // @[RegFile.scala 66:20:@127664.4]
  wire  regs_191_io_reset; // @[RegFile.scala 66:20:@127664.4]
  wire [63:0] regs_191_io_out; // @[RegFile.scala 66:20:@127664.4]
  wire  regs_191_io_enable; // @[RegFile.scala 66:20:@127664.4]
  wire  regs_192_clock; // @[RegFile.scala 66:20:@127678.4]
  wire  regs_192_reset; // @[RegFile.scala 66:20:@127678.4]
  wire [63:0] regs_192_io_in; // @[RegFile.scala 66:20:@127678.4]
  wire  regs_192_io_reset; // @[RegFile.scala 66:20:@127678.4]
  wire [63:0] regs_192_io_out; // @[RegFile.scala 66:20:@127678.4]
  wire  regs_192_io_enable; // @[RegFile.scala 66:20:@127678.4]
  wire  regs_193_clock; // @[RegFile.scala 66:20:@127692.4]
  wire  regs_193_reset; // @[RegFile.scala 66:20:@127692.4]
  wire [63:0] regs_193_io_in; // @[RegFile.scala 66:20:@127692.4]
  wire  regs_193_io_reset; // @[RegFile.scala 66:20:@127692.4]
  wire [63:0] regs_193_io_out; // @[RegFile.scala 66:20:@127692.4]
  wire  regs_193_io_enable; // @[RegFile.scala 66:20:@127692.4]
  wire  regs_194_clock; // @[RegFile.scala 66:20:@127706.4]
  wire  regs_194_reset; // @[RegFile.scala 66:20:@127706.4]
  wire [63:0] regs_194_io_in; // @[RegFile.scala 66:20:@127706.4]
  wire  regs_194_io_reset; // @[RegFile.scala 66:20:@127706.4]
  wire [63:0] regs_194_io_out; // @[RegFile.scala 66:20:@127706.4]
  wire  regs_194_io_enable; // @[RegFile.scala 66:20:@127706.4]
  wire  regs_195_clock; // @[RegFile.scala 66:20:@127720.4]
  wire  regs_195_reset; // @[RegFile.scala 66:20:@127720.4]
  wire [63:0] regs_195_io_in; // @[RegFile.scala 66:20:@127720.4]
  wire  regs_195_io_reset; // @[RegFile.scala 66:20:@127720.4]
  wire [63:0] regs_195_io_out; // @[RegFile.scala 66:20:@127720.4]
  wire  regs_195_io_enable; // @[RegFile.scala 66:20:@127720.4]
  wire  regs_196_clock; // @[RegFile.scala 66:20:@127734.4]
  wire  regs_196_reset; // @[RegFile.scala 66:20:@127734.4]
  wire [63:0] regs_196_io_in; // @[RegFile.scala 66:20:@127734.4]
  wire  regs_196_io_reset; // @[RegFile.scala 66:20:@127734.4]
  wire [63:0] regs_196_io_out; // @[RegFile.scala 66:20:@127734.4]
  wire  regs_196_io_enable; // @[RegFile.scala 66:20:@127734.4]
  wire  regs_197_clock; // @[RegFile.scala 66:20:@127748.4]
  wire  regs_197_reset; // @[RegFile.scala 66:20:@127748.4]
  wire [63:0] regs_197_io_in; // @[RegFile.scala 66:20:@127748.4]
  wire  regs_197_io_reset; // @[RegFile.scala 66:20:@127748.4]
  wire [63:0] regs_197_io_out; // @[RegFile.scala 66:20:@127748.4]
  wire  regs_197_io_enable; // @[RegFile.scala 66:20:@127748.4]
  wire  regs_198_clock; // @[RegFile.scala 66:20:@127762.4]
  wire  regs_198_reset; // @[RegFile.scala 66:20:@127762.4]
  wire [63:0] regs_198_io_in; // @[RegFile.scala 66:20:@127762.4]
  wire  regs_198_io_reset; // @[RegFile.scala 66:20:@127762.4]
  wire [63:0] regs_198_io_out; // @[RegFile.scala 66:20:@127762.4]
  wire  regs_198_io_enable; // @[RegFile.scala 66:20:@127762.4]
  wire  regs_199_clock; // @[RegFile.scala 66:20:@127776.4]
  wire  regs_199_reset; // @[RegFile.scala 66:20:@127776.4]
  wire [63:0] regs_199_io_in; // @[RegFile.scala 66:20:@127776.4]
  wire  regs_199_io_reset; // @[RegFile.scala 66:20:@127776.4]
  wire [63:0] regs_199_io_out; // @[RegFile.scala 66:20:@127776.4]
  wire  regs_199_io_enable; // @[RegFile.scala 66:20:@127776.4]
  wire  regs_200_clock; // @[RegFile.scala 66:20:@127790.4]
  wire  regs_200_reset; // @[RegFile.scala 66:20:@127790.4]
  wire [63:0] regs_200_io_in; // @[RegFile.scala 66:20:@127790.4]
  wire  regs_200_io_reset; // @[RegFile.scala 66:20:@127790.4]
  wire [63:0] regs_200_io_out; // @[RegFile.scala 66:20:@127790.4]
  wire  regs_200_io_enable; // @[RegFile.scala 66:20:@127790.4]
  wire  regs_201_clock; // @[RegFile.scala 66:20:@127804.4]
  wire  regs_201_reset; // @[RegFile.scala 66:20:@127804.4]
  wire [63:0] regs_201_io_in; // @[RegFile.scala 66:20:@127804.4]
  wire  regs_201_io_reset; // @[RegFile.scala 66:20:@127804.4]
  wire [63:0] regs_201_io_out; // @[RegFile.scala 66:20:@127804.4]
  wire  regs_201_io_enable; // @[RegFile.scala 66:20:@127804.4]
  wire  regs_202_clock; // @[RegFile.scala 66:20:@127818.4]
  wire  regs_202_reset; // @[RegFile.scala 66:20:@127818.4]
  wire [63:0] regs_202_io_in; // @[RegFile.scala 66:20:@127818.4]
  wire  regs_202_io_reset; // @[RegFile.scala 66:20:@127818.4]
  wire [63:0] regs_202_io_out; // @[RegFile.scala 66:20:@127818.4]
  wire  regs_202_io_enable; // @[RegFile.scala 66:20:@127818.4]
  wire  regs_203_clock; // @[RegFile.scala 66:20:@127832.4]
  wire  regs_203_reset; // @[RegFile.scala 66:20:@127832.4]
  wire [63:0] regs_203_io_in; // @[RegFile.scala 66:20:@127832.4]
  wire  regs_203_io_reset; // @[RegFile.scala 66:20:@127832.4]
  wire [63:0] regs_203_io_out; // @[RegFile.scala 66:20:@127832.4]
  wire  regs_203_io_enable; // @[RegFile.scala 66:20:@127832.4]
  wire  regs_204_clock; // @[RegFile.scala 66:20:@127846.4]
  wire  regs_204_reset; // @[RegFile.scala 66:20:@127846.4]
  wire [63:0] regs_204_io_in; // @[RegFile.scala 66:20:@127846.4]
  wire  regs_204_io_reset; // @[RegFile.scala 66:20:@127846.4]
  wire [63:0] regs_204_io_out; // @[RegFile.scala 66:20:@127846.4]
  wire  regs_204_io_enable; // @[RegFile.scala 66:20:@127846.4]
  wire  regs_205_clock; // @[RegFile.scala 66:20:@127860.4]
  wire  regs_205_reset; // @[RegFile.scala 66:20:@127860.4]
  wire [63:0] regs_205_io_in; // @[RegFile.scala 66:20:@127860.4]
  wire  regs_205_io_reset; // @[RegFile.scala 66:20:@127860.4]
  wire [63:0] regs_205_io_out; // @[RegFile.scala 66:20:@127860.4]
  wire  regs_205_io_enable; // @[RegFile.scala 66:20:@127860.4]
  wire  regs_206_clock; // @[RegFile.scala 66:20:@127874.4]
  wire  regs_206_reset; // @[RegFile.scala 66:20:@127874.4]
  wire [63:0] regs_206_io_in; // @[RegFile.scala 66:20:@127874.4]
  wire  regs_206_io_reset; // @[RegFile.scala 66:20:@127874.4]
  wire [63:0] regs_206_io_out; // @[RegFile.scala 66:20:@127874.4]
  wire  regs_206_io_enable; // @[RegFile.scala 66:20:@127874.4]
  wire  regs_207_clock; // @[RegFile.scala 66:20:@127888.4]
  wire  regs_207_reset; // @[RegFile.scala 66:20:@127888.4]
  wire [63:0] regs_207_io_in; // @[RegFile.scala 66:20:@127888.4]
  wire  regs_207_io_reset; // @[RegFile.scala 66:20:@127888.4]
  wire [63:0] regs_207_io_out; // @[RegFile.scala 66:20:@127888.4]
  wire  regs_207_io_enable; // @[RegFile.scala 66:20:@127888.4]
  wire  regs_208_clock; // @[RegFile.scala 66:20:@127902.4]
  wire  regs_208_reset; // @[RegFile.scala 66:20:@127902.4]
  wire [63:0] regs_208_io_in; // @[RegFile.scala 66:20:@127902.4]
  wire  regs_208_io_reset; // @[RegFile.scala 66:20:@127902.4]
  wire [63:0] regs_208_io_out; // @[RegFile.scala 66:20:@127902.4]
  wire  regs_208_io_enable; // @[RegFile.scala 66:20:@127902.4]
  wire  regs_209_clock; // @[RegFile.scala 66:20:@127916.4]
  wire  regs_209_reset; // @[RegFile.scala 66:20:@127916.4]
  wire [63:0] regs_209_io_in; // @[RegFile.scala 66:20:@127916.4]
  wire  regs_209_io_reset; // @[RegFile.scala 66:20:@127916.4]
  wire [63:0] regs_209_io_out; // @[RegFile.scala 66:20:@127916.4]
  wire  regs_209_io_enable; // @[RegFile.scala 66:20:@127916.4]
  wire  regs_210_clock; // @[RegFile.scala 66:20:@127930.4]
  wire  regs_210_reset; // @[RegFile.scala 66:20:@127930.4]
  wire [63:0] regs_210_io_in; // @[RegFile.scala 66:20:@127930.4]
  wire  regs_210_io_reset; // @[RegFile.scala 66:20:@127930.4]
  wire [63:0] regs_210_io_out; // @[RegFile.scala 66:20:@127930.4]
  wire  regs_210_io_enable; // @[RegFile.scala 66:20:@127930.4]
  wire  regs_211_clock; // @[RegFile.scala 66:20:@127944.4]
  wire  regs_211_reset; // @[RegFile.scala 66:20:@127944.4]
  wire [63:0] regs_211_io_in; // @[RegFile.scala 66:20:@127944.4]
  wire  regs_211_io_reset; // @[RegFile.scala 66:20:@127944.4]
  wire [63:0] regs_211_io_out; // @[RegFile.scala 66:20:@127944.4]
  wire  regs_211_io_enable; // @[RegFile.scala 66:20:@127944.4]
  wire  regs_212_clock; // @[RegFile.scala 66:20:@127958.4]
  wire  regs_212_reset; // @[RegFile.scala 66:20:@127958.4]
  wire [63:0] regs_212_io_in; // @[RegFile.scala 66:20:@127958.4]
  wire  regs_212_io_reset; // @[RegFile.scala 66:20:@127958.4]
  wire [63:0] regs_212_io_out; // @[RegFile.scala 66:20:@127958.4]
  wire  regs_212_io_enable; // @[RegFile.scala 66:20:@127958.4]
  wire  regs_213_clock; // @[RegFile.scala 66:20:@127972.4]
  wire  regs_213_reset; // @[RegFile.scala 66:20:@127972.4]
  wire [63:0] regs_213_io_in; // @[RegFile.scala 66:20:@127972.4]
  wire  regs_213_io_reset; // @[RegFile.scala 66:20:@127972.4]
  wire [63:0] regs_213_io_out; // @[RegFile.scala 66:20:@127972.4]
  wire  regs_213_io_enable; // @[RegFile.scala 66:20:@127972.4]
  wire  regs_214_clock; // @[RegFile.scala 66:20:@127986.4]
  wire  regs_214_reset; // @[RegFile.scala 66:20:@127986.4]
  wire [63:0] regs_214_io_in; // @[RegFile.scala 66:20:@127986.4]
  wire  regs_214_io_reset; // @[RegFile.scala 66:20:@127986.4]
  wire [63:0] regs_214_io_out; // @[RegFile.scala 66:20:@127986.4]
  wire  regs_214_io_enable; // @[RegFile.scala 66:20:@127986.4]
  wire  regs_215_clock; // @[RegFile.scala 66:20:@128000.4]
  wire  regs_215_reset; // @[RegFile.scala 66:20:@128000.4]
  wire [63:0] regs_215_io_in; // @[RegFile.scala 66:20:@128000.4]
  wire  regs_215_io_reset; // @[RegFile.scala 66:20:@128000.4]
  wire [63:0] regs_215_io_out; // @[RegFile.scala 66:20:@128000.4]
  wire  regs_215_io_enable; // @[RegFile.scala 66:20:@128000.4]
  wire  regs_216_clock; // @[RegFile.scala 66:20:@128014.4]
  wire  regs_216_reset; // @[RegFile.scala 66:20:@128014.4]
  wire [63:0] regs_216_io_in; // @[RegFile.scala 66:20:@128014.4]
  wire  regs_216_io_reset; // @[RegFile.scala 66:20:@128014.4]
  wire [63:0] regs_216_io_out; // @[RegFile.scala 66:20:@128014.4]
  wire  regs_216_io_enable; // @[RegFile.scala 66:20:@128014.4]
  wire  regs_217_clock; // @[RegFile.scala 66:20:@128028.4]
  wire  regs_217_reset; // @[RegFile.scala 66:20:@128028.4]
  wire [63:0] regs_217_io_in; // @[RegFile.scala 66:20:@128028.4]
  wire  regs_217_io_reset; // @[RegFile.scala 66:20:@128028.4]
  wire [63:0] regs_217_io_out; // @[RegFile.scala 66:20:@128028.4]
  wire  regs_217_io_enable; // @[RegFile.scala 66:20:@128028.4]
  wire  regs_218_clock; // @[RegFile.scala 66:20:@128042.4]
  wire  regs_218_reset; // @[RegFile.scala 66:20:@128042.4]
  wire [63:0] regs_218_io_in; // @[RegFile.scala 66:20:@128042.4]
  wire  regs_218_io_reset; // @[RegFile.scala 66:20:@128042.4]
  wire [63:0] regs_218_io_out; // @[RegFile.scala 66:20:@128042.4]
  wire  regs_218_io_enable; // @[RegFile.scala 66:20:@128042.4]
  wire  regs_219_clock; // @[RegFile.scala 66:20:@128056.4]
  wire  regs_219_reset; // @[RegFile.scala 66:20:@128056.4]
  wire [63:0] regs_219_io_in; // @[RegFile.scala 66:20:@128056.4]
  wire  regs_219_io_reset; // @[RegFile.scala 66:20:@128056.4]
  wire [63:0] regs_219_io_out; // @[RegFile.scala 66:20:@128056.4]
  wire  regs_219_io_enable; // @[RegFile.scala 66:20:@128056.4]
  wire  regs_220_clock; // @[RegFile.scala 66:20:@128070.4]
  wire  regs_220_reset; // @[RegFile.scala 66:20:@128070.4]
  wire [63:0] regs_220_io_in; // @[RegFile.scala 66:20:@128070.4]
  wire  regs_220_io_reset; // @[RegFile.scala 66:20:@128070.4]
  wire [63:0] regs_220_io_out; // @[RegFile.scala 66:20:@128070.4]
  wire  regs_220_io_enable; // @[RegFile.scala 66:20:@128070.4]
  wire  regs_221_clock; // @[RegFile.scala 66:20:@128084.4]
  wire  regs_221_reset; // @[RegFile.scala 66:20:@128084.4]
  wire [63:0] regs_221_io_in; // @[RegFile.scala 66:20:@128084.4]
  wire  regs_221_io_reset; // @[RegFile.scala 66:20:@128084.4]
  wire [63:0] regs_221_io_out; // @[RegFile.scala 66:20:@128084.4]
  wire  regs_221_io_enable; // @[RegFile.scala 66:20:@128084.4]
  wire  regs_222_clock; // @[RegFile.scala 66:20:@128098.4]
  wire  regs_222_reset; // @[RegFile.scala 66:20:@128098.4]
  wire [63:0] regs_222_io_in; // @[RegFile.scala 66:20:@128098.4]
  wire  regs_222_io_reset; // @[RegFile.scala 66:20:@128098.4]
  wire [63:0] regs_222_io_out; // @[RegFile.scala 66:20:@128098.4]
  wire  regs_222_io_enable; // @[RegFile.scala 66:20:@128098.4]
  wire  regs_223_clock; // @[RegFile.scala 66:20:@128112.4]
  wire  regs_223_reset; // @[RegFile.scala 66:20:@128112.4]
  wire [63:0] regs_223_io_in; // @[RegFile.scala 66:20:@128112.4]
  wire  regs_223_io_reset; // @[RegFile.scala 66:20:@128112.4]
  wire [63:0] regs_223_io_out; // @[RegFile.scala 66:20:@128112.4]
  wire  regs_223_io_enable; // @[RegFile.scala 66:20:@128112.4]
  wire  regs_224_clock; // @[RegFile.scala 66:20:@128126.4]
  wire  regs_224_reset; // @[RegFile.scala 66:20:@128126.4]
  wire [63:0] regs_224_io_in; // @[RegFile.scala 66:20:@128126.4]
  wire  regs_224_io_reset; // @[RegFile.scala 66:20:@128126.4]
  wire [63:0] regs_224_io_out; // @[RegFile.scala 66:20:@128126.4]
  wire  regs_224_io_enable; // @[RegFile.scala 66:20:@128126.4]
  wire  regs_225_clock; // @[RegFile.scala 66:20:@128140.4]
  wire  regs_225_reset; // @[RegFile.scala 66:20:@128140.4]
  wire [63:0] regs_225_io_in; // @[RegFile.scala 66:20:@128140.4]
  wire  regs_225_io_reset; // @[RegFile.scala 66:20:@128140.4]
  wire [63:0] regs_225_io_out; // @[RegFile.scala 66:20:@128140.4]
  wire  regs_225_io_enable; // @[RegFile.scala 66:20:@128140.4]
  wire  regs_226_clock; // @[RegFile.scala 66:20:@128154.4]
  wire  regs_226_reset; // @[RegFile.scala 66:20:@128154.4]
  wire [63:0] regs_226_io_in; // @[RegFile.scala 66:20:@128154.4]
  wire  regs_226_io_reset; // @[RegFile.scala 66:20:@128154.4]
  wire [63:0] regs_226_io_out; // @[RegFile.scala 66:20:@128154.4]
  wire  regs_226_io_enable; // @[RegFile.scala 66:20:@128154.4]
  wire  regs_227_clock; // @[RegFile.scala 66:20:@128168.4]
  wire  regs_227_reset; // @[RegFile.scala 66:20:@128168.4]
  wire [63:0] regs_227_io_in; // @[RegFile.scala 66:20:@128168.4]
  wire  regs_227_io_reset; // @[RegFile.scala 66:20:@128168.4]
  wire [63:0] regs_227_io_out; // @[RegFile.scala 66:20:@128168.4]
  wire  regs_227_io_enable; // @[RegFile.scala 66:20:@128168.4]
  wire  regs_228_clock; // @[RegFile.scala 66:20:@128182.4]
  wire  regs_228_reset; // @[RegFile.scala 66:20:@128182.4]
  wire [63:0] regs_228_io_in; // @[RegFile.scala 66:20:@128182.4]
  wire  regs_228_io_reset; // @[RegFile.scala 66:20:@128182.4]
  wire [63:0] regs_228_io_out; // @[RegFile.scala 66:20:@128182.4]
  wire  regs_228_io_enable; // @[RegFile.scala 66:20:@128182.4]
  wire  regs_229_clock; // @[RegFile.scala 66:20:@128196.4]
  wire  regs_229_reset; // @[RegFile.scala 66:20:@128196.4]
  wire [63:0] regs_229_io_in; // @[RegFile.scala 66:20:@128196.4]
  wire  regs_229_io_reset; // @[RegFile.scala 66:20:@128196.4]
  wire [63:0] regs_229_io_out; // @[RegFile.scala 66:20:@128196.4]
  wire  regs_229_io_enable; // @[RegFile.scala 66:20:@128196.4]
  wire  regs_230_clock; // @[RegFile.scala 66:20:@128210.4]
  wire  regs_230_reset; // @[RegFile.scala 66:20:@128210.4]
  wire [63:0] regs_230_io_in; // @[RegFile.scala 66:20:@128210.4]
  wire  regs_230_io_reset; // @[RegFile.scala 66:20:@128210.4]
  wire [63:0] regs_230_io_out; // @[RegFile.scala 66:20:@128210.4]
  wire  regs_230_io_enable; // @[RegFile.scala 66:20:@128210.4]
  wire  regs_231_clock; // @[RegFile.scala 66:20:@128224.4]
  wire  regs_231_reset; // @[RegFile.scala 66:20:@128224.4]
  wire [63:0] regs_231_io_in; // @[RegFile.scala 66:20:@128224.4]
  wire  regs_231_io_reset; // @[RegFile.scala 66:20:@128224.4]
  wire [63:0] regs_231_io_out; // @[RegFile.scala 66:20:@128224.4]
  wire  regs_231_io_enable; // @[RegFile.scala 66:20:@128224.4]
  wire  regs_232_clock; // @[RegFile.scala 66:20:@128238.4]
  wire  regs_232_reset; // @[RegFile.scala 66:20:@128238.4]
  wire [63:0] regs_232_io_in; // @[RegFile.scala 66:20:@128238.4]
  wire  regs_232_io_reset; // @[RegFile.scala 66:20:@128238.4]
  wire [63:0] regs_232_io_out; // @[RegFile.scala 66:20:@128238.4]
  wire  regs_232_io_enable; // @[RegFile.scala 66:20:@128238.4]
  wire  regs_233_clock; // @[RegFile.scala 66:20:@128252.4]
  wire  regs_233_reset; // @[RegFile.scala 66:20:@128252.4]
  wire [63:0] regs_233_io_in; // @[RegFile.scala 66:20:@128252.4]
  wire  regs_233_io_reset; // @[RegFile.scala 66:20:@128252.4]
  wire [63:0] regs_233_io_out; // @[RegFile.scala 66:20:@128252.4]
  wire  regs_233_io_enable; // @[RegFile.scala 66:20:@128252.4]
  wire  regs_234_clock; // @[RegFile.scala 66:20:@128266.4]
  wire  regs_234_reset; // @[RegFile.scala 66:20:@128266.4]
  wire [63:0] regs_234_io_in; // @[RegFile.scala 66:20:@128266.4]
  wire  regs_234_io_reset; // @[RegFile.scala 66:20:@128266.4]
  wire [63:0] regs_234_io_out; // @[RegFile.scala 66:20:@128266.4]
  wire  regs_234_io_enable; // @[RegFile.scala 66:20:@128266.4]
  wire  regs_235_clock; // @[RegFile.scala 66:20:@128280.4]
  wire  regs_235_reset; // @[RegFile.scala 66:20:@128280.4]
  wire [63:0] regs_235_io_in; // @[RegFile.scala 66:20:@128280.4]
  wire  regs_235_io_reset; // @[RegFile.scala 66:20:@128280.4]
  wire [63:0] regs_235_io_out; // @[RegFile.scala 66:20:@128280.4]
  wire  regs_235_io_enable; // @[RegFile.scala 66:20:@128280.4]
  wire  regs_236_clock; // @[RegFile.scala 66:20:@128294.4]
  wire  regs_236_reset; // @[RegFile.scala 66:20:@128294.4]
  wire [63:0] regs_236_io_in; // @[RegFile.scala 66:20:@128294.4]
  wire  regs_236_io_reset; // @[RegFile.scala 66:20:@128294.4]
  wire [63:0] regs_236_io_out; // @[RegFile.scala 66:20:@128294.4]
  wire  regs_236_io_enable; // @[RegFile.scala 66:20:@128294.4]
  wire  regs_237_clock; // @[RegFile.scala 66:20:@128308.4]
  wire  regs_237_reset; // @[RegFile.scala 66:20:@128308.4]
  wire [63:0] regs_237_io_in; // @[RegFile.scala 66:20:@128308.4]
  wire  regs_237_io_reset; // @[RegFile.scala 66:20:@128308.4]
  wire [63:0] regs_237_io_out; // @[RegFile.scala 66:20:@128308.4]
  wire  regs_237_io_enable; // @[RegFile.scala 66:20:@128308.4]
  wire  regs_238_clock; // @[RegFile.scala 66:20:@128322.4]
  wire  regs_238_reset; // @[RegFile.scala 66:20:@128322.4]
  wire [63:0] regs_238_io_in; // @[RegFile.scala 66:20:@128322.4]
  wire  regs_238_io_reset; // @[RegFile.scala 66:20:@128322.4]
  wire [63:0] regs_238_io_out; // @[RegFile.scala 66:20:@128322.4]
  wire  regs_238_io_enable; // @[RegFile.scala 66:20:@128322.4]
  wire  regs_239_clock; // @[RegFile.scala 66:20:@128336.4]
  wire  regs_239_reset; // @[RegFile.scala 66:20:@128336.4]
  wire [63:0] regs_239_io_in; // @[RegFile.scala 66:20:@128336.4]
  wire  regs_239_io_reset; // @[RegFile.scala 66:20:@128336.4]
  wire [63:0] regs_239_io_out; // @[RegFile.scala 66:20:@128336.4]
  wire  regs_239_io_enable; // @[RegFile.scala 66:20:@128336.4]
  wire  regs_240_clock; // @[RegFile.scala 66:20:@128350.4]
  wire  regs_240_reset; // @[RegFile.scala 66:20:@128350.4]
  wire [63:0] regs_240_io_in; // @[RegFile.scala 66:20:@128350.4]
  wire  regs_240_io_reset; // @[RegFile.scala 66:20:@128350.4]
  wire [63:0] regs_240_io_out; // @[RegFile.scala 66:20:@128350.4]
  wire  regs_240_io_enable; // @[RegFile.scala 66:20:@128350.4]
  wire  regs_241_clock; // @[RegFile.scala 66:20:@128364.4]
  wire  regs_241_reset; // @[RegFile.scala 66:20:@128364.4]
  wire [63:0] regs_241_io_in; // @[RegFile.scala 66:20:@128364.4]
  wire  regs_241_io_reset; // @[RegFile.scala 66:20:@128364.4]
  wire [63:0] regs_241_io_out; // @[RegFile.scala 66:20:@128364.4]
  wire  regs_241_io_enable; // @[RegFile.scala 66:20:@128364.4]
  wire  regs_242_clock; // @[RegFile.scala 66:20:@128378.4]
  wire  regs_242_reset; // @[RegFile.scala 66:20:@128378.4]
  wire [63:0] regs_242_io_in; // @[RegFile.scala 66:20:@128378.4]
  wire  regs_242_io_reset; // @[RegFile.scala 66:20:@128378.4]
  wire [63:0] regs_242_io_out; // @[RegFile.scala 66:20:@128378.4]
  wire  regs_242_io_enable; // @[RegFile.scala 66:20:@128378.4]
  wire  regs_243_clock; // @[RegFile.scala 66:20:@128392.4]
  wire  regs_243_reset; // @[RegFile.scala 66:20:@128392.4]
  wire [63:0] regs_243_io_in; // @[RegFile.scala 66:20:@128392.4]
  wire  regs_243_io_reset; // @[RegFile.scala 66:20:@128392.4]
  wire [63:0] regs_243_io_out; // @[RegFile.scala 66:20:@128392.4]
  wire  regs_243_io_enable; // @[RegFile.scala 66:20:@128392.4]
  wire  regs_244_clock; // @[RegFile.scala 66:20:@128406.4]
  wire  regs_244_reset; // @[RegFile.scala 66:20:@128406.4]
  wire [63:0] regs_244_io_in; // @[RegFile.scala 66:20:@128406.4]
  wire  regs_244_io_reset; // @[RegFile.scala 66:20:@128406.4]
  wire [63:0] regs_244_io_out; // @[RegFile.scala 66:20:@128406.4]
  wire  regs_244_io_enable; // @[RegFile.scala 66:20:@128406.4]
  wire  regs_245_clock; // @[RegFile.scala 66:20:@128420.4]
  wire  regs_245_reset; // @[RegFile.scala 66:20:@128420.4]
  wire [63:0] regs_245_io_in; // @[RegFile.scala 66:20:@128420.4]
  wire  regs_245_io_reset; // @[RegFile.scala 66:20:@128420.4]
  wire [63:0] regs_245_io_out; // @[RegFile.scala 66:20:@128420.4]
  wire  regs_245_io_enable; // @[RegFile.scala 66:20:@128420.4]
  wire  regs_246_clock; // @[RegFile.scala 66:20:@128434.4]
  wire  regs_246_reset; // @[RegFile.scala 66:20:@128434.4]
  wire [63:0] regs_246_io_in; // @[RegFile.scala 66:20:@128434.4]
  wire  regs_246_io_reset; // @[RegFile.scala 66:20:@128434.4]
  wire [63:0] regs_246_io_out; // @[RegFile.scala 66:20:@128434.4]
  wire  regs_246_io_enable; // @[RegFile.scala 66:20:@128434.4]
  wire  regs_247_clock; // @[RegFile.scala 66:20:@128448.4]
  wire  regs_247_reset; // @[RegFile.scala 66:20:@128448.4]
  wire [63:0] regs_247_io_in; // @[RegFile.scala 66:20:@128448.4]
  wire  regs_247_io_reset; // @[RegFile.scala 66:20:@128448.4]
  wire [63:0] regs_247_io_out; // @[RegFile.scala 66:20:@128448.4]
  wire  regs_247_io_enable; // @[RegFile.scala 66:20:@128448.4]
  wire  regs_248_clock; // @[RegFile.scala 66:20:@128462.4]
  wire  regs_248_reset; // @[RegFile.scala 66:20:@128462.4]
  wire [63:0] regs_248_io_in; // @[RegFile.scala 66:20:@128462.4]
  wire  regs_248_io_reset; // @[RegFile.scala 66:20:@128462.4]
  wire [63:0] regs_248_io_out; // @[RegFile.scala 66:20:@128462.4]
  wire  regs_248_io_enable; // @[RegFile.scala 66:20:@128462.4]
  wire  regs_249_clock; // @[RegFile.scala 66:20:@128476.4]
  wire  regs_249_reset; // @[RegFile.scala 66:20:@128476.4]
  wire [63:0] regs_249_io_in; // @[RegFile.scala 66:20:@128476.4]
  wire  regs_249_io_reset; // @[RegFile.scala 66:20:@128476.4]
  wire [63:0] regs_249_io_out; // @[RegFile.scala 66:20:@128476.4]
  wire  regs_249_io_enable; // @[RegFile.scala 66:20:@128476.4]
  wire  regs_250_clock; // @[RegFile.scala 66:20:@128490.4]
  wire  regs_250_reset; // @[RegFile.scala 66:20:@128490.4]
  wire [63:0] regs_250_io_in; // @[RegFile.scala 66:20:@128490.4]
  wire  regs_250_io_reset; // @[RegFile.scala 66:20:@128490.4]
  wire [63:0] regs_250_io_out; // @[RegFile.scala 66:20:@128490.4]
  wire  regs_250_io_enable; // @[RegFile.scala 66:20:@128490.4]
  wire  regs_251_clock; // @[RegFile.scala 66:20:@128504.4]
  wire  regs_251_reset; // @[RegFile.scala 66:20:@128504.4]
  wire [63:0] regs_251_io_in; // @[RegFile.scala 66:20:@128504.4]
  wire  regs_251_io_reset; // @[RegFile.scala 66:20:@128504.4]
  wire [63:0] regs_251_io_out; // @[RegFile.scala 66:20:@128504.4]
  wire  regs_251_io_enable; // @[RegFile.scala 66:20:@128504.4]
  wire  regs_252_clock; // @[RegFile.scala 66:20:@128518.4]
  wire  regs_252_reset; // @[RegFile.scala 66:20:@128518.4]
  wire [63:0] regs_252_io_in; // @[RegFile.scala 66:20:@128518.4]
  wire  regs_252_io_reset; // @[RegFile.scala 66:20:@128518.4]
  wire [63:0] regs_252_io_out; // @[RegFile.scala 66:20:@128518.4]
  wire  regs_252_io_enable; // @[RegFile.scala 66:20:@128518.4]
  wire  regs_253_clock; // @[RegFile.scala 66:20:@128532.4]
  wire  regs_253_reset; // @[RegFile.scala 66:20:@128532.4]
  wire [63:0] regs_253_io_in; // @[RegFile.scala 66:20:@128532.4]
  wire  regs_253_io_reset; // @[RegFile.scala 66:20:@128532.4]
  wire [63:0] regs_253_io_out; // @[RegFile.scala 66:20:@128532.4]
  wire  regs_253_io_enable; // @[RegFile.scala 66:20:@128532.4]
  wire  regs_254_clock; // @[RegFile.scala 66:20:@128546.4]
  wire  regs_254_reset; // @[RegFile.scala 66:20:@128546.4]
  wire [63:0] regs_254_io_in; // @[RegFile.scala 66:20:@128546.4]
  wire  regs_254_io_reset; // @[RegFile.scala 66:20:@128546.4]
  wire [63:0] regs_254_io_out; // @[RegFile.scala 66:20:@128546.4]
  wire  regs_254_io_enable; // @[RegFile.scala 66:20:@128546.4]
  wire  regs_255_clock; // @[RegFile.scala 66:20:@128560.4]
  wire  regs_255_reset; // @[RegFile.scala 66:20:@128560.4]
  wire [63:0] regs_255_io_in; // @[RegFile.scala 66:20:@128560.4]
  wire  regs_255_io_reset; // @[RegFile.scala 66:20:@128560.4]
  wire [63:0] regs_255_io_out; // @[RegFile.scala 66:20:@128560.4]
  wire  regs_255_io_enable; // @[RegFile.scala 66:20:@128560.4]
  wire  regs_256_clock; // @[RegFile.scala 66:20:@128574.4]
  wire  regs_256_reset; // @[RegFile.scala 66:20:@128574.4]
  wire [63:0] regs_256_io_in; // @[RegFile.scala 66:20:@128574.4]
  wire  regs_256_io_reset; // @[RegFile.scala 66:20:@128574.4]
  wire [63:0] regs_256_io_out; // @[RegFile.scala 66:20:@128574.4]
  wire  regs_256_io_enable; // @[RegFile.scala 66:20:@128574.4]
  wire  regs_257_clock; // @[RegFile.scala 66:20:@128588.4]
  wire  regs_257_reset; // @[RegFile.scala 66:20:@128588.4]
  wire [63:0] regs_257_io_in; // @[RegFile.scala 66:20:@128588.4]
  wire  regs_257_io_reset; // @[RegFile.scala 66:20:@128588.4]
  wire [63:0] regs_257_io_out; // @[RegFile.scala 66:20:@128588.4]
  wire  regs_257_io_enable; // @[RegFile.scala 66:20:@128588.4]
  wire  regs_258_clock; // @[RegFile.scala 66:20:@128602.4]
  wire  regs_258_reset; // @[RegFile.scala 66:20:@128602.4]
  wire [63:0] regs_258_io_in; // @[RegFile.scala 66:20:@128602.4]
  wire  regs_258_io_reset; // @[RegFile.scala 66:20:@128602.4]
  wire [63:0] regs_258_io_out; // @[RegFile.scala 66:20:@128602.4]
  wire  regs_258_io_enable; // @[RegFile.scala 66:20:@128602.4]
  wire  regs_259_clock; // @[RegFile.scala 66:20:@128616.4]
  wire  regs_259_reset; // @[RegFile.scala 66:20:@128616.4]
  wire [63:0] regs_259_io_in; // @[RegFile.scala 66:20:@128616.4]
  wire  regs_259_io_reset; // @[RegFile.scala 66:20:@128616.4]
  wire [63:0] regs_259_io_out; // @[RegFile.scala 66:20:@128616.4]
  wire  regs_259_io_enable; // @[RegFile.scala 66:20:@128616.4]
  wire  regs_260_clock; // @[RegFile.scala 66:20:@128630.4]
  wire  regs_260_reset; // @[RegFile.scala 66:20:@128630.4]
  wire [63:0] regs_260_io_in; // @[RegFile.scala 66:20:@128630.4]
  wire  regs_260_io_reset; // @[RegFile.scala 66:20:@128630.4]
  wire [63:0] regs_260_io_out; // @[RegFile.scala 66:20:@128630.4]
  wire  regs_260_io_enable; // @[RegFile.scala 66:20:@128630.4]
  wire  regs_261_clock; // @[RegFile.scala 66:20:@128644.4]
  wire  regs_261_reset; // @[RegFile.scala 66:20:@128644.4]
  wire [63:0] regs_261_io_in; // @[RegFile.scala 66:20:@128644.4]
  wire  regs_261_io_reset; // @[RegFile.scala 66:20:@128644.4]
  wire [63:0] regs_261_io_out; // @[RegFile.scala 66:20:@128644.4]
  wire  regs_261_io_enable; // @[RegFile.scala 66:20:@128644.4]
  wire  regs_262_clock; // @[RegFile.scala 66:20:@128658.4]
  wire  regs_262_reset; // @[RegFile.scala 66:20:@128658.4]
  wire [63:0] regs_262_io_in; // @[RegFile.scala 66:20:@128658.4]
  wire  regs_262_io_reset; // @[RegFile.scala 66:20:@128658.4]
  wire [63:0] regs_262_io_out; // @[RegFile.scala 66:20:@128658.4]
  wire  regs_262_io_enable; // @[RegFile.scala 66:20:@128658.4]
  wire  regs_263_clock; // @[RegFile.scala 66:20:@128672.4]
  wire  regs_263_reset; // @[RegFile.scala 66:20:@128672.4]
  wire [63:0] regs_263_io_in; // @[RegFile.scala 66:20:@128672.4]
  wire  regs_263_io_reset; // @[RegFile.scala 66:20:@128672.4]
  wire [63:0] regs_263_io_out; // @[RegFile.scala 66:20:@128672.4]
  wire  regs_263_io_enable; // @[RegFile.scala 66:20:@128672.4]
  wire  regs_264_clock; // @[RegFile.scala 66:20:@128686.4]
  wire  regs_264_reset; // @[RegFile.scala 66:20:@128686.4]
  wire [63:0] regs_264_io_in; // @[RegFile.scala 66:20:@128686.4]
  wire  regs_264_io_reset; // @[RegFile.scala 66:20:@128686.4]
  wire [63:0] regs_264_io_out; // @[RegFile.scala 66:20:@128686.4]
  wire  regs_264_io_enable; // @[RegFile.scala 66:20:@128686.4]
  wire  regs_265_clock; // @[RegFile.scala 66:20:@128700.4]
  wire  regs_265_reset; // @[RegFile.scala 66:20:@128700.4]
  wire [63:0] regs_265_io_in; // @[RegFile.scala 66:20:@128700.4]
  wire  regs_265_io_reset; // @[RegFile.scala 66:20:@128700.4]
  wire [63:0] regs_265_io_out; // @[RegFile.scala 66:20:@128700.4]
  wire  regs_265_io_enable; // @[RegFile.scala 66:20:@128700.4]
  wire  regs_266_clock; // @[RegFile.scala 66:20:@128714.4]
  wire  regs_266_reset; // @[RegFile.scala 66:20:@128714.4]
  wire [63:0] regs_266_io_in; // @[RegFile.scala 66:20:@128714.4]
  wire  regs_266_io_reset; // @[RegFile.scala 66:20:@128714.4]
  wire [63:0] regs_266_io_out; // @[RegFile.scala 66:20:@128714.4]
  wire  regs_266_io_enable; // @[RegFile.scala 66:20:@128714.4]
  wire  regs_267_clock; // @[RegFile.scala 66:20:@128728.4]
  wire  regs_267_reset; // @[RegFile.scala 66:20:@128728.4]
  wire [63:0] regs_267_io_in; // @[RegFile.scala 66:20:@128728.4]
  wire  regs_267_io_reset; // @[RegFile.scala 66:20:@128728.4]
  wire [63:0] regs_267_io_out; // @[RegFile.scala 66:20:@128728.4]
  wire  regs_267_io_enable; // @[RegFile.scala 66:20:@128728.4]
  wire  regs_268_clock; // @[RegFile.scala 66:20:@128742.4]
  wire  regs_268_reset; // @[RegFile.scala 66:20:@128742.4]
  wire [63:0] regs_268_io_in; // @[RegFile.scala 66:20:@128742.4]
  wire  regs_268_io_reset; // @[RegFile.scala 66:20:@128742.4]
  wire [63:0] regs_268_io_out; // @[RegFile.scala 66:20:@128742.4]
  wire  regs_268_io_enable; // @[RegFile.scala 66:20:@128742.4]
  wire  regs_269_clock; // @[RegFile.scala 66:20:@128756.4]
  wire  regs_269_reset; // @[RegFile.scala 66:20:@128756.4]
  wire [63:0] regs_269_io_in; // @[RegFile.scala 66:20:@128756.4]
  wire  regs_269_io_reset; // @[RegFile.scala 66:20:@128756.4]
  wire [63:0] regs_269_io_out; // @[RegFile.scala 66:20:@128756.4]
  wire  regs_269_io_enable; // @[RegFile.scala 66:20:@128756.4]
  wire  regs_270_clock; // @[RegFile.scala 66:20:@128770.4]
  wire  regs_270_reset; // @[RegFile.scala 66:20:@128770.4]
  wire [63:0] regs_270_io_in; // @[RegFile.scala 66:20:@128770.4]
  wire  regs_270_io_reset; // @[RegFile.scala 66:20:@128770.4]
  wire [63:0] regs_270_io_out; // @[RegFile.scala 66:20:@128770.4]
  wire  regs_270_io_enable; // @[RegFile.scala 66:20:@128770.4]
  wire  regs_271_clock; // @[RegFile.scala 66:20:@128784.4]
  wire  regs_271_reset; // @[RegFile.scala 66:20:@128784.4]
  wire [63:0] regs_271_io_in; // @[RegFile.scala 66:20:@128784.4]
  wire  regs_271_io_reset; // @[RegFile.scala 66:20:@128784.4]
  wire [63:0] regs_271_io_out; // @[RegFile.scala 66:20:@128784.4]
  wire  regs_271_io_enable; // @[RegFile.scala 66:20:@128784.4]
  wire  regs_272_clock; // @[RegFile.scala 66:20:@128798.4]
  wire  regs_272_reset; // @[RegFile.scala 66:20:@128798.4]
  wire [63:0] regs_272_io_in; // @[RegFile.scala 66:20:@128798.4]
  wire  regs_272_io_reset; // @[RegFile.scala 66:20:@128798.4]
  wire [63:0] regs_272_io_out; // @[RegFile.scala 66:20:@128798.4]
  wire  regs_272_io_enable; // @[RegFile.scala 66:20:@128798.4]
  wire  regs_273_clock; // @[RegFile.scala 66:20:@128812.4]
  wire  regs_273_reset; // @[RegFile.scala 66:20:@128812.4]
  wire [63:0] regs_273_io_in; // @[RegFile.scala 66:20:@128812.4]
  wire  regs_273_io_reset; // @[RegFile.scala 66:20:@128812.4]
  wire [63:0] regs_273_io_out; // @[RegFile.scala 66:20:@128812.4]
  wire  regs_273_io_enable; // @[RegFile.scala 66:20:@128812.4]
  wire  regs_274_clock; // @[RegFile.scala 66:20:@128826.4]
  wire  regs_274_reset; // @[RegFile.scala 66:20:@128826.4]
  wire [63:0] regs_274_io_in; // @[RegFile.scala 66:20:@128826.4]
  wire  regs_274_io_reset; // @[RegFile.scala 66:20:@128826.4]
  wire [63:0] regs_274_io_out; // @[RegFile.scala 66:20:@128826.4]
  wire  regs_274_io_enable; // @[RegFile.scala 66:20:@128826.4]
  wire  regs_275_clock; // @[RegFile.scala 66:20:@128840.4]
  wire  regs_275_reset; // @[RegFile.scala 66:20:@128840.4]
  wire [63:0] regs_275_io_in; // @[RegFile.scala 66:20:@128840.4]
  wire  regs_275_io_reset; // @[RegFile.scala 66:20:@128840.4]
  wire [63:0] regs_275_io_out; // @[RegFile.scala 66:20:@128840.4]
  wire  regs_275_io_enable; // @[RegFile.scala 66:20:@128840.4]
  wire  regs_276_clock; // @[RegFile.scala 66:20:@128854.4]
  wire  regs_276_reset; // @[RegFile.scala 66:20:@128854.4]
  wire [63:0] regs_276_io_in; // @[RegFile.scala 66:20:@128854.4]
  wire  regs_276_io_reset; // @[RegFile.scala 66:20:@128854.4]
  wire [63:0] regs_276_io_out; // @[RegFile.scala 66:20:@128854.4]
  wire  regs_276_io_enable; // @[RegFile.scala 66:20:@128854.4]
  wire  regs_277_clock; // @[RegFile.scala 66:20:@128868.4]
  wire  regs_277_reset; // @[RegFile.scala 66:20:@128868.4]
  wire [63:0] regs_277_io_in; // @[RegFile.scala 66:20:@128868.4]
  wire  regs_277_io_reset; // @[RegFile.scala 66:20:@128868.4]
  wire [63:0] regs_277_io_out; // @[RegFile.scala 66:20:@128868.4]
  wire  regs_277_io_enable; // @[RegFile.scala 66:20:@128868.4]
  wire  regs_278_clock; // @[RegFile.scala 66:20:@128882.4]
  wire  regs_278_reset; // @[RegFile.scala 66:20:@128882.4]
  wire [63:0] regs_278_io_in; // @[RegFile.scala 66:20:@128882.4]
  wire  regs_278_io_reset; // @[RegFile.scala 66:20:@128882.4]
  wire [63:0] regs_278_io_out; // @[RegFile.scala 66:20:@128882.4]
  wire  regs_278_io_enable; // @[RegFile.scala 66:20:@128882.4]
  wire  regs_279_clock; // @[RegFile.scala 66:20:@128896.4]
  wire  regs_279_reset; // @[RegFile.scala 66:20:@128896.4]
  wire [63:0] regs_279_io_in; // @[RegFile.scala 66:20:@128896.4]
  wire  regs_279_io_reset; // @[RegFile.scala 66:20:@128896.4]
  wire [63:0] regs_279_io_out; // @[RegFile.scala 66:20:@128896.4]
  wire  regs_279_io_enable; // @[RegFile.scala 66:20:@128896.4]
  wire  regs_280_clock; // @[RegFile.scala 66:20:@128910.4]
  wire  regs_280_reset; // @[RegFile.scala 66:20:@128910.4]
  wire [63:0] regs_280_io_in; // @[RegFile.scala 66:20:@128910.4]
  wire  regs_280_io_reset; // @[RegFile.scala 66:20:@128910.4]
  wire [63:0] regs_280_io_out; // @[RegFile.scala 66:20:@128910.4]
  wire  regs_280_io_enable; // @[RegFile.scala 66:20:@128910.4]
  wire  regs_281_clock; // @[RegFile.scala 66:20:@128924.4]
  wire  regs_281_reset; // @[RegFile.scala 66:20:@128924.4]
  wire [63:0] regs_281_io_in; // @[RegFile.scala 66:20:@128924.4]
  wire  regs_281_io_reset; // @[RegFile.scala 66:20:@128924.4]
  wire [63:0] regs_281_io_out; // @[RegFile.scala 66:20:@128924.4]
  wire  regs_281_io_enable; // @[RegFile.scala 66:20:@128924.4]
  wire  regs_282_clock; // @[RegFile.scala 66:20:@128938.4]
  wire  regs_282_reset; // @[RegFile.scala 66:20:@128938.4]
  wire [63:0] regs_282_io_in; // @[RegFile.scala 66:20:@128938.4]
  wire  regs_282_io_reset; // @[RegFile.scala 66:20:@128938.4]
  wire [63:0] regs_282_io_out; // @[RegFile.scala 66:20:@128938.4]
  wire  regs_282_io_enable; // @[RegFile.scala 66:20:@128938.4]
  wire  regs_283_clock; // @[RegFile.scala 66:20:@128952.4]
  wire  regs_283_reset; // @[RegFile.scala 66:20:@128952.4]
  wire [63:0] regs_283_io_in; // @[RegFile.scala 66:20:@128952.4]
  wire  regs_283_io_reset; // @[RegFile.scala 66:20:@128952.4]
  wire [63:0] regs_283_io_out; // @[RegFile.scala 66:20:@128952.4]
  wire  regs_283_io_enable; // @[RegFile.scala 66:20:@128952.4]
  wire  regs_284_clock; // @[RegFile.scala 66:20:@128966.4]
  wire  regs_284_reset; // @[RegFile.scala 66:20:@128966.4]
  wire [63:0] regs_284_io_in; // @[RegFile.scala 66:20:@128966.4]
  wire  regs_284_io_reset; // @[RegFile.scala 66:20:@128966.4]
  wire [63:0] regs_284_io_out; // @[RegFile.scala 66:20:@128966.4]
  wire  regs_284_io_enable; // @[RegFile.scala 66:20:@128966.4]
  wire  regs_285_clock; // @[RegFile.scala 66:20:@128980.4]
  wire  regs_285_reset; // @[RegFile.scala 66:20:@128980.4]
  wire [63:0] regs_285_io_in; // @[RegFile.scala 66:20:@128980.4]
  wire  regs_285_io_reset; // @[RegFile.scala 66:20:@128980.4]
  wire [63:0] regs_285_io_out; // @[RegFile.scala 66:20:@128980.4]
  wire  regs_285_io_enable; // @[RegFile.scala 66:20:@128980.4]
  wire  regs_286_clock; // @[RegFile.scala 66:20:@128994.4]
  wire  regs_286_reset; // @[RegFile.scala 66:20:@128994.4]
  wire [63:0] regs_286_io_in; // @[RegFile.scala 66:20:@128994.4]
  wire  regs_286_io_reset; // @[RegFile.scala 66:20:@128994.4]
  wire [63:0] regs_286_io_out; // @[RegFile.scala 66:20:@128994.4]
  wire  regs_286_io_enable; // @[RegFile.scala 66:20:@128994.4]
  wire  regs_287_clock; // @[RegFile.scala 66:20:@129008.4]
  wire  regs_287_reset; // @[RegFile.scala 66:20:@129008.4]
  wire [63:0] regs_287_io_in; // @[RegFile.scala 66:20:@129008.4]
  wire  regs_287_io_reset; // @[RegFile.scala 66:20:@129008.4]
  wire [63:0] regs_287_io_out; // @[RegFile.scala 66:20:@129008.4]
  wire  regs_287_io_enable; // @[RegFile.scala 66:20:@129008.4]
  wire  regs_288_clock; // @[RegFile.scala 66:20:@129022.4]
  wire  regs_288_reset; // @[RegFile.scala 66:20:@129022.4]
  wire [63:0] regs_288_io_in; // @[RegFile.scala 66:20:@129022.4]
  wire  regs_288_io_reset; // @[RegFile.scala 66:20:@129022.4]
  wire [63:0] regs_288_io_out; // @[RegFile.scala 66:20:@129022.4]
  wire  regs_288_io_enable; // @[RegFile.scala 66:20:@129022.4]
  wire  regs_289_clock; // @[RegFile.scala 66:20:@129036.4]
  wire  regs_289_reset; // @[RegFile.scala 66:20:@129036.4]
  wire [63:0] regs_289_io_in; // @[RegFile.scala 66:20:@129036.4]
  wire  regs_289_io_reset; // @[RegFile.scala 66:20:@129036.4]
  wire [63:0] regs_289_io_out; // @[RegFile.scala 66:20:@129036.4]
  wire  regs_289_io_enable; // @[RegFile.scala 66:20:@129036.4]
  wire  regs_290_clock; // @[RegFile.scala 66:20:@129050.4]
  wire  regs_290_reset; // @[RegFile.scala 66:20:@129050.4]
  wire [63:0] regs_290_io_in; // @[RegFile.scala 66:20:@129050.4]
  wire  regs_290_io_reset; // @[RegFile.scala 66:20:@129050.4]
  wire [63:0] regs_290_io_out; // @[RegFile.scala 66:20:@129050.4]
  wire  regs_290_io_enable; // @[RegFile.scala 66:20:@129050.4]
  wire  regs_291_clock; // @[RegFile.scala 66:20:@129064.4]
  wire  regs_291_reset; // @[RegFile.scala 66:20:@129064.4]
  wire [63:0] regs_291_io_in; // @[RegFile.scala 66:20:@129064.4]
  wire  regs_291_io_reset; // @[RegFile.scala 66:20:@129064.4]
  wire [63:0] regs_291_io_out; // @[RegFile.scala 66:20:@129064.4]
  wire  regs_291_io_enable; // @[RegFile.scala 66:20:@129064.4]
  wire  regs_292_clock; // @[RegFile.scala 66:20:@129078.4]
  wire  regs_292_reset; // @[RegFile.scala 66:20:@129078.4]
  wire [63:0] regs_292_io_in; // @[RegFile.scala 66:20:@129078.4]
  wire  regs_292_io_reset; // @[RegFile.scala 66:20:@129078.4]
  wire [63:0] regs_292_io_out; // @[RegFile.scala 66:20:@129078.4]
  wire  regs_292_io_enable; // @[RegFile.scala 66:20:@129078.4]
  wire  regs_293_clock; // @[RegFile.scala 66:20:@129092.4]
  wire  regs_293_reset; // @[RegFile.scala 66:20:@129092.4]
  wire [63:0] regs_293_io_in; // @[RegFile.scala 66:20:@129092.4]
  wire  regs_293_io_reset; // @[RegFile.scala 66:20:@129092.4]
  wire [63:0] regs_293_io_out; // @[RegFile.scala 66:20:@129092.4]
  wire  regs_293_io_enable; // @[RegFile.scala 66:20:@129092.4]
  wire  regs_294_clock; // @[RegFile.scala 66:20:@129106.4]
  wire  regs_294_reset; // @[RegFile.scala 66:20:@129106.4]
  wire [63:0] regs_294_io_in; // @[RegFile.scala 66:20:@129106.4]
  wire  regs_294_io_reset; // @[RegFile.scala 66:20:@129106.4]
  wire [63:0] regs_294_io_out; // @[RegFile.scala 66:20:@129106.4]
  wire  regs_294_io_enable; // @[RegFile.scala 66:20:@129106.4]
  wire  regs_295_clock; // @[RegFile.scala 66:20:@129120.4]
  wire  regs_295_reset; // @[RegFile.scala 66:20:@129120.4]
  wire [63:0] regs_295_io_in; // @[RegFile.scala 66:20:@129120.4]
  wire  regs_295_io_reset; // @[RegFile.scala 66:20:@129120.4]
  wire [63:0] regs_295_io_out; // @[RegFile.scala 66:20:@129120.4]
  wire  regs_295_io_enable; // @[RegFile.scala 66:20:@129120.4]
  wire  regs_296_clock; // @[RegFile.scala 66:20:@129134.4]
  wire  regs_296_reset; // @[RegFile.scala 66:20:@129134.4]
  wire [63:0] regs_296_io_in; // @[RegFile.scala 66:20:@129134.4]
  wire  regs_296_io_reset; // @[RegFile.scala 66:20:@129134.4]
  wire [63:0] regs_296_io_out; // @[RegFile.scala 66:20:@129134.4]
  wire  regs_296_io_enable; // @[RegFile.scala 66:20:@129134.4]
  wire  regs_297_clock; // @[RegFile.scala 66:20:@129148.4]
  wire  regs_297_reset; // @[RegFile.scala 66:20:@129148.4]
  wire [63:0] regs_297_io_in; // @[RegFile.scala 66:20:@129148.4]
  wire  regs_297_io_reset; // @[RegFile.scala 66:20:@129148.4]
  wire [63:0] regs_297_io_out; // @[RegFile.scala 66:20:@129148.4]
  wire  regs_297_io_enable; // @[RegFile.scala 66:20:@129148.4]
  wire  regs_298_clock; // @[RegFile.scala 66:20:@129162.4]
  wire  regs_298_reset; // @[RegFile.scala 66:20:@129162.4]
  wire [63:0] regs_298_io_in; // @[RegFile.scala 66:20:@129162.4]
  wire  regs_298_io_reset; // @[RegFile.scala 66:20:@129162.4]
  wire [63:0] regs_298_io_out; // @[RegFile.scala 66:20:@129162.4]
  wire  regs_298_io_enable; // @[RegFile.scala 66:20:@129162.4]
  wire  regs_299_clock; // @[RegFile.scala 66:20:@129176.4]
  wire  regs_299_reset; // @[RegFile.scala 66:20:@129176.4]
  wire [63:0] regs_299_io_in; // @[RegFile.scala 66:20:@129176.4]
  wire  regs_299_io_reset; // @[RegFile.scala 66:20:@129176.4]
  wire [63:0] regs_299_io_out; // @[RegFile.scala 66:20:@129176.4]
  wire  regs_299_io_enable; // @[RegFile.scala 66:20:@129176.4]
  wire  regs_300_clock; // @[RegFile.scala 66:20:@129190.4]
  wire  regs_300_reset; // @[RegFile.scala 66:20:@129190.4]
  wire [63:0] regs_300_io_in; // @[RegFile.scala 66:20:@129190.4]
  wire  regs_300_io_reset; // @[RegFile.scala 66:20:@129190.4]
  wire [63:0] regs_300_io_out; // @[RegFile.scala 66:20:@129190.4]
  wire  regs_300_io_enable; // @[RegFile.scala 66:20:@129190.4]
  wire  regs_301_clock; // @[RegFile.scala 66:20:@129204.4]
  wire  regs_301_reset; // @[RegFile.scala 66:20:@129204.4]
  wire [63:0] regs_301_io_in; // @[RegFile.scala 66:20:@129204.4]
  wire  regs_301_io_reset; // @[RegFile.scala 66:20:@129204.4]
  wire [63:0] regs_301_io_out; // @[RegFile.scala 66:20:@129204.4]
  wire  regs_301_io_enable; // @[RegFile.scala 66:20:@129204.4]
  wire  regs_302_clock; // @[RegFile.scala 66:20:@129218.4]
  wire  regs_302_reset; // @[RegFile.scala 66:20:@129218.4]
  wire [63:0] regs_302_io_in; // @[RegFile.scala 66:20:@129218.4]
  wire  regs_302_io_reset; // @[RegFile.scala 66:20:@129218.4]
  wire [63:0] regs_302_io_out; // @[RegFile.scala 66:20:@129218.4]
  wire  regs_302_io_enable; // @[RegFile.scala 66:20:@129218.4]
  wire  regs_303_clock; // @[RegFile.scala 66:20:@129232.4]
  wire  regs_303_reset; // @[RegFile.scala 66:20:@129232.4]
  wire [63:0] regs_303_io_in; // @[RegFile.scala 66:20:@129232.4]
  wire  regs_303_io_reset; // @[RegFile.scala 66:20:@129232.4]
  wire [63:0] regs_303_io_out; // @[RegFile.scala 66:20:@129232.4]
  wire  regs_303_io_enable; // @[RegFile.scala 66:20:@129232.4]
  wire  regs_304_clock; // @[RegFile.scala 66:20:@129246.4]
  wire  regs_304_reset; // @[RegFile.scala 66:20:@129246.4]
  wire [63:0] regs_304_io_in; // @[RegFile.scala 66:20:@129246.4]
  wire  regs_304_io_reset; // @[RegFile.scala 66:20:@129246.4]
  wire [63:0] regs_304_io_out; // @[RegFile.scala 66:20:@129246.4]
  wire  regs_304_io_enable; // @[RegFile.scala 66:20:@129246.4]
  wire  regs_305_clock; // @[RegFile.scala 66:20:@129260.4]
  wire  regs_305_reset; // @[RegFile.scala 66:20:@129260.4]
  wire [63:0] regs_305_io_in; // @[RegFile.scala 66:20:@129260.4]
  wire  regs_305_io_reset; // @[RegFile.scala 66:20:@129260.4]
  wire [63:0] regs_305_io_out; // @[RegFile.scala 66:20:@129260.4]
  wire  regs_305_io_enable; // @[RegFile.scala 66:20:@129260.4]
  wire  regs_306_clock; // @[RegFile.scala 66:20:@129274.4]
  wire  regs_306_reset; // @[RegFile.scala 66:20:@129274.4]
  wire [63:0] regs_306_io_in; // @[RegFile.scala 66:20:@129274.4]
  wire  regs_306_io_reset; // @[RegFile.scala 66:20:@129274.4]
  wire [63:0] regs_306_io_out; // @[RegFile.scala 66:20:@129274.4]
  wire  regs_306_io_enable; // @[RegFile.scala 66:20:@129274.4]
  wire  regs_307_clock; // @[RegFile.scala 66:20:@129288.4]
  wire  regs_307_reset; // @[RegFile.scala 66:20:@129288.4]
  wire [63:0] regs_307_io_in; // @[RegFile.scala 66:20:@129288.4]
  wire  regs_307_io_reset; // @[RegFile.scala 66:20:@129288.4]
  wire [63:0] regs_307_io_out; // @[RegFile.scala 66:20:@129288.4]
  wire  regs_307_io_enable; // @[RegFile.scala 66:20:@129288.4]
  wire  regs_308_clock; // @[RegFile.scala 66:20:@129302.4]
  wire  regs_308_reset; // @[RegFile.scala 66:20:@129302.4]
  wire [63:0] regs_308_io_in; // @[RegFile.scala 66:20:@129302.4]
  wire  regs_308_io_reset; // @[RegFile.scala 66:20:@129302.4]
  wire [63:0] regs_308_io_out; // @[RegFile.scala 66:20:@129302.4]
  wire  regs_308_io_enable; // @[RegFile.scala 66:20:@129302.4]
  wire  regs_309_clock; // @[RegFile.scala 66:20:@129316.4]
  wire  regs_309_reset; // @[RegFile.scala 66:20:@129316.4]
  wire [63:0] regs_309_io_in; // @[RegFile.scala 66:20:@129316.4]
  wire  regs_309_io_reset; // @[RegFile.scala 66:20:@129316.4]
  wire [63:0] regs_309_io_out; // @[RegFile.scala 66:20:@129316.4]
  wire  regs_309_io_enable; // @[RegFile.scala 66:20:@129316.4]
  wire  regs_310_clock; // @[RegFile.scala 66:20:@129330.4]
  wire  regs_310_reset; // @[RegFile.scala 66:20:@129330.4]
  wire [63:0] regs_310_io_in; // @[RegFile.scala 66:20:@129330.4]
  wire  regs_310_io_reset; // @[RegFile.scala 66:20:@129330.4]
  wire [63:0] regs_310_io_out; // @[RegFile.scala 66:20:@129330.4]
  wire  regs_310_io_enable; // @[RegFile.scala 66:20:@129330.4]
  wire  regs_311_clock; // @[RegFile.scala 66:20:@129344.4]
  wire  regs_311_reset; // @[RegFile.scala 66:20:@129344.4]
  wire [63:0] regs_311_io_in; // @[RegFile.scala 66:20:@129344.4]
  wire  regs_311_io_reset; // @[RegFile.scala 66:20:@129344.4]
  wire [63:0] regs_311_io_out; // @[RegFile.scala 66:20:@129344.4]
  wire  regs_311_io_enable; // @[RegFile.scala 66:20:@129344.4]
  wire  regs_312_clock; // @[RegFile.scala 66:20:@129358.4]
  wire  regs_312_reset; // @[RegFile.scala 66:20:@129358.4]
  wire [63:0] regs_312_io_in; // @[RegFile.scala 66:20:@129358.4]
  wire  regs_312_io_reset; // @[RegFile.scala 66:20:@129358.4]
  wire [63:0] regs_312_io_out; // @[RegFile.scala 66:20:@129358.4]
  wire  regs_312_io_enable; // @[RegFile.scala 66:20:@129358.4]
  wire  regs_313_clock; // @[RegFile.scala 66:20:@129372.4]
  wire  regs_313_reset; // @[RegFile.scala 66:20:@129372.4]
  wire [63:0] regs_313_io_in; // @[RegFile.scala 66:20:@129372.4]
  wire  regs_313_io_reset; // @[RegFile.scala 66:20:@129372.4]
  wire [63:0] regs_313_io_out; // @[RegFile.scala 66:20:@129372.4]
  wire  regs_313_io_enable; // @[RegFile.scala 66:20:@129372.4]
  wire  regs_314_clock; // @[RegFile.scala 66:20:@129386.4]
  wire  regs_314_reset; // @[RegFile.scala 66:20:@129386.4]
  wire [63:0] regs_314_io_in; // @[RegFile.scala 66:20:@129386.4]
  wire  regs_314_io_reset; // @[RegFile.scala 66:20:@129386.4]
  wire [63:0] regs_314_io_out; // @[RegFile.scala 66:20:@129386.4]
  wire  regs_314_io_enable; // @[RegFile.scala 66:20:@129386.4]
  wire  regs_315_clock; // @[RegFile.scala 66:20:@129400.4]
  wire  regs_315_reset; // @[RegFile.scala 66:20:@129400.4]
  wire [63:0] regs_315_io_in; // @[RegFile.scala 66:20:@129400.4]
  wire  regs_315_io_reset; // @[RegFile.scala 66:20:@129400.4]
  wire [63:0] regs_315_io_out; // @[RegFile.scala 66:20:@129400.4]
  wire  regs_315_io_enable; // @[RegFile.scala 66:20:@129400.4]
  wire  regs_316_clock; // @[RegFile.scala 66:20:@129414.4]
  wire  regs_316_reset; // @[RegFile.scala 66:20:@129414.4]
  wire [63:0] regs_316_io_in; // @[RegFile.scala 66:20:@129414.4]
  wire  regs_316_io_reset; // @[RegFile.scala 66:20:@129414.4]
  wire [63:0] regs_316_io_out; // @[RegFile.scala 66:20:@129414.4]
  wire  regs_316_io_enable; // @[RegFile.scala 66:20:@129414.4]
  wire  regs_317_clock; // @[RegFile.scala 66:20:@129428.4]
  wire  regs_317_reset; // @[RegFile.scala 66:20:@129428.4]
  wire [63:0] regs_317_io_in; // @[RegFile.scala 66:20:@129428.4]
  wire  regs_317_io_reset; // @[RegFile.scala 66:20:@129428.4]
  wire [63:0] regs_317_io_out; // @[RegFile.scala 66:20:@129428.4]
  wire  regs_317_io_enable; // @[RegFile.scala 66:20:@129428.4]
  wire  regs_318_clock; // @[RegFile.scala 66:20:@129442.4]
  wire  regs_318_reset; // @[RegFile.scala 66:20:@129442.4]
  wire [63:0] regs_318_io_in; // @[RegFile.scala 66:20:@129442.4]
  wire  regs_318_io_reset; // @[RegFile.scala 66:20:@129442.4]
  wire [63:0] regs_318_io_out; // @[RegFile.scala 66:20:@129442.4]
  wire  regs_318_io_enable; // @[RegFile.scala 66:20:@129442.4]
  wire  regs_319_clock; // @[RegFile.scala 66:20:@129456.4]
  wire  regs_319_reset; // @[RegFile.scala 66:20:@129456.4]
  wire [63:0] regs_319_io_in; // @[RegFile.scala 66:20:@129456.4]
  wire  regs_319_io_reset; // @[RegFile.scala 66:20:@129456.4]
  wire [63:0] regs_319_io_out; // @[RegFile.scala 66:20:@129456.4]
  wire  regs_319_io_enable; // @[RegFile.scala 66:20:@129456.4]
  wire  regs_320_clock; // @[RegFile.scala 66:20:@129470.4]
  wire  regs_320_reset; // @[RegFile.scala 66:20:@129470.4]
  wire [63:0] regs_320_io_in; // @[RegFile.scala 66:20:@129470.4]
  wire  regs_320_io_reset; // @[RegFile.scala 66:20:@129470.4]
  wire [63:0] regs_320_io_out; // @[RegFile.scala 66:20:@129470.4]
  wire  regs_320_io_enable; // @[RegFile.scala 66:20:@129470.4]
  wire  regs_321_clock; // @[RegFile.scala 66:20:@129484.4]
  wire  regs_321_reset; // @[RegFile.scala 66:20:@129484.4]
  wire [63:0] regs_321_io_in; // @[RegFile.scala 66:20:@129484.4]
  wire  regs_321_io_reset; // @[RegFile.scala 66:20:@129484.4]
  wire [63:0] regs_321_io_out; // @[RegFile.scala 66:20:@129484.4]
  wire  regs_321_io_enable; // @[RegFile.scala 66:20:@129484.4]
  wire  regs_322_clock; // @[RegFile.scala 66:20:@129498.4]
  wire  regs_322_reset; // @[RegFile.scala 66:20:@129498.4]
  wire [63:0] regs_322_io_in; // @[RegFile.scala 66:20:@129498.4]
  wire  regs_322_io_reset; // @[RegFile.scala 66:20:@129498.4]
  wire [63:0] regs_322_io_out; // @[RegFile.scala 66:20:@129498.4]
  wire  regs_322_io_enable; // @[RegFile.scala 66:20:@129498.4]
  wire  regs_323_clock; // @[RegFile.scala 66:20:@129512.4]
  wire  regs_323_reset; // @[RegFile.scala 66:20:@129512.4]
  wire [63:0] regs_323_io_in; // @[RegFile.scala 66:20:@129512.4]
  wire  regs_323_io_reset; // @[RegFile.scala 66:20:@129512.4]
  wire [63:0] regs_323_io_out; // @[RegFile.scala 66:20:@129512.4]
  wire  regs_323_io_enable; // @[RegFile.scala 66:20:@129512.4]
  wire  regs_324_clock; // @[RegFile.scala 66:20:@129526.4]
  wire  regs_324_reset; // @[RegFile.scala 66:20:@129526.4]
  wire [63:0] regs_324_io_in; // @[RegFile.scala 66:20:@129526.4]
  wire  regs_324_io_reset; // @[RegFile.scala 66:20:@129526.4]
  wire [63:0] regs_324_io_out; // @[RegFile.scala 66:20:@129526.4]
  wire  regs_324_io_enable; // @[RegFile.scala 66:20:@129526.4]
  wire  regs_325_clock; // @[RegFile.scala 66:20:@129540.4]
  wire  regs_325_reset; // @[RegFile.scala 66:20:@129540.4]
  wire [63:0] regs_325_io_in; // @[RegFile.scala 66:20:@129540.4]
  wire  regs_325_io_reset; // @[RegFile.scala 66:20:@129540.4]
  wire [63:0] regs_325_io_out; // @[RegFile.scala 66:20:@129540.4]
  wire  regs_325_io_enable; // @[RegFile.scala 66:20:@129540.4]
  wire  regs_326_clock; // @[RegFile.scala 66:20:@129554.4]
  wire  regs_326_reset; // @[RegFile.scala 66:20:@129554.4]
  wire [63:0] regs_326_io_in; // @[RegFile.scala 66:20:@129554.4]
  wire  regs_326_io_reset; // @[RegFile.scala 66:20:@129554.4]
  wire [63:0] regs_326_io_out; // @[RegFile.scala 66:20:@129554.4]
  wire  regs_326_io_enable; // @[RegFile.scala 66:20:@129554.4]
  wire  regs_327_clock; // @[RegFile.scala 66:20:@129568.4]
  wire  regs_327_reset; // @[RegFile.scala 66:20:@129568.4]
  wire [63:0] regs_327_io_in; // @[RegFile.scala 66:20:@129568.4]
  wire  regs_327_io_reset; // @[RegFile.scala 66:20:@129568.4]
  wire [63:0] regs_327_io_out; // @[RegFile.scala 66:20:@129568.4]
  wire  regs_327_io_enable; // @[RegFile.scala 66:20:@129568.4]
  wire  regs_328_clock; // @[RegFile.scala 66:20:@129582.4]
  wire  regs_328_reset; // @[RegFile.scala 66:20:@129582.4]
  wire [63:0] regs_328_io_in; // @[RegFile.scala 66:20:@129582.4]
  wire  regs_328_io_reset; // @[RegFile.scala 66:20:@129582.4]
  wire [63:0] regs_328_io_out; // @[RegFile.scala 66:20:@129582.4]
  wire  regs_328_io_enable; // @[RegFile.scala 66:20:@129582.4]
  wire  regs_329_clock; // @[RegFile.scala 66:20:@129596.4]
  wire  regs_329_reset; // @[RegFile.scala 66:20:@129596.4]
  wire [63:0] regs_329_io_in; // @[RegFile.scala 66:20:@129596.4]
  wire  regs_329_io_reset; // @[RegFile.scala 66:20:@129596.4]
  wire [63:0] regs_329_io_out; // @[RegFile.scala 66:20:@129596.4]
  wire  regs_329_io_enable; // @[RegFile.scala 66:20:@129596.4]
  wire  regs_330_clock; // @[RegFile.scala 66:20:@129610.4]
  wire  regs_330_reset; // @[RegFile.scala 66:20:@129610.4]
  wire [63:0] regs_330_io_in; // @[RegFile.scala 66:20:@129610.4]
  wire  regs_330_io_reset; // @[RegFile.scala 66:20:@129610.4]
  wire [63:0] regs_330_io_out; // @[RegFile.scala 66:20:@129610.4]
  wire  regs_330_io_enable; // @[RegFile.scala 66:20:@129610.4]
  wire  regs_331_clock; // @[RegFile.scala 66:20:@129624.4]
  wire  regs_331_reset; // @[RegFile.scala 66:20:@129624.4]
  wire [63:0] regs_331_io_in; // @[RegFile.scala 66:20:@129624.4]
  wire  regs_331_io_reset; // @[RegFile.scala 66:20:@129624.4]
  wire [63:0] regs_331_io_out; // @[RegFile.scala 66:20:@129624.4]
  wire  regs_331_io_enable; // @[RegFile.scala 66:20:@129624.4]
  wire  regs_332_clock; // @[RegFile.scala 66:20:@129638.4]
  wire  regs_332_reset; // @[RegFile.scala 66:20:@129638.4]
  wire [63:0] regs_332_io_in; // @[RegFile.scala 66:20:@129638.4]
  wire  regs_332_io_reset; // @[RegFile.scala 66:20:@129638.4]
  wire [63:0] regs_332_io_out; // @[RegFile.scala 66:20:@129638.4]
  wire  regs_332_io_enable; // @[RegFile.scala 66:20:@129638.4]
  wire  regs_333_clock; // @[RegFile.scala 66:20:@129652.4]
  wire  regs_333_reset; // @[RegFile.scala 66:20:@129652.4]
  wire [63:0] regs_333_io_in; // @[RegFile.scala 66:20:@129652.4]
  wire  regs_333_io_reset; // @[RegFile.scala 66:20:@129652.4]
  wire [63:0] regs_333_io_out; // @[RegFile.scala 66:20:@129652.4]
  wire  regs_333_io_enable; // @[RegFile.scala 66:20:@129652.4]
  wire  regs_334_clock; // @[RegFile.scala 66:20:@129666.4]
  wire  regs_334_reset; // @[RegFile.scala 66:20:@129666.4]
  wire [63:0] regs_334_io_in; // @[RegFile.scala 66:20:@129666.4]
  wire  regs_334_io_reset; // @[RegFile.scala 66:20:@129666.4]
  wire [63:0] regs_334_io_out; // @[RegFile.scala 66:20:@129666.4]
  wire  regs_334_io_enable; // @[RegFile.scala 66:20:@129666.4]
  wire  regs_335_clock; // @[RegFile.scala 66:20:@129680.4]
  wire  regs_335_reset; // @[RegFile.scala 66:20:@129680.4]
  wire [63:0] regs_335_io_in; // @[RegFile.scala 66:20:@129680.4]
  wire  regs_335_io_reset; // @[RegFile.scala 66:20:@129680.4]
  wire [63:0] regs_335_io_out; // @[RegFile.scala 66:20:@129680.4]
  wire  regs_335_io_enable; // @[RegFile.scala 66:20:@129680.4]
  wire  regs_336_clock; // @[RegFile.scala 66:20:@129694.4]
  wire  regs_336_reset; // @[RegFile.scala 66:20:@129694.4]
  wire [63:0] regs_336_io_in; // @[RegFile.scala 66:20:@129694.4]
  wire  regs_336_io_reset; // @[RegFile.scala 66:20:@129694.4]
  wire [63:0] regs_336_io_out; // @[RegFile.scala 66:20:@129694.4]
  wire  regs_336_io_enable; // @[RegFile.scala 66:20:@129694.4]
  wire  regs_337_clock; // @[RegFile.scala 66:20:@129708.4]
  wire  regs_337_reset; // @[RegFile.scala 66:20:@129708.4]
  wire [63:0] regs_337_io_in; // @[RegFile.scala 66:20:@129708.4]
  wire  regs_337_io_reset; // @[RegFile.scala 66:20:@129708.4]
  wire [63:0] regs_337_io_out; // @[RegFile.scala 66:20:@129708.4]
  wire  regs_337_io_enable; // @[RegFile.scala 66:20:@129708.4]
  wire  regs_338_clock; // @[RegFile.scala 66:20:@129722.4]
  wire  regs_338_reset; // @[RegFile.scala 66:20:@129722.4]
  wire [63:0] regs_338_io_in; // @[RegFile.scala 66:20:@129722.4]
  wire  regs_338_io_reset; // @[RegFile.scala 66:20:@129722.4]
  wire [63:0] regs_338_io_out; // @[RegFile.scala 66:20:@129722.4]
  wire  regs_338_io_enable; // @[RegFile.scala 66:20:@129722.4]
  wire  regs_339_clock; // @[RegFile.scala 66:20:@129736.4]
  wire  regs_339_reset; // @[RegFile.scala 66:20:@129736.4]
  wire [63:0] regs_339_io_in; // @[RegFile.scala 66:20:@129736.4]
  wire  regs_339_io_reset; // @[RegFile.scala 66:20:@129736.4]
  wire [63:0] regs_339_io_out; // @[RegFile.scala 66:20:@129736.4]
  wire  regs_339_io_enable; // @[RegFile.scala 66:20:@129736.4]
  wire  regs_340_clock; // @[RegFile.scala 66:20:@129750.4]
  wire  regs_340_reset; // @[RegFile.scala 66:20:@129750.4]
  wire [63:0] regs_340_io_in; // @[RegFile.scala 66:20:@129750.4]
  wire  regs_340_io_reset; // @[RegFile.scala 66:20:@129750.4]
  wire [63:0] regs_340_io_out; // @[RegFile.scala 66:20:@129750.4]
  wire  regs_340_io_enable; // @[RegFile.scala 66:20:@129750.4]
  wire  regs_341_clock; // @[RegFile.scala 66:20:@129764.4]
  wire  regs_341_reset; // @[RegFile.scala 66:20:@129764.4]
  wire [63:0] regs_341_io_in; // @[RegFile.scala 66:20:@129764.4]
  wire  regs_341_io_reset; // @[RegFile.scala 66:20:@129764.4]
  wire [63:0] regs_341_io_out; // @[RegFile.scala 66:20:@129764.4]
  wire  regs_341_io_enable; // @[RegFile.scala 66:20:@129764.4]
  wire  regs_342_clock; // @[RegFile.scala 66:20:@129778.4]
  wire  regs_342_reset; // @[RegFile.scala 66:20:@129778.4]
  wire [63:0] regs_342_io_in; // @[RegFile.scala 66:20:@129778.4]
  wire  regs_342_io_reset; // @[RegFile.scala 66:20:@129778.4]
  wire [63:0] regs_342_io_out; // @[RegFile.scala 66:20:@129778.4]
  wire  regs_342_io_enable; // @[RegFile.scala 66:20:@129778.4]
  wire  regs_343_clock; // @[RegFile.scala 66:20:@129792.4]
  wire  regs_343_reset; // @[RegFile.scala 66:20:@129792.4]
  wire [63:0] regs_343_io_in; // @[RegFile.scala 66:20:@129792.4]
  wire  regs_343_io_reset; // @[RegFile.scala 66:20:@129792.4]
  wire [63:0] regs_343_io_out; // @[RegFile.scala 66:20:@129792.4]
  wire  regs_343_io_enable; // @[RegFile.scala 66:20:@129792.4]
  wire  regs_344_clock; // @[RegFile.scala 66:20:@129806.4]
  wire  regs_344_reset; // @[RegFile.scala 66:20:@129806.4]
  wire [63:0] regs_344_io_in; // @[RegFile.scala 66:20:@129806.4]
  wire  regs_344_io_reset; // @[RegFile.scala 66:20:@129806.4]
  wire [63:0] regs_344_io_out; // @[RegFile.scala 66:20:@129806.4]
  wire  regs_344_io_enable; // @[RegFile.scala 66:20:@129806.4]
  wire  regs_345_clock; // @[RegFile.scala 66:20:@129820.4]
  wire  regs_345_reset; // @[RegFile.scala 66:20:@129820.4]
  wire [63:0] regs_345_io_in; // @[RegFile.scala 66:20:@129820.4]
  wire  regs_345_io_reset; // @[RegFile.scala 66:20:@129820.4]
  wire [63:0] regs_345_io_out; // @[RegFile.scala 66:20:@129820.4]
  wire  regs_345_io_enable; // @[RegFile.scala 66:20:@129820.4]
  wire  regs_346_clock; // @[RegFile.scala 66:20:@129834.4]
  wire  regs_346_reset; // @[RegFile.scala 66:20:@129834.4]
  wire [63:0] regs_346_io_in; // @[RegFile.scala 66:20:@129834.4]
  wire  regs_346_io_reset; // @[RegFile.scala 66:20:@129834.4]
  wire [63:0] regs_346_io_out; // @[RegFile.scala 66:20:@129834.4]
  wire  regs_346_io_enable; // @[RegFile.scala 66:20:@129834.4]
  wire  regs_347_clock; // @[RegFile.scala 66:20:@129848.4]
  wire  regs_347_reset; // @[RegFile.scala 66:20:@129848.4]
  wire [63:0] regs_347_io_in; // @[RegFile.scala 66:20:@129848.4]
  wire  regs_347_io_reset; // @[RegFile.scala 66:20:@129848.4]
  wire [63:0] regs_347_io_out; // @[RegFile.scala 66:20:@129848.4]
  wire  regs_347_io_enable; // @[RegFile.scala 66:20:@129848.4]
  wire  regs_348_clock; // @[RegFile.scala 66:20:@129862.4]
  wire  regs_348_reset; // @[RegFile.scala 66:20:@129862.4]
  wire [63:0] regs_348_io_in; // @[RegFile.scala 66:20:@129862.4]
  wire  regs_348_io_reset; // @[RegFile.scala 66:20:@129862.4]
  wire [63:0] regs_348_io_out; // @[RegFile.scala 66:20:@129862.4]
  wire  regs_348_io_enable; // @[RegFile.scala 66:20:@129862.4]
  wire  regs_349_clock; // @[RegFile.scala 66:20:@129876.4]
  wire  regs_349_reset; // @[RegFile.scala 66:20:@129876.4]
  wire [63:0] regs_349_io_in; // @[RegFile.scala 66:20:@129876.4]
  wire  regs_349_io_reset; // @[RegFile.scala 66:20:@129876.4]
  wire [63:0] regs_349_io_out; // @[RegFile.scala 66:20:@129876.4]
  wire  regs_349_io_enable; // @[RegFile.scala 66:20:@129876.4]
  wire  regs_350_clock; // @[RegFile.scala 66:20:@129890.4]
  wire  regs_350_reset; // @[RegFile.scala 66:20:@129890.4]
  wire [63:0] regs_350_io_in; // @[RegFile.scala 66:20:@129890.4]
  wire  regs_350_io_reset; // @[RegFile.scala 66:20:@129890.4]
  wire [63:0] regs_350_io_out; // @[RegFile.scala 66:20:@129890.4]
  wire  regs_350_io_enable; // @[RegFile.scala 66:20:@129890.4]
  wire  regs_351_clock; // @[RegFile.scala 66:20:@129904.4]
  wire  regs_351_reset; // @[RegFile.scala 66:20:@129904.4]
  wire [63:0] regs_351_io_in; // @[RegFile.scala 66:20:@129904.4]
  wire  regs_351_io_reset; // @[RegFile.scala 66:20:@129904.4]
  wire [63:0] regs_351_io_out; // @[RegFile.scala 66:20:@129904.4]
  wire  regs_351_io_enable; // @[RegFile.scala 66:20:@129904.4]
  wire  regs_352_clock; // @[RegFile.scala 66:20:@129918.4]
  wire  regs_352_reset; // @[RegFile.scala 66:20:@129918.4]
  wire [63:0] regs_352_io_in; // @[RegFile.scala 66:20:@129918.4]
  wire  regs_352_io_reset; // @[RegFile.scala 66:20:@129918.4]
  wire [63:0] regs_352_io_out; // @[RegFile.scala 66:20:@129918.4]
  wire  regs_352_io_enable; // @[RegFile.scala 66:20:@129918.4]
  wire  regs_353_clock; // @[RegFile.scala 66:20:@129932.4]
  wire  regs_353_reset; // @[RegFile.scala 66:20:@129932.4]
  wire [63:0] regs_353_io_in; // @[RegFile.scala 66:20:@129932.4]
  wire  regs_353_io_reset; // @[RegFile.scala 66:20:@129932.4]
  wire [63:0] regs_353_io_out; // @[RegFile.scala 66:20:@129932.4]
  wire  regs_353_io_enable; // @[RegFile.scala 66:20:@129932.4]
  wire  regs_354_clock; // @[RegFile.scala 66:20:@129946.4]
  wire  regs_354_reset; // @[RegFile.scala 66:20:@129946.4]
  wire [63:0] regs_354_io_in; // @[RegFile.scala 66:20:@129946.4]
  wire  regs_354_io_reset; // @[RegFile.scala 66:20:@129946.4]
  wire [63:0] regs_354_io_out; // @[RegFile.scala 66:20:@129946.4]
  wire  regs_354_io_enable; // @[RegFile.scala 66:20:@129946.4]
  wire  regs_355_clock; // @[RegFile.scala 66:20:@129960.4]
  wire  regs_355_reset; // @[RegFile.scala 66:20:@129960.4]
  wire [63:0] regs_355_io_in; // @[RegFile.scala 66:20:@129960.4]
  wire  regs_355_io_reset; // @[RegFile.scala 66:20:@129960.4]
  wire [63:0] regs_355_io_out; // @[RegFile.scala 66:20:@129960.4]
  wire  regs_355_io_enable; // @[RegFile.scala 66:20:@129960.4]
  wire  regs_356_clock; // @[RegFile.scala 66:20:@129974.4]
  wire  regs_356_reset; // @[RegFile.scala 66:20:@129974.4]
  wire [63:0] regs_356_io_in; // @[RegFile.scala 66:20:@129974.4]
  wire  regs_356_io_reset; // @[RegFile.scala 66:20:@129974.4]
  wire [63:0] regs_356_io_out; // @[RegFile.scala 66:20:@129974.4]
  wire  regs_356_io_enable; // @[RegFile.scala 66:20:@129974.4]
  wire  regs_357_clock; // @[RegFile.scala 66:20:@129988.4]
  wire  regs_357_reset; // @[RegFile.scala 66:20:@129988.4]
  wire [63:0] regs_357_io_in; // @[RegFile.scala 66:20:@129988.4]
  wire  regs_357_io_reset; // @[RegFile.scala 66:20:@129988.4]
  wire [63:0] regs_357_io_out; // @[RegFile.scala 66:20:@129988.4]
  wire  regs_357_io_enable; // @[RegFile.scala 66:20:@129988.4]
  wire  regs_358_clock; // @[RegFile.scala 66:20:@130002.4]
  wire  regs_358_reset; // @[RegFile.scala 66:20:@130002.4]
  wire [63:0] regs_358_io_in; // @[RegFile.scala 66:20:@130002.4]
  wire  regs_358_io_reset; // @[RegFile.scala 66:20:@130002.4]
  wire [63:0] regs_358_io_out; // @[RegFile.scala 66:20:@130002.4]
  wire  regs_358_io_enable; // @[RegFile.scala 66:20:@130002.4]
  wire  regs_359_clock; // @[RegFile.scala 66:20:@130016.4]
  wire  regs_359_reset; // @[RegFile.scala 66:20:@130016.4]
  wire [63:0] regs_359_io_in; // @[RegFile.scala 66:20:@130016.4]
  wire  regs_359_io_reset; // @[RegFile.scala 66:20:@130016.4]
  wire [63:0] regs_359_io_out; // @[RegFile.scala 66:20:@130016.4]
  wire  regs_359_io_enable; // @[RegFile.scala 66:20:@130016.4]
  wire  regs_360_clock; // @[RegFile.scala 66:20:@130030.4]
  wire  regs_360_reset; // @[RegFile.scala 66:20:@130030.4]
  wire [63:0] regs_360_io_in; // @[RegFile.scala 66:20:@130030.4]
  wire  regs_360_io_reset; // @[RegFile.scala 66:20:@130030.4]
  wire [63:0] regs_360_io_out; // @[RegFile.scala 66:20:@130030.4]
  wire  regs_360_io_enable; // @[RegFile.scala 66:20:@130030.4]
  wire  regs_361_clock; // @[RegFile.scala 66:20:@130044.4]
  wire  regs_361_reset; // @[RegFile.scala 66:20:@130044.4]
  wire [63:0] regs_361_io_in; // @[RegFile.scala 66:20:@130044.4]
  wire  regs_361_io_reset; // @[RegFile.scala 66:20:@130044.4]
  wire [63:0] regs_361_io_out; // @[RegFile.scala 66:20:@130044.4]
  wire  regs_361_io_enable; // @[RegFile.scala 66:20:@130044.4]
  wire  regs_362_clock; // @[RegFile.scala 66:20:@130058.4]
  wire  regs_362_reset; // @[RegFile.scala 66:20:@130058.4]
  wire [63:0] regs_362_io_in; // @[RegFile.scala 66:20:@130058.4]
  wire  regs_362_io_reset; // @[RegFile.scala 66:20:@130058.4]
  wire [63:0] regs_362_io_out; // @[RegFile.scala 66:20:@130058.4]
  wire  regs_362_io_enable; // @[RegFile.scala 66:20:@130058.4]
  wire  regs_363_clock; // @[RegFile.scala 66:20:@130072.4]
  wire  regs_363_reset; // @[RegFile.scala 66:20:@130072.4]
  wire [63:0] regs_363_io_in; // @[RegFile.scala 66:20:@130072.4]
  wire  regs_363_io_reset; // @[RegFile.scala 66:20:@130072.4]
  wire [63:0] regs_363_io_out; // @[RegFile.scala 66:20:@130072.4]
  wire  regs_363_io_enable; // @[RegFile.scala 66:20:@130072.4]
  wire  regs_364_clock; // @[RegFile.scala 66:20:@130086.4]
  wire  regs_364_reset; // @[RegFile.scala 66:20:@130086.4]
  wire [63:0] regs_364_io_in; // @[RegFile.scala 66:20:@130086.4]
  wire  regs_364_io_reset; // @[RegFile.scala 66:20:@130086.4]
  wire [63:0] regs_364_io_out; // @[RegFile.scala 66:20:@130086.4]
  wire  regs_364_io_enable; // @[RegFile.scala 66:20:@130086.4]
  wire  regs_365_clock; // @[RegFile.scala 66:20:@130100.4]
  wire  regs_365_reset; // @[RegFile.scala 66:20:@130100.4]
  wire [63:0] regs_365_io_in; // @[RegFile.scala 66:20:@130100.4]
  wire  regs_365_io_reset; // @[RegFile.scala 66:20:@130100.4]
  wire [63:0] regs_365_io_out; // @[RegFile.scala 66:20:@130100.4]
  wire  regs_365_io_enable; // @[RegFile.scala 66:20:@130100.4]
  wire  regs_366_clock; // @[RegFile.scala 66:20:@130114.4]
  wire  regs_366_reset; // @[RegFile.scala 66:20:@130114.4]
  wire [63:0] regs_366_io_in; // @[RegFile.scala 66:20:@130114.4]
  wire  regs_366_io_reset; // @[RegFile.scala 66:20:@130114.4]
  wire [63:0] regs_366_io_out; // @[RegFile.scala 66:20:@130114.4]
  wire  regs_366_io_enable; // @[RegFile.scala 66:20:@130114.4]
  wire  regs_367_clock; // @[RegFile.scala 66:20:@130128.4]
  wire  regs_367_reset; // @[RegFile.scala 66:20:@130128.4]
  wire [63:0] regs_367_io_in; // @[RegFile.scala 66:20:@130128.4]
  wire  regs_367_io_reset; // @[RegFile.scala 66:20:@130128.4]
  wire [63:0] regs_367_io_out; // @[RegFile.scala 66:20:@130128.4]
  wire  regs_367_io_enable; // @[RegFile.scala 66:20:@130128.4]
  wire  regs_368_clock; // @[RegFile.scala 66:20:@130142.4]
  wire  regs_368_reset; // @[RegFile.scala 66:20:@130142.4]
  wire [63:0] regs_368_io_in; // @[RegFile.scala 66:20:@130142.4]
  wire  regs_368_io_reset; // @[RegFile.scala 66:20:@130142.4]
  wire [63:0] regs_368_io_out; // @[RegFile.scala 66:20:@130142.4]
  wire  regs_368_io_enable; // @[RegFile.scala 66:20:@130142.4]
  wire  regs_369_clock; // @[RegFile.scala 66:20:@130156.4]
  wire  regs_369_reset; // @[RegFile.scala 66:20:@130156.4]
  wire [63:0] regs_369_io_in; // @[RegFile.scala 66:20:@130156.4]
  wire  regs_369_io_reset; // @[RegFile.scala 66:20:@130156.4]
  wire [63:0] regs_369_io_out; // @[RegFile.scala 66:20:@130156.4]
  wire  regs_369_io_enable; // @[RegFile.scala 66:20:@130156.4]
  wire  regs_370_clock; // @[RegFile.scala 66:20:@130170.4]
  wire  regs_370_reset; // @[RegFile.scala 66:20:@130170.4]
  wire [63:0] regs_370_io_in; // @[RegFile.scala 66:20:@130170.4]
  wire  regs_370_io_reset; // @[RegFile.scala 66:20:@130170.4]
  wire [63:0] regs_370_io_out; // @[RegFile.scala 66:20:@130170.4]
  wire  regs_370_io_enable; // @[RegFile.scala 66:20:@130170.4]
  wire  regs_371_clock; // @[RegFile.scala 66:20:@130184.4]
  wire  regs_371_reset; // @[RegFile.scala 66:20:@130184.4]
  wire [63:0] regs_371_io_in; // @[RegFile.scala 66:20:@130184.4]
  wire  regs_371_io_reset; // @[RegFile.scala 66:20:@130184.4]
  wire [63:0] regs_371_io_out; // @[RegFile.scala 66:20:@130184.4]
  wire  regs_371_io_enable; // @[RegFile.scala 66:20:@130184.4]
  wire  regs_372_clock; // @[RegFile.scala 66:20:@130198.4]
  wire  regs_372_reset; // @[RegFile.scala 66:20:@130198.4]
  wire [63:0] regs_372_io_in; // @[RegFile.scala 66:20:@130198.4]
  wire  regs_372_io_reset; // @[RegFile.scala 66:20:@130198.4]
  wire [63:0] regs_372_io_out; // @[RegFile.scala 66:20:@130198.4]
  wire  regs_372_io_enable; // @[RegFile.scala 66:20:@130198.4]
  wire  regs_373_clock; // @[RegFile.scala 66:20:@130212.4]
  wire  regs_373_reset; // @[RegFile.scala 66:20:@130212.4]
  wire [63:0] regs_373_io_in; // @[RegFile.scala 66:20:@130212.4]
  wire  regs_373_io_reset; // @[RegFile.scala 66:20:@130212.4]
  wire [63:0] regs_373_io_out; // @[RegFile.scala 66:20:@130212.4]
  wire  regs_373_io_enable; // @[RegFile.scala 66:20:@130212.4]
  wire  regs_374_clock; // @[RegFile.scala 66:20:@130226.4]
  wire  regs_374_reset; // @[RegFile.scala 66:20:@130226.4]
  wire [63:0] regs_374_io_in; // @[RegFile.scala 66:20:@130226.4]
  wire  regs_374_io_reset; // @[RegFile.scala 66:20:@130226.4]
  wire [63:0] regs_374_io_out; // @[RegFile.scala 66:20:@130226.4]
  wire  regs_374_io_enable; // @[RegFile.scala 66:20:@130226.4]
  wire  regs_375_clock; // @[RegFile.scala 66:20:@130240.4]
  wire  regs_375_reset; // @[RegFile.scala 66:20:@130240.4]
  wire [63:0] regs_375_io_in; // @[RegFile.scala 66:20:@130240.4]
  wire  regs_375_io_reset; // @[RegFile.scala 66:20:@130240.4]
  wire [63:0] regs_375_io_out; // @[RegFile.scala 66:20:@130240.4]
  wire  regs_375_io_enable; // @[RegFile.scala 66:20:@130240.4]
  wire  regs_376_clock; // @[RegFile.scala 66:20:@130254.4]
  wire  regs_376_reset; // @[RegFile.scala 66:20:@130254.4]
  wire [63:0] regs_376_io_in; // @[RegFile.scala 66:20:@130254.4]
  wire  regs_376_io_reset; // @[RegFile.scala 66:20:@130254.4]
  wire [63:0] regs_376_io_out; // @[RegFile.scala 66:20:@130254.4]
  wire  regs_376_io_enable; // @[RegFile.scala 66:20:@130254.4]
  wire  regs_377_clock; // @[RegFile.scala 66:20:@130268.4]
  wire  regs_377_reset; // @[RegFile.scala 66:20:@130268.4]
  wire [63:0] regs_377_io_in; // @[RegFile.scala 66:20:@130268.4]
  wire  regs_377_io_reset; // @[RegFile.scala 66:20:@130268.4]
  wire [63:0] regs_377_io_out; // @[RegFile.scala 66:20:@130268.4]
  wire  regs_377_io_enable; // @[RegFile.scala 66:20:@130268.4]
  wire  regs_378_clock; // @[RegFile.scala 66:20:@130282.4]
  wire  regs_378_reset; // @[RegFile.scala 66:20:@130282.4]
  wire [63:0] regs_378_io_in; // @[RegFile.scala 66:20:@130282.4]
  wire  regs_378_io_reset; // @[RegFile.scala 66:20:@130282.4]
  wire [63:0] regs_378_io_out; // @[RegFile.scala 66:20:@130282.4]
  wire  regs_378_io_enable; // @[RegFile.scala 66:20:@130282.4]
  wire  regs_379_clock; // @[RegFile.scala 66:20:@130296.4]
  wire  regs_379_reset; // @[RegFile.scala 66:20:@130296.4]
  wire [63:0] regs_379_io_in; // @[RegFile.scala 66:20:@130296.4]
  wire  regs_379_io_reset; // @[RegFile.scala 66:20:@130296.4]
  wire [63:0] regs_379_io_out; // @[RegFile.scala 66:20:@130296.4]
  wire  regs_379_io_enable; // @[RegFile.scala 66:20:@130296.4]
  wire  regs_380_clock; // @[RegFile.scala 66:20:@130310.4]
  wire  regs_380_reset; // @[RegFile.scala 66:20:@130310.4]
  wire [63:0] regs_380_io_in; // @[RegFile.scala 66:20:@130310.4]
  wire  regs_380_io_reset; // @[RegFile.scala 66:20:@130310.4]
  wire [63:0] regs_380_io_out; // @[RegFile.scala 66:20:@130310.4]
  wire  regs_380_io_enable; // @[RegFile.scala 66:20:@130310.4]
  wire  regs_381_clock; // @[RegFile.scala 66:20:@130324.4]
  wire  regs_381_reset; // @[RegFile.scala 66:20:@130324.4]
  wire [63:0] regs_381_io_in; // @[RegFile.scala 66:20:@130324.4]
  wire  regs_381_io_reset; // @[RegFile.scala 66:20:@130324.4]
  wire [63:0] regs_381_io_out; // @[RegFile.scala 66:20:@130324.4]
  wire  regs_381_io_enable; // @[RegFile.scala 66:20:@130324.4]
  wire  regs_382_clock; // @[RegFile.scala 66:20:@130338.4]
  wire  regs_382_reset; // @[RegFile.scala 66:20:@130338.4]
  wire [63:0] regs_382_io_in; // @[RegFile.scala 66:20:@130338.4]
  wire  regs_382_io_reset; // @[RegFile.scala 66:20:@130338.4]
  wire [63:0] regs_382_io_out; // @[RegFile.scala 66:20:@130338.4]
  wire  regs_382_io_enable; // @[RegFile.scala 66:20:@130338.4]
  wire  regs_383_clock; // @[RegFile.scala 66:20:@130352.4]
  wire  regs_383_reset; // @[RegFile.scala 66:20:@130352.4]
  wire [63:0] regs_383_io_in; // @[RegFile.scala 66:20:@130352.4]
  wire  regs_383_io_reset; // @[RegFile.scala 66:20:@130352.4]
  wire [63:0] regs_383_io_out; // @[RegFile.scala 66:20:@130352.4]
  wire  regs_383_io_enable; // @[RegFile.scala 66:20:@130352.4]
  wire  regs_384_clock; // @[RegFile.scala 66:20:@130366.4]
  wire  regs_384_reset; // @[RegFile.scala 66:20:@130366.4]
  wire [63:0] regs_384_io_in; // @[RegFile.scala 66:20:@130366.4]
  wire  regs_384_io_reset; // @[RegFile.scala 66:20:@130366.4]
  wire [63:0] regs_384_io_out; // @[RegFile.scala 66:20:@130366.4]
  wire  regs_384_io_enable; // @[RegFile.scala 66:20:@130366.4]
  wire  regs_385_clock; // @[RegFile.scala 66:20:@130380.4]
  wire  regs_385_reset; // @[RegFile.scala 66:20:@130380.4]
  wire [63:0] regs_385_io_in; // @[RegFile.scala 66:20:@130380.4]
  wire  regs_385_io_reset; // @[RegFile.scala 66:20:@130380.4]
  wire [63:0] regs_385_io_out; // @[RegFile.scala 66:20:@130380.4]
  wire  regs_385_io_enable; // @[RegFile.scala 66:20:@130380.4]
  wire  regs_386_clock; // @[RegFile.scala 66:20:@130394.4]
  wire  regs_386_reset; // @[RegFile.scala 66:20:@130394.4]
  wire [63:0] regs_386_io_in; // @[RegFile.scala 66:20:@130394.4]
  wire  regs_386_io_reset; // @[RegFile.scala 66:20:@130394.4]
  wire [63:0] regs_386_io_out; // @[RegFile.scala 66:20:@130394.4]
  wire  regs_386_io_enable; // @[RegFile.scala 66:20:@130394.4]
  wire  regs_387_clock; // @[RegFile.scala 66:20:@130408.4]
  wire  regs_387_reset; // @[RegFile.scala 66:20:@130408.4]
  wire [63:0] regs_387_io_in; // @[RegFile.scala 66:20:@130408.4]
  wire  regs_387_io_reset; // @[RegFile.scala 66:20:@130408.4]
  wire [63:0] regs_387_io_out; // @[RegFile.scala 66:20:@130408.4]
  wire  regs_387_io_enable; // @[RegFile.scala 66:20:@130408.4]
  wire  regs_388_clock; // @[RegFile.scala 66:20:@130422.4]
  wire  regs_388_reset; // @[RegFile.scala 66:20:@130422.4]
  wire [63:0] regs_388_io_in; // @[RegFile.scala 66:20:@130422.4]
  wire  regs_388_io_reset; // @[RegFile.scala 66:20:@130422.4]
  wire [63:0] regs_388_io_out; // @[RegFile.scala 66:20:@130422.4]
  wire  regs_388_io_enable; // @[RegFile.scala 66:20:@130422.4]
  wire  regs_389_clock; // @[RegFile.scala 66:20:@130436.4]
  wire  regs_389_reset; // @[RegFile.scala 66:20:@130436.4]
  wire [63:0] regs_389_io_in; // @[RegFile.scala 66:20:@130436.4]
  wire  regs_389_io_reset; // @[RegFile.scala 66:20:@130436.4]
  wire [63:0] regs_389_io_out; // @[RegFile.scala 66:20:@130436.4]
  wire  regs_389_io_enable; // @[RegFile.scala 66:20:@130436.4]
  wire  regs_390_clock; // @[RegFile.scala 66:20:@130450.4]
  wire  regs_390_reset; // @[RegFile.scala 66:20:@130450.4]
  wire [63:0] regs_390_io_in; // @[RegFile.scala 66:20:@130450.4]
  wire  regs_390_io_reset; // @[RegFile.scala 66:20:@130450.4]
  wire [63:0] regs_390_io_out; // @[RegFile.scala 66:20:@130450.4]
  wire  regs_390_io_enable; // @[RegFile.scala 66:20:@130450.4]
  wire  regs_391_clock; // @[RegFile.scala 66:20:@130464.4]
  wire  regs_391_reset; // @[RegFile.scala 66:20:@130464.4]
  wire [63:0] regs_391_io_in; // @[RegFile.scala 66:20:@130464.4]
  wire  regs_391_io_reset; // @[RegFile.scala 66:20:@130464.4]
  wire [63:0] regs_391_io_out; // @[RegFile.scala 66:20:@130464.4]
  wire  regs_391_io_enable; // @[RegFile.scala 66:20:@130464.4]
  wire  regs_392_clock; // @[RegFile.scala 66:20:@130478.4]
  wire  regs_392_reset; // @[RegFile.scala 66:20:@130478.4]
  wire [63:0] regs_392_io_in; // @[RegFile.scala 66:20:@130478.4]
  wire  regs_392_io_reset; // @[RegFile.scala 66:20:@130478.4]
  wire [63:0] regs_392_io_out; // @[RegFile.scala 66:20:@130478.4]
  wire  regs_392_io_enable; // @[RegFile.scala 66:20:@130478.4]
  wire  regs_393_clock; // @[RegFile.scala 66:20:@130492.4]
  wire  regs_393_reset; // @[RegFile.scala 66:20:@130492.4]
  wire [63:0] regs_393_io_in; // @[RegFile.scala 66:20:@130492.4]
  wire  regs_393_io_reset; // @[RegFile.scala 66:20:@130492.4]
  wire [63:0] regs_393_io_out; // @[RegFile.scala 66:20:@130492.4]
  wire  regs_393_io_enable; // @[RegFile.scala 66:20:@130492.4]
  wire  regs_394_clock; // @[RegFile.scala 66:20:@130506.4]
  wire  regs_394_reset; // @[RegFile.scala 66:20:@130506.4]
  wire [63:0] regs_394_io_in; // @[RegFile.scala 66:20:@130506.4]
  wire  regs_394_io_reset; // @[RegFile.scala 66:20:@130506.4]
  wire [63:0] regs_394_io_out; // @[RegFile.scala 66:20:@130506.4]
  wire  regs_394_io_enable; // @[RegFile.scala 66:20:@130506.4]
  wire  regs_395_clock; // @[RegFile.scala 66:20:@130520.4]
  wire  regs_395_reset; // @[RegFile.scala 66:20:@130520.4]
  wire [63:0] regs_395_io_in; // @[RegFile.scala 66:20:@130520.4]
  wire  regs_395_io_reset; // @[RegFile.scala 66:20:@130520.4]
  wire [63:0] regs_395_io_out; // @[RegFile.scala 66:20:@130520.4]
  wire  regs_395_io_enable; // @[RegFile.scala 66:20:@130520.4]
  wire  regs_396_clock; // @[RegFile.scala 66:20:@130534.4]
  wire  regs_396_reset; // @[RegFile.scala 66:20:@130534.4]
  wire [63:0] regs_396_io_in; // @[RegFile.scala 66:20:@130534.4]
  wire  regs_396_io_reset; // @[RegFile.scala 66:20:@130534.4]
  wire [63:0] regs_396_io_out; // @[RegFile.scala 66:20:@130534.4]
  wire  regs_396_io_enable; // @[RegFile.scala 66:20:@130534.4]
  wire  regs_397_clock; // @[RegFile.scala 66:20:@130548.4]
  wire  regs_397_reset; // @[RegFile.scala 66:20:@130548.4]
  wire [63:0] regs_397_io_in; // @[RegFile.scala 66:20:@130548.4]
  wire  regs_397_io_reset; // @[RegFile.scala 66:20:@130548.4]
  wire [63:0] regs_397_io_out; // @[RegFile.scala 66:20:@130548.4]
  wire  regs_397_io_enable; // @[RegFile.scala 66:20:@130548.4]
  wire  regs_398_clock; // @[RegFile.scala 66:20:@130562.4]
  wire  regs_398_reset; // @[RegFile.scala 66:20:@130562.4]
  wire [63:0] regs_398_io_in; // @[RegFile.scala 66:20:@130562.4]
  wire  regs_398_io_reset; // @[RegFile.scala 66:20:@130562.4]
  wire [63:0] regs_398_io_out; // @[RegFile.scala 66:20:@130562.4]
  wire  regs_398_io_enable; // @[RegFile.scala 66:20:@130562.4]
  wire  regs_399_clock; // @[RegFile.scala 66:20:@130576.4]
  wire  regs_399_reset; // @[RegFile.scala 66:20:@130576.4]
  wire [63:0] regs_399_io_in; // @[RegFile.scala 66:20:@130576.4]
  wire  regs_399_io_reset; // @[RegFile.scala 66:20:@130576.4]
  wire [63:0] regs_399_io_out; // @[RegFile.scala 66:20:@130576.4]
  wire  regs_399_io_enable; // @[RegFile.scala 66:20:@130576.4]
  wire  regs_400_clock; // @[RegFile.scala 66:20:@130590.4]
  wire  regs_400_reset; // @[RegFile.scala 66:20:@130590.4]
  wire [63:0] regs_400_io_in; // @[RegFile.scala 66:20:@130590.4]
  wire  regs_400_io_reset; // @[RegFile.scala 66:20:@130590.4]
  wire [63:0] regs_400_io_out; // @[RegFile.scala 66:20:@130590.4]
  wire  regs_400_io_enable; // @[RegFile.scala 66:20:@130590.4]
  wire  regs_401_clock; // @[RegFile.scala 66:20:@130604.4]
  wire  regs_401_reset; // @[RegFile.scala 66:20:@130604.4]
  wire [63:0] regs_401_io_in; // @[RegFile.scala 66:20:@130604.4]
  wire  regs_401_io_reset; // @[RegFile.scala 66:20:@130604.4]
  wire [63:0] regs_401_io_out; // @[RegFile.scala 66:20:@130604.4]
  wire  regs_401_io_enable; // @[RegFile.scala 66:20:@130604.4]
  wire  regs_402_clock; // @[RegFile.scala 66:20:@130618.4]
  wire  regs_402_reset; // @[RegFile.scala 66:20:@130618.4]
  wire [63:0] regs_402_io_in; // @[RegFile.scala 66:20:@130618.4]
  wire  regs_402_io_reset; // @[RegFile.scala 66:20:@130618.4]
  wire [63:0] regs_402_io_out; // @[RegFile.scala 66:20:@130618.4]
  wire  regs_402_io_enable; // @[RegFile.scala 66:20:@130618.4]
  wire  regs_403_clock; // @[RegFile.scala 66:20:@130632.4]
  wire  regs_403_reset; // @[RegFile.scala 66:20:@130632.4]
  wire [63:0] regs_403_io_in; // @[RegFile.scala 66:20:@130632.4]
  wire  regs_403_io_reset; // @[RegFile.scala 66:20:@130632.4]
  wire [63:0] regs_403_io_out; // @[RegFile.scala 66:20:@130632.4]
  wire  regs_403_io_enable; // @[RegFile.scala 66:20:@130632.4]
  wire  regs_404_clock; // @[RegFile.scala 66:20:@130646.4]
  wire  regs_404_reset; // @[RegFile.scala 66:20:@130646.4]
  wire [63:0] regs_404_io_in; // @[RegFile.scala 66:20:@130646.4]
  wire  regs_404_io_reset; // @[RegFile.scala 66:20:@130646.4]
  wire [63:0] regs_404_io_out; // @[RegFile.scala 66:20:@130646.4]
  wire  regs_404_io_enable; // @[RegFile.scala 66:20:@130646.4]
  wire  regs_405_clock; // @[RegFile.scala 66:20:@130660.4]
  wire  regs_405_reset; // @[RegFile.scala 66:20:@130660.4]
  wire [63:0] regs_405_io_in; // @[RegFile.scala 66:20:@130660.4]
  wire  regs_405_io_reset; // @[RegFile.scala 66:20:@130660.4]
  wire [63:0] regs_405_io_out; // @[RegFile.scala 66:20:@130660.4]
  wire  regs_405_io_enable; // @[RegFile.scala 66:20:@130660.4]
  wire  regs_406_clock; // @[RegFile.scala 66:20:@130674.4]
  wire  regs_406_reset; // @[RegFile.scala 66:20:@130674.4]
  wire [63:0] regs_406_io_in; // @[RegFile.scala 66:20:@130674.4]
  wire  regs_406_io_reset; // @[RegFile.scala 66:20:@130674.4]
  wire [63:0] regs_406_io_out; // @[RegFile.scala 66:20:@130674.4]
  wire  regs_406_io_enable; // @[RegFile.scala 66:20:@130674.4]
  wire  regs_407_clock; // @[RegFile.scala 66:20:@130688.4]
  wire  regs_407_reset; // @[RegFile.scala 66:20:@130688.4]
  wire [63:0] regs_407_io_in; // @[RegFile.scala 66:20:@130688.4]
  wire  regs_407_io_reset; // @[RegFile.scala 66:20:@130688.4]
  wire [63:0] regs_407_io_out; // @[RegFile.scala 66:20:@130688.4]
  wire  regs_407_io_enable; // @[RegFile.scala 66:20:@130688.4]
  wire  regs_408_clock; // @[RegFile.scala 66:20:@130702.4]
  wire  regs_408_reset; // @[RegFile.scala 66:20:@130702.4]
  wire [63:0] regs_408_io_in; // @[RegFile.scala 66:20:@130702.4]
  wire  regs_408_io_reset; // @[RegFile.scala 66:20:@130702.4]
  wire [63:0] regs_408_io_out; // @[RegFile.scala 66:20:@130702.4]
  wire  regs_408_io_enable; // @[RegFile.scala 66:20:@130702.4]
  wire  regs_409_clock; // @[RegFile.scala 66:20:@130716.4]
  wire  regs_409_reset; // @[RegFile.scala 66:20:@130716.4]
  wire [63:0] regs_409_io_in; // @[RegFile.scala 66:20:@130716.4]
  wire  regs_409_io_reset; // @[RegFile.scala 66:20:@130716.4]
  wire [63:0] regs_409_io_out; // @[RegFile.scala 66:20:@130716.4]
  wire  regs_409_io_enable; // @[RegFile.scala 66:20:@130716.4]
  wire  regs_410_clock; // @[RegFile.scala 66:20:@130730.4]
  wire  regs_410_reset; // @[RegFile.scala 66:20:@130730.4]
  wire [63:0] regs_410_io_in; // @[RegFile.scala 66:20:@130730.4]
  wire  regs_410_io_reset; // @[RegFile.scala 66:20:@130730.4]
  wire [63:0] regs_410_io_out; // @[RegFile.scala 66:20:@130730.4]
  wire  regs_410_io_enable; // @[RegFile.scala 66:20:@130730.4]
  wire  regs_411_clock; // @[RegFile.scala 66:20:@130744.4]
  wire  regs_411_reset; // @[RegFile.scala 66:20:@130744.4]
  wire [63:0] regs_411_io_in; // @[RegFile.scala 66:20:@130744.4]
  wire  regs_411_io_reset; // @[RegFile.scala 66:20:@130744.4]
  wire [63:0] regs_411_io_out; // @[RegFile.scala 66:20:@130744.4]
  wire  regs_411_io_enable; // @[RegFile.scala 66:20:@130744.4]
  wire  regs_412_clock; // @[RegFile.scala 66:20:@130758.4]
  wire  regs_412_reset; // @[RegFile.scala 66:20:@130758.4]
  wire [63:0] regs_412_io_in; // @[RegFile.scala 66:20:@130758.4]
  wire  regs_412_io_reset; // @[RegFile.scala 66:20:@130758.4]
  wire [63:0] regs_412_io_out; // @[RegFile.scala 66:20:@130758.4]
  wire  regs_412_io_enable; // @[RegFile.scala 66:20:@130758.4]
  wire  regs_413_clock; // @[RegFile.scala 66:20:@130772.4]
  wire  regs_413_reset; // @[RegFile.scala 66:20:@130772.4]
  wire [63:0] regs_413_io_in; // @[RegFile.scala 66:20:@130772.4]
  wire  regs_413_io_reset; // @[RegFile.scala 66:20:@130772.4]
  wire [63:0] regs_413_io_out; // @[RegFile.scala 66:20:@130772.4]
  wire  regs_413_io_enable; // @[RegFile.scala 66:20:@130772.4]
  wire  regs_414_clock; // @[RegFile.scala 66:20:@130786.4]
  wire  regs_414_reset; // @[RegFile.scala 66:20:@130786.4]
  wire [63:0] regs_414_io_in; // @[RegFile.scala 66:20:@130786.4]
  wire  regs_414_io_reset; // @[RegFile.scala 66:20:@130786.4]
  wire [63:0] regs_414_io_out; // @[RegFile.scala 66:20:@130786.4]
  wire  regs_414_io_enable; // @[RegFile.scala 66:20:@130786.4]
  wire  regs_415_clock; // @[RegFile.scala 66:20:@130800.4]
  wire  regs_415_reset; // @[RegFile.scala 66:20:@130800.4]
  wire [63:0] regs_415_io_in; // @[RegFile.scala 66:20:@130800.4]
  wire  regs_415_io_reset; // @[RegFile.scala 66:20:@130800.4]
  wire [63:0] regs_415_io_out; // @[RegFile.scala 66:20:@130800.4]
  wire  regs_415_io_enable; // @[RegFile.scala 66:20:@130800.4]
  wire  regs_416_clock; // @[RegFile.scala 66:20:@130814.4]
  wire  regs_416_reset; // @[RegFile.scala 66:20:@130814.4]
  wire [63:0] regs_416_io_in; // @[RegFile.scala 66:20:@130814.4]
  wire  regs_416_io_reset; // @[RegFile.scala 66:20:@130814.4]
  wire [63:0] regs_416_io_out; // @[RegFile.scala 66:20:@130814.4]
  wire  regs_416_io_enable; // @[RegFile.scala 66:20:@130814.4]
  wire  regs_417_clock; // @[RegFile.scala 66:20:@130828.4]
  wire  regs_417_reset; // @[RegFile.scala 66:20:@130828.4]
  wire [63:0] regs_417_io_in; // @[RegFile.scala 66:20:@130828.4]
  wire  regs_417_io_reset; // @[RegFile.scala 66:20:@130828.4]
  wire [63:0] regs_417_io_out; // @[RegFile.scala 66:20:@130828.4]
  wire  regs_417_io_enable; // @[RegFile.scala 66:20:@130828.4]
  wire  regs_418_clock; // @[RegFile.scala 66:20:@130842.4]
  wire  regs_418_reset; // @[RegFile.scala 66:20:@130842.4]
  wire [63:0] regs_418_io_in; // @[RegFile.scala 66:20:@130842.4]
  wire  regs_418_io_reset; // @[RegFile.scala 66:20:@130842.4]
  wire [63:0] regs_418_io_out; // @[RegFile.scala 66:20:@130842.4]
  wire  regs_418_io_enable; // @[RegFile.scala 66:20:@130842.4]
  wire  regs_419_clock; // @[RegFile.scala 66:20:@130856.4]
  wire  regs_419_reset; // @[RegFile.scala 66:20:@130856.4]
  wire [63:0] regs_419_io_in; // @[RegFile.scala 66:20:@130856.4]
  wire  regs_419_io_reset; // @[RegFile.scala 66:20:@130856.4]
  wire [63:0] regs_419_io_out; // @[RegFile.scala 66:20:@130856.4]
  wire  regs_419_io_enable; // @[RegFile.scala 66:20:@130856.4]
  wire  regs_420_clock; // @[RegFile.scala 66:20:@130870.4]
  wire  regs_420_reset; // @[RegFile.scala 66:20:@130870.4]
  wire [63:0] regs_420_io_in; // @[RegFile.scala 66:20:@130870.4]
  wire  regs_420_io_reset; // @[RegFile.scala 66:20:@130870.4]
  wire [63:0] regs_420_io_out; // @[RegFile.scala 66:20:@130870.4]
  wire  regs_420_io_enable; // @[RegFile.scala 66:20:@130870.4]
  wire  regs_421_clock; // @[RegFile.scala 66:20:@130884.4]
  wire  regs_421_reset; // @[RegFile.scala 66:20:@130884.4]
  wire [63:0] regs_421_io_in; // @[RegFile.scala 66:20:@130884.4]
  wire  regs_421_io_reset; // @[RegFile.scala 66:20:@130884.4]
  wire [63:0] regs_421_io_out; // @[RegFile.scala 66:20:@130884.4]
  wire  regs_421_io_enable; // @[RegFile.scala 66:20:@130884.4]
  wire  regs_422_clock; // @[RegFile.scala 66:20:@130898.4]
  wire  regs_422_reset; // @[RegFile.scala 66:20:@130898.4]
  wire [63:0] regs_422_io_in; // @[RegFile.scala 66:20:@130898.4]
  wire  regs_422_io_reset; // @[RegFile.scala 66:20:@130898.4]
  wire [63:0] regs_422_io_out; // @[RegFile.scala 66:20:@130898.4]
  wire  regs_422_io_enable; // @[RegFile.scala 66:20:@130898.4]
  wire  regs_423_clock; // @[RegFile.scala 66:20:@130912.4]
  wire  regs_423_reset; // @[RegFile.scala 66:20:@130912.4]
  wire [63:0] regs_423_io_in; // @[RegFile.scala 66:20:@130912.4]
  wire  regs_423_io_reset; // @[RegFile.scala 66:20:@130912.4]
  wire [63:0] regs_423_io_out; // @[RegFile.scala 66:20:@130912.4]
  wire  regs_423_io_enable; // @[RegFile.scala 66:20:@130912.4]
  wire  regs_424_clock; // @[RegFile.scala 66:20:@130926.4]
  wire  regs_424_reset; // @[RegFile.scala 66:20:@130926.4]
  wire [63:0] regs_424_io_in; // @[RegFile.scala 66:20:@130926.4]
  wire  regs_424_io_reset; // @[RegFile.scala 66:20:@130926.4]
  wire [63:0] regs_424_io_out; // @[RegFile.scala 66:20:@130926.4]
  wire  regs_424_io_enable; // @[RegFile.scala 66:20:@130926.4]
  wire  regs_425_clock; // @[RegFile.scala 66:20:@130940.4]
  wire  regs_425_reset; // @[RegFile.scala 66:20:@130940.4]
  wire [63:0] regs_425_io_in; // @[RegFile.scala 66:20:@130940.4]
  wire  regs_425_io_reset; // @[RegFile.scala 66:20:@130940.4]
  wire [63:0] regs_425_io_out; // @[RegFile.scala 66:20:@130940.4]
  wire  regs_425_io_enable; // @[RegFile.scala 66:20:@130940.4]
  wire  regs_426_clock; // @[RegFile.scala 66:20:@130954.4]
  wire  regs_426_reset; // @[RegFile.scala 66:20:@130954.4]
  wire [63:0] regs_426_io_in; // @[RegFile.scala 66:20:@130954.4]
  wire  regs_426_io_reset; // @[RegFile.scala 66:20:@130954.4]
  wire [63:0] regs_426_io_out; // @[RegFile.scala 66:20:@130954.4]
  wire  regs_426_io_enable; // @[RegFile.scala 66:20:@130954.4]
  wire  regs_427_clock; // @[RegFile.scala 66:20:@130968.4]
  wire  regs_427_reset; // @[RegFile.scala 66:20:@130968.4]
  wire [63:0] regs_427_io_in; // @[RegFile.scala 66:20:@130968.4]
  wire  regs_427_io_reset; // @[RegFile.scala 66:20:@130968.4]
  wire [63:0] regs_427_io_out; // @[RegFile.scala 66:20:@130968.4]
  wire  regs_427_io_enable; // @[RegFile.scala 66:20:@130968.4]
  wire  regs_428_clock; // @[RegFile.scala 66:20:@130982.4]
  wire  regs_428_reset; // @[RegFile.scala 66:20:@130982.4]
  wire [63:0] regs_428_io_in; // @[RegFile.scala 66:20:@130982.4]
  wire  regs_428_io_reset; // @[RegFile.scala 66:20:@130982.4]
  wire [63:0] regs_428_io_out; // @[RegFile.scala 66:20:@130982.4]
  wire  regs_428_io_enable; // @[RegFile.scala 66:20:@130982.4]
  wire  regs_429_clock; // @[RegFile.scala 66:20:@130996.4]
  wire  regs_429_reset; // @[RegFile.scala 66:20:@130996.4]
  wire [63:0] regs_429_io_in; // @[RegFile.scala 66:20:@130996.4]
  wire  regs_429_io_reset; // @[RegFile.scala 66:20:@130996.4]
  wire [63:0] regs_429_io_out; // @[RegFile.scala 66:20:@130996.4]
  wire  regs_429_io_enable; // @[RegFile.scala 66:20:@130996.4]
  wire  regs_430_clock; // @[RegFile.scala 66:20:@131010.4]
  wire  regs_430_reset; // @[RegFile.scala 66:20:@131010.4]
  wire [63:0] regs_430_io_in; // @[RegFile.scala 66:20:@131010.4]
  wire  regs_430_io_reset; // @[RegFile.scala 66:20:@131010.4]
  wire [63:0] regs_430_io_out; // @[RegFile.scala 66:20:@131010.4]
  wire  regs_430_io_enable; // @[RegFile.scala 66:20:@131010.4]
  wire  regs_431_clock; // @[RegFile.scala 66:20:@131024.4]
  wire  regs_431_reset; // @[RegFile.scala 66:20:@131024.4]
  wire [63:0] regs_431_io_in; // @[RegFile.scala 66:20:@131024.4]
  wire  regs_431_io_reset; // @[RegFile.scala 66:20:@131024.4]
  wire [63:0] regs_431_io_out; // @[RegFile.scala 66:20:@131024.4]
  wire  regs_431_io_enable; // @[RegFile.scala 66:20:@131024.4]
  wire  regs_432_clock; // @[RegFile.scala 66:20:@131038.4]
  wire  regs_432_reset; // @[RegFile.scala 66:20:@131038.4]
  wire [63:0] regs_432_io_in; // @[RegFile.scala 66:20:@131038.4]
  wire  regs_432_io_reset; // @[RegFile.scala 66:20:@131038.4]
  wire [63:0] regs_432_io_out; // @[RegFile.scala 66:20:@131038.4]
  wire  regs_432_io_enable; // @[RegFile.scala 66:20:@131038.4]
  wire  regs_433_clock; // @[RegFile.scala 66:20:@131052.4]
  wire  regs_433_reset; // @[RegFile.scala 66:20:@131052.4]
  wire [63:0] regs_433_io_in; // @[RegFile.scala 66:20:@131052.4]
  wire  regs_433_io_reset; // @[RegFile.scala 66:20:@131052.4]
  wire [63:0] regs_433_io_out; // @[RegFile.scala 66:20:@131052.4]
  wire  regs_433_io_enable; // @[RegFile.scala 66:20:@131052.4]
  wire  regs_434_clock; // @[RegFile.scala 66:20:@131066.4]
  wire  regs_434_reset; // @[RegFile.scala 66:20:@131066.4]
  wire [63:0] regs_434_io_in; // @[RegFile.scala 66:20:@131066.4]
  wire  regs_434_io_reset; // @[RegFile.scala 66:20:@131066.4]
  wire [63:0] regs_434_io_out; // @[RegFile.scala 66:20:@131066.4]
  wire  regs_434_io_enable; // @[RegFile.scala 66:20:@131066.4]
  wire  regs_435_clock; // @[RegFile.scala 66:20:@131080.4]
  wire  regs_435_reset; // @[RegFile.scala 66:20:@131080.4]
  wire [63:0] regs_435_io_in; // @[RegFile.scala 66:20:@131080.4]
  wire  regs_435_io_reset; // @[RegFile.scala 66:20:@131080.4]
  wire [63:0] regs_435_io_out; // @[RegFile.scala 66:20:@131080.4]
  wire  regs_435_io_enable; // @[RegFile.scala 66:20:@131080.4]
  wire  regs_436_clock; // @[RegFile.scala 66:20:@131094.4]
  wire  regs_436_reset; // @[RegFile.scala 66:20:@131094.4]
  wire [63:0] regs_436_io_in; // @[RegFile.scala 66:20:@131094.4]
  wire  regs_436_io_reset; // @[RegFile.scala 66:20:@131094.4]
  wire [63:0] regs_436_io_out; // @[RegFile.scala 66:20:@131094.4]
  wire  regs_436_io_enable; // @[RegFile.scala 66:20:@131094.4]
  wire  regs_437_clock; // @[RegFile.scala 66:20:@131108.4]
  wire  regs_437_reset; // @[RegFile.scala 66:20:@131108.4]
  wire [63:0] regs_437_io_in; // @[RegFile.scala 66:20:@131108.4]
  wire  regs_437_io_reset; // @[RegFile.scala 66:20:@131108.4]
  wire [63:0] regs_437_io_out; // @[RegFile.scala 66:20:@131108.4]
  wire  regs_437_io_enable; // @[RegFile.scala 66:20:@131108.4]
  wire  regs_438_clock; // @[RegFile.scala 66:20:@131122.4]
  wire  regs_438_reset; // @[RegFile.scala 66:20:@131122.4]
  wire [63:0] regs_438_io_in; // @[RegFile.scala 66:20:@131122.4]
  wire  regs_438_io_reset; // @[RegFile.scala 66:20:@131122.4]
  wire [63:0] regs_438_io_out; // @[RegFile.scala 66:20:@131122.4]
  wire  regs_438_io_enable; // @[RegFile.scala 66:20:@131122.4]
  wire  regs_439_clock; // @[RegFile.scala 66:20:@131136.4]
  wire  regs_439_reset; // @[RegFile.scala 66:20:@131136.4]
  wire [63:0] regs_439_io_in; // @[RegFile.scala 66:20:@131136.4]
  wire  regs_439_io_reset; // @[RegFile.scala 66:20:@131136.4]
  wire [63:0] regs_439_io_out; // @[RegFile.scala 66:20:@131136.4]
  wire  regs_439_io_enable; // @[RegFile.scala 66:20:@131136.4]
  wire  regs_440_clock; // @[RegFile.scala 66:20:@131150.4]
  wire  regs_440_reset; // @[RegFile.scala 66:20:@131150.4]
  wire [63:0] regs_440_io_in; // @[RegFile.scala 66:20:@131150.4]
  wire  regs_440_io_reset; // @[RegFile.scala 66:20:@131150.4]
  wire [63:0] regs_440_io_out; // @[RegFile.scala 66:20:@131150.4]
  wire  regs_440_io_enable; // @[RegFile.scala 66:20:@131150.4]
  wire  regs_441_clock; // @[RegFile.scala 66:20:@131164.4]
  wire  regs_441_reset; // @[RegFile.scala 66:20:@131164.4]
  wire [63:0] regs_441_io_in; // @[RegFile.scala 66:20:@131164.4]
  wire  regs_441_io_reset; // @[RegFile.scala 66:20:@131164.4]
  wire [63:0] regs_441_io_out; // @[RegFile.scala 66:20:@131164.4]
  wire  regs_441_io_enable; // @[RegFile.scala 66:20:@131164.4]
  wire  regs_442_clock; // @[RegFile.scala 66:20:@131178.4]
  wire  regs_442_reset; // @[RegFile.scala 66:20:@131178.4]
  wire [63:0] regs_442_io_in; // @[RegFile.scala 66:20:@131178.4]
  wire  regs_442_io_reset; // @[RegFile.scala 66:20:@131178.4]
  wire [63:0] regs_442_io_out; // @[RegFile.scala 66:20:@131178.4]
  wire  regs_442_io_enable; // @[RegFile.scala 66:20:@131178.4]
  wire  regs_443_clock; // @[RegFile.scala 66:20:@131192.4]
  wire  regs_443_reset; // @[RegFile.scala 66:20:@131192.4]
  wire [63:0] regs_443_io_in; // @[RegFile.scala 66:20:@131192.4]
  wire  regs_443_io_reset; // @[RegFile.scala 66:20:@131192.4]
  wire [63:0] regs_443_io_out; // @[RegFile.scala 66:20:@131192.4]
  wire  regs_443_io_enable; // @[RegFile.scala 66:20:@131192.4]
  wire  regs_444_clock; // @[RegFile.scala 66:20:@131206.4]
  wire  regs_444_reset; // @[RegFile.scala 66:20:@131206.4]
  wire [63:0] regs_444_io_in; // @[RegFile.scala 66:20:@131206.4]
  wire  regs_444_io_reset; // @[RegFile.scala 66:20:@131206.4]
  wire [63:0] regs_444_io_out; // @[RegFile.scala 66:20:@131206.4]
  wire  regs_444_io_enable; // @[RegFile.scala 66:20:@131206.4]
  wire  regs_445_clock; // @[RegFile.scala 66:20:@131220.4]
  wire  regs_445_reset; // @[RegFile.scala 66:20:@131220.4]
  wire [63:0] regs_445_io_in; // @[RegFile.scala 66:20:@131220.4]
  wire  regs_445_io_reset; // @[RegFile.scala 66:20:@131220.4]
  wire [63:0] regs_445_io_out; // @[RegFile.scala 66:20:@131220.4]
  wire  regs_445_io_enable; // @[RegFile.scala 66:20:@131220.4]
  wire  regs_446_clock; // @[RegFile.scala 66:20:@131234.4]
  wire  regs_446_reset; // @[RegFile.scala 66:20:@131234.4]
  wire [63:0] regs_446_io_in; // @[RegFile.scala 66:20:@131234.4]
  wire  regs_446_io_reset; // @[RegFile.scala 66:20:@131234.4]
  wire [63:0] regs_446_io_out; // @[RegFile.scala 66:20:@131234.4]
  wire  regs_446_io_enable; // @[RegFile.scala 66:20:@131234.4]
  wire  regs_447_clock; // @[RegFile.scala 66:20:@131248.4]
  wire  regs_447_reset; // @[RegFile.scala 66:20:@131248.4]
  wire [63:0] regs_447_io_in; // @[RegFile.scala 66:20:@131248.4]
  wire  regs_447_io_reset; // @[RegFile.scala 66:20:@131248.4]
  wire [63:0] regs_447_io_out; // @[RegFile.scala 66:20:@131248.4]
  wire  regs_447_io_enable; // @[RegFile.scala 66:20:@131248.4]
  wire  regs_448_clock; // @[RegFile.scala 66:20:@131262.4]
  wire  regs_448_reset; // @[RegFile.scala 66:20:@131262.4]
  wire [63:0] regs_448_io_in; // @[RegFile.scala 66:20:@131262.4]
  wire  regs_448_io_reset; // @[RegFile.scala 66:20:@131262.4]
  wire [63:0] regs_448_io_out; // @[RegFile.scala 66:20:@131262.4]
  wire  regs_448_io_enable; // @[RegFile.scala 66:20:@131262.4]
  wire  regs_449_clock; // @[RegFile.scala 66:20:@131276.4]
  wire  regs_449_reset; // @[RegFile.scala 66:20:@131276.4]
  wire [63:0] regs_449_io_in; // @[RegFile.scala 66:20:@131276.4]
  wire  regs_449_io_reset; // @[RegFile.scala 66:20:@131276.4]
  wire [63:0] regs_449_io_out; // @[RegFile.scala 66:20:@131276.4]
  wire  regs_449_io_enable; // @[RegFile.scala 66:20:@131276.4]
  wire  regs_450_clock; // @[RegFile.scala 66:20:@131290.4]
  wire  regs_450_reset; // @[RegFile.scala 66:20:@131290.4]
  wire [63:0] regs_450_io_in; // @[RegFile.scala 66:20:@131290.4]
  wire  regs_450_io_reset; // @[RegFile.scala 66:20:@131290.4]
  wire [63:0] regs_450_io_out; // @[RegFile.scala 66:20:@131290.4]
  wire  regs_450_io_enable; // @[RegFile.scala 66:20:@131290.4]
  wire  regs_451_clock; // @[RegFile.scala 66:20:@131304.4]
  wire  regs_451_reset; // @[RegFile.scala 66:20:@131304.4]
  wire [63:0] regs_451_io_in; // @[RegFile.scala 66:20:@131304.4]
  wire  regs_451_io_reset; // @[RegFile.scala 66:20:@131304.4]
  wire [63:0] regs_451_io_out; // @[RegFile.scala 66:20:@131304.4]
  wire  regs_451_io_enable; // @[RegFile.scala 66:20:@131304.4]
  wire  regs_452_clock; // @[RegFile.scala 66:20:@131318.4]
  wire  regs_452_reset; // @[RegFile.scala 66:20:@131318.4]
  wire [63:0] regs_452_io_in; // @[RegFile.scala 66:20:@131318.4]
  wire  regs_452_io_reset; // @[RegFile.scala 66:20:@131318.4]
  wire [63:0] regs_452_io_out; // @[RegFile.scala 66:20:@131318.4]
  wire  regs_452_io_enable; // @[RegFile.scala 66:20:@131318.4]
  wire  regs_453_clock; // @[RegFile.scala 66:20:@131332.4]
  wire  regs_453_reset; // @[RegFile.scala 66:20:@131332.4]
  wire [63:0] regs_453_io_in; // @[RegFile.scala 66:20:@131332.4]
  wire  regs_453_io_reset; // @[RegFile.scala 66:20:@131332.4]
  wire [63:0] regs_453_io_out; // @[RegFile.scala 66:20:@131332.4]
  wire  regs_453_io_enable; // @[RegFile.scala 66:20:@131332.4]
  wire  regs_454_clock; // @[RegFile.scala 66:20:@131346.4]
  wire  regs_454_reset; // @[RegFile.scala 66:20:@131346.4]
  wire [63:0] regs_454_io_in; // @[RegFile.scala 66:20:@131346.4]
  wire  regs_454_io_reset; // @[RegFile.scala 66:20:@131346.4]
  wire [63:0] regs_454_io_out; // @[RegFile.scala 66:20:@131346.4]
  wire  regs_454_io_enable; // @[RegFile.scala 66:20:@131346.4]
  wire  regs_455_clock; // @[RegFile.scala 66:20:@131360.4]
  wire  regs_455_reset; // @[RegFile.scala 66:20:@131360.4]
  wire [63:0] regs_455_io_in; // @[RegFile.scala 66:20:@131360.4]
  wire  regs_455_io_reset; // @[RegFile.scala 66:20:@131360.4]
  wire [63:0] regs_455_io_out; // @[RegFile.scala 66:20:@131360.4]
  wire  regs_455_io_enable; // @[RegFile.scala 66:20:@131360.4]
  wire  regs_456_clock; // @[RegFile.scala 66:20:@131374.4]
  wire  regs_456_reset; // @[RegFile.scala 66:20:@131374.4]
  wire [63:0] regs_456_io_in; // @[RegFile.scala 66:20:@131374.4]
  wire  regs_456_io_reset; // @[RegFile.scala 66:20:@131374.4]
  wire [63:0] regs_456_io_out; // @[RegFile.scala 66:20:@131374.4]
  wire  regs_456_io_enable; // @[RegFile.scala 66:20:@131374.4]
  wire  regs_457_clock; // @[RegFile.scala 66:20:@131388.4]
  wire  regs_457_reset; // @[RegFile.scala 66:20:@131388.4]
  wire [63:0] regs_457_io_in; // @[RegFile.scala 66:20:@131388.4]
  wire  regs_457_io_reset; // @[RegFile.scala 66:20:@131388.4]
  wire [63:0] regs_457_io_out; // @[RegFile.scala 66:20:@131388.4]
  wire  regs_457_io_enable; // @[RegFile.scala 66:20:@131388.4]
  wire  regs_458_clock; // @[RegFile.scala 66:20:@131402.4]
  wire  regs_458_reset; // @[RegFile.scala 66:20:@131402.4]
  wire [63:0] regs_458_io_in; // @[RegFile.scala 66:20:@131402.4]
  wire  regs_458_io_reset; // @[RegFile.scala 66:20:@131402.4]
  wire [63:0] regs_458_io_out; // @[RegFile.scala 66:20:@131402.4]
  wire  regs_458_io_enable; // @[RegFile.scala 66:20:@131402.4]
  wire  regs_459_clock; // @[RegFile.scala 66:20:@131416.4]
  wire  regs_459_reset; // @[RegFile.scala 66:20:@131416.4]
  wire [63:0] regs_459_io_in; // @[RegFile.scala 66:20:@131416.4]
  wire  regs_459_io_reset; // @[RegFile.scala 66:20:@131416.4]
  wire [63:0] regs_459_io_out; // @[RegFile.scala 66:20:@131416.4]
  wire  regs_459_io_enable; // @[RegFile.scala 66:20:@131416.4]
  wire  regs_460_clock; // @[RegFile.scala 66:20:@131430.4]
  wire  regs_460_reset; // @[RegFile.scala 66:20:@131430.4]
  wire [63:0] regs_460_io_in; // @[RegFile.scala 66:20:@131430.4]
  wire  regs_460_io_reset; // @[RegFile.scala 66:20:@131430.4]
  wire [63:0] regs_460_io_out; // @[RegFile.scala 66:20:@131430.4]
  wire  regs_460_io_enable; // @[RegFile.scala 66:20:@131430.4]
  wire  regs_461_clock; // @[RegFile.scala 66:20:@131444.4]
  wire  regs_461_reset; // @[RegFile.scala 66:20:@131444.4]
  wire [63:0] regs_461_io_in; // @[RegFile.scala 66:20:@131444.4]
  wire  regs_461_io_reset; // @[RegFile.scala 66:20:@131444.4]
  wire [63:0] regs_461_io_out; // @[RegFile.scala 66:20:@131444.4]
  wire  regs_461_io_enable; // @[RegFile.scala 66:20:@131444.4]
  wire  regs_462_clock; // @[RegFile.scala 66:20:@131458.4]
  wire  regs_462_reset; // @[RegFile.scala 66:20:@131458.4]
  wire [63:0] regs_462_io_in; // @[RegFile.scala 66:20:@131458.4]
  wire  regs_462_io_reset; // @[RegFile.scala 66:20:@131458.4]
  wire [63:0] regs_462_io_out; // @[RegFile.scala 66:20:@131458.4]
  wire  regs_462_io_enable; // @[RegFile.scala 66:20:@131458.4]
  wire  regs_463_clock; // @[RegFile.scala 66:20:@131472.4]
  wire  regs_463_reset; // @[RegFile.scala 66:20:@131472.4]
  wire [63:0] regs_463_io_in; // @[RegFile.scala 66:20:@131472.4]
  wire  regs_463_io_reset; // @[RegFile.scala 66:20:@131472.4]
  wire [63:0] regs_463_io_out; // @[RegFile.scala 66:20:@131472.4]
  wire  regs_463_io_enable; // @[RegFile.scala 66:20:@131472.4]
  wire  regs_464_clock; // @[RegFile.scala 66:20:@131486.4]
  wire  regs_464_reset; // @[RegFile.scala 66:20:@131486.4]
  wire [63:0] regs_464_io_in; // @[RegFile.scala 66:20:@131486.4]
  wire  regs_464_io_reset; // @[RegFile.scala 66:20:@131486.4]
  wire [63:0] regs_464_io_out; // @[RegFile.scala 66:20:@131486.4]
  wire  regs_464_io_enable; // @[RegFile.scala 66:20:@131486.4]
  wire  regs_465_clock; // @[RegFile.scala 66:20:@131500.4]
  wire  regs_465_reset; // @[RegFile.scala 66:20:@131500.4]
  wire [63:0] regs_465_io_in; // @[RegFile.scala 66:20:@131500.4]
  wire  regs_465_io_reset; // @[RegFile.scala 66:20:@131500.4]
  wire [63:0] regs_465_io_out; // @[RegFile.scala 66:20:@131500.4]
  wire  regs_465_io_enable; // @[RegFile.scala 66:20:@131500.4]
  wire  regs_466_clock; // @[RegFile.scala 66:20:@131514.4]
  wire  regs_466_reset; // @[RegFile.scala 66:20:@131514.4]
  wire [63:0] regs_466_io_in; // @[RegFile.scala 66:20:@131514.4]
  wire  regs_466_io_reset; // @[RegFile.scala 66:20:@131514.4]
  wire [63:0] regs_466_io_out; // @[RegFile.scala 66:20:@131514.4]
  wire  regs_466_io_enable; // @[RegFile.scala 66:20:@131514.4]
  wire  regs_467_clock; // @[RegFile.scala 66:20:@131528.4]
  wire  regs_467_reset; // @[RegFile.scala 66:20:@131528.4]
  wire [63:0] regs_467_io_in; // @[RegFile.scala 66:20:@131528.4]
  wire  regs_467_io_reset; // @[RegFile.scala 66:20:@131528.4]
  wire [63:0] regs_467_io_out; // @[RegFile.scala 66:20:@131528.4]
  wire  regs_467_io_enable; // @[RegFile.scala 66:20:@131528.4]
  wire  regs_468_clock; // @[RegFile.scala 66:20:@131542.4]
  wire  regs_468_reset; // @[RegFile.scala 66:20:@131542.4]
  wire [63:0] regs_468_io_in; // @[RegFile.scala 66:20:@131542.4]
  wire  regs_468_io_reset; // @[RegFile.scala 66:20:@131542.4]
  wire [63:0] regs_468_io_out; // @[RegFile.scala 66:20:@131542.4]
  wire  regs_468_io_enable; // @[RegFile.scala 66:20:@131542.4]
  wire  regs_469_clock; // @[RegFile.scala 66:20:@131556.4]
  wire  regs_469_reset; // @[RegFile.scala 66:20:@131556.4]
  wire [63:0] regs_469_io_in; // @[RegFile.scala 66:20:@131556.4]
  wire  regs_469_io_reset; // @[RegFile.scala 66:20:@131556.4]
  wire [63:0] regs_469_io_out; // @[RegFile.scala 66:20:@131556.4]
  wire  regs_469_io_enable; // @[RegFile.scala 66:20:@131556.4]
  wire  regs_470_clock; // @[RegFile.scala 66:20:@131570.4]
  wire  regs_470_reset; // @[RegFile.scala 66:20:@131570.4]
  wire [63:0] regs_470_io_in; // @[RegFile.scala 66:20:@131570.4]
  wire  regs_470_io_reset; // @[RegFile.scala 66:20:@131570.4]
  wire [63:0] regs_470_io_out; // @[RegFile.scala 66:20:@131570.4]
  wire  regs_470_io_enable; // @[RegFile.scala 66:20:@131570.4]
  wire  regs_471_clock; // @[RegFile.scala 66:20:@131584.4]
  wire  regs_471_reset; // @[RegFile.scala 66:20:@131584.4]
  wire [63:0] regs_471_io_in; // @[RegFile.scala 66:20:@131584.4]
  wire  regs_471_io_reset; // @[RegFile.scala 66:20:@131584.4]
  wire [63:0] regs_471_io_out; // @[RegFile.scala 66:20:@131584.4]
  wire  regs_471_io_enable; // @[RegFile.scala 66:20:@131584.4]
  wire  regs_472_clock; // @[RegFile.scala 66:20:@131598.4]
  wire  regs_472_reset; // @[RegFile.scala 66:20:@131598.4]
  wire [63:0] regs_472_io_in; // @[RegFile.scala 66:20:@131598.4]
  wire  regs_472_io_reset; // @[RegFile.scala 66:20:@131598.4]
  wire [63:0] regs_472_io_out; // @[RegFile.scala 66:20:@131598.4]
  wire  regs_472_io_enable; // @[RegFile.scala 66:20:@131598.4]
  wire  regs_473_clock; // @[RegFile.scala 66:20:@131612.4]
  wire  regs_473_reset; // @[RegFile.scala 66:20:@131612.4]
  wire [63:0] regs_473_io_in; // @[RegFile.scala 66:20:@131612.4]
  wire  regs_473_io_reset; // @[RegFile.scala 66:20:@131612.4]
  wire [63:0] regs_473_io_out; // @[RegFile.scala 66:20:@131612.4]
  wire  regs_473_io_enable; // @[RegFile.scala 66:20:@131612.4]
  wire  regs_474_clock; // @[RegFile.scala 66:20:@131626.4]
  wire  regs_474_reset; // @[RegFile.scala 66:20:@131626.4]
  wire [63:0] regs_474_io_in; // @[RegFile.scala 66:20:@131626.4]
  wire  regs_474_io_reset; // @[RegFile.scala 66:20:@131626.4]
  wire [63:0] regs_474_io_out; // @[RegFile.scala 66:20:@131626.4]
  wire  regs_474_io_enable; // @[RegFile.scala 66:20:@131626.4]
  wire  regs_475_clock; // @[RegFile.scala 66:20:@131640.4]
  wire  regs_475_reset; // @[RegFile.scala 66:20:@131640.4]
  wire [63:0] regs_475_io_in; // @[RegFile.scala 66:20:@131640.4]
  wire  regs_475_io_reset; // @[RegFile.scala 66:20:@131640.4]
  wire [63:0] regs_475_io_out; // @[RegFile.scala 66:20:@131640.4]
  wire  regs_475_io_enable; // @[RegFile.scala 66:20:@131640.4]
  wire  regs_476_clock; // @[RegFile.scala 66:20:@131654.4]
  wire  regs_476_reset; // @[RegFile.scala 66:20:@131654.4]
  wire [63:0] regs_476_io_in; // @[RegFile.scala 66:20:@131654.4]
  wire  regs_476_io_reset; // @[RegFile.scala 66:20:@131654.4]
  wire [63:0] regs_476_io_out; // @[RegFile.scala 66:20:@131654.4]
  wire  regs_476_io_enable; // @[RegFile.scala 66:20:@131654.4]
  wire  regs_477_clock; // @[RegFile.scala 66:20:@131668.4]
  wire  regs_477_reset; // @[RegFile.scala 66:20:@131668.4]
  wire [63:0] regs_477_io_in; // @[RegFile.scala 66:20:@131668.4]
  wire  regs_477_io_reset; // @[RegFile.scala 66:20:@131668.4]
  wire [63:0] regs_477_io_out; // @[RegFile.scala 66:20:@131668.4]
  wire  regs_477_io_enable; // @[RegFile.scala 66:20:@131668.4]
  wire  regs_478_clock; // @[RegFile.scala 66:20:@131682.4]
  wire  regs_478_reset; // @[RegFile.scala 66:20:@131682.4]
  wire [63:0] regs_478_io_in; // @[RegFile.scala 66:20:@131682.4]
  wire  regs_478_io_reset; // @[RegFile.scala 66:20:@131682.4]
  wire [63:0] regs_478_io_out; // @[RegFile.scala 66:20:@131682.4]
  wire  regs_478_io_enable; // @[RegFile.scala 66:20:@131682.4]
  wire  regs_479_clock; // @[RegFile.scala 66:20:@131696.4]
  wire  regs_479_reset; // @[RegFile.scala 66:20:@131696.4]
  wire [63:0] regs_479_io_in; // @[RegFile.scala 66:20:@131696.4]
  wire  regs_479_io_reset; // @[RegFile.scala 66:20:@131696.4]
  wire [63:0] regs_479_io_out; // @[RegFile.scala 66:20:@131696.4]
  wire  regs_479_io_enable; // @[RegFile.scala 66:20:@131696.4]
  wire  regs_480_clock; // @[RegFile.scala 66:20:@131710.4]
  wire  regs_480_reset; // @[RegFile.scala 66:20:@131710.4]
  wire [63:0] regs_480_io_in; // @[RegFile.scala 66:20:@131710.4]
  wire  regs_480_io_reset; // @[RegFile.scala 66:20:@131710.4]
  wire [63:0] regs_480_io_out; // @[RegFile.scala 66:20:@131710.4]
  wire  regs_480_io_enable; // @[RegFile.scala 66:20:@131710.4]
  wire  regs_481_clock; // @[RegFile.scala 66:20:@131724.4]
  wire  regs_481_reset; // @[RegFile.scala 66:20:@131724.4]
  wire [63:0] regs_481_io_in; // @[RegFile.scala 66:20:@131724.4]
  wire  regs_481_io_reset; // @[RegFile.scala 66:20:@131724.4]
  wire [63:0] regs_481_io_out; // @[RegFile.scala 66:20:@131724.4]
  wire  regs_481_io_enable; // @[RegFile.scala 66:20:@131724.4]
  wire  regs_482_clock; // @[RegFile.scala 66:20:@131738.4]
  wire  regs_482_reset; // @[RegFile.scala 66:20:@131738.4]
  wire [63:0] regs_482_io_in; // @[RegFile.scala 66:20:@131738.4]
  wire  regs_482_io_reset; // @[RegFile.scala 66:20:@131738.4]
  wire [63:0] regs_482_io_out; // @[RegFile.scala 66:20:@131738.4]
  wire  regs_482_io_enable; // @[RegFile.scala 66:20:@131738.4]
  wire  regs_483_clock; // @[RegFile.scala 66:20:@131752.4]
  wire  regs_483_reset; // @[RegFile.scala 66:20:@131752.4]
  wire [63:0] regs_483_io_in; // @[RegFile.scala 66:20:@131752.4]
  wire  regs_483_io_reset; // @[RegFile.scala 66:20:@131752.4]
  wire [63:0] regs_483_io_out; // @[RegFile.scala 66:20:@131752.4]
  wire  regs_483_io_enable; // @[RegFile.scala 66:20:@131752.4]
  wire  regs_484_clock; // @[RegFile.scala 66:20:@131766.4]
  wire  regs_484_reset; // @[RegFile.scala 66:20:@131766.4]
  wire [63:0] regs_484_io_in; // @[RegFile.scala 66:20:@131766.4]
  wire  regs_484_io_reset; // @[RegFile.scala 66:20:@131766.4]
  wire [63:0] regs_484_io_out; // @[RegFile.scala 66:20:@131766.4]
  wire  regs_484_io_enable; // @[RegFile.scala 66:20:@131766.4]
  wire  regs_485_clock; // @[RegFile.scala 66:20:@131780.4]
  wire  regs_485_reset; // @[RegFile.scala 66:20:@131780.4]
  wire [63:0] regs_485_io_in; // @[RegFile.scala 66:20:@131780.4]
  wire  regs_485_io_reset; // @[RegFile.scala 66:20:@131780.4]
  wire [63:0] regs_485_io_out; // @[RegFile.scala 66:20:@131780.4]
  wire  regs_485_io_enable; // @[RegFile.scala 66:20:@131780.4]
  wire  regs_486_clock; // @[RegFile.scala 66:20:@131794.4]
  wire  regs_486_reset; // @[RegFile.scala 66:20:@131794.4]
  wire [63:0] regs_486_io_in; // @[RegFile.scala 66:20:@131794.4]
  wire  regs_486_io_reset; // @[RegFile.scala 66:20:@131794.4]
  wire [63:0] regs_486_io_out; // @[RegFile.scala 66:20:@131794.4]
  wire  regs_486_io_enable; // @[RegFile.scala 66:20:@131794.4]
  wire  regs_487_clock; // @[RegFile.scala 66:20:@131808.4]
  wire  regs_487_reset; // @[RegFile.scala 66:20:@131808.4]
  wire [63:0] regs_487_io_in; // @[RegFile.scala 66:20:@131808.4]
  wire  regs_487_io_reset; // @[RegFile.scala 66:20:@131808.4]
  wire [63:0] regs_487_io_out; // @[RegFile.scala 66:20:@131808.4]
  wire  regs_487_io_enable; // @[RegFile.scala 66:20:@131808.4]
  wire  regs_488_clock; // @[RegFile.scala 66:20:@131822.4]
  wire  regs_488_reset; // @[RegFile.scala 66:20:@131822.4]
  wire [63:0] regs_488_io_in; // @[RegFile.scala 66:20:@131822.4]
  wire  regs_488_io_reset; // @[RegFile.scala 66:20:@131822.4]
  wire [63:0] regs_488_io_out; // @[RegFile.scala 66:20:@131822.4]
  wire  regs_488_io_enable; // @[RegFile.scala 66:20:@131822.4]
  wire  regs_489_clock; // @[RegFile.scala 66:20:@131836.4]
  wire  regs_489_reset; // @[RegFile.scala 66:20:@131836.4]
  wire [63:0] regs_489_io_in; // @[RegFile.scala 66:20:@131836.4]
  wire  regs_489_io_reset; // @[RegFile.scala 66:20:@131836.4]
  wire [63:0] regs_489_io_out; // @[RegFile.scala 66:20:@131836.4]
  wire  regs_489_io_enable; // @[RegFile.scala 66:20:@131836.4]
  wire  regs_490_clock; // @[RegFile.scala 66:20:@131850.4]
  wire  regs_490_reset; // @[RegFile.scala 66:20:@131850.4]
  wire [63:0] regs_490_io_in; // @[RegFile.scala 66:20:@131850.4]
  wire  regs_490_io_reset; // @[RegFile.scala 66:20:@131850.4]
  wire [63:0] regs_490_io_out; // @[RegFile.scala 66:20:@131850.4]
  wire  regs_490_io_enable; // @[RegFile.scala 66:20:@131850.4]
  wire  regs_491_clock; // @[RegFile.scala 66:20:@131864.4]
  wire  regs_491_reset; // @[RegFile.scala 66:20:@131864.4]
  wire [63:0] regs_491_io_in; // @[RegFile.scala 66:20:@131864.4]
  wire  regs_491_io_reset; // @[RegFile.scala 66:20:@131864.4]
  wire [63:0] regs_491_io_out; // @[RegFile.scala 66:20:@131864.4]
  wire  regs_491_io_enable; // @[RegFile.scala 66:20:@131864.4]
  wire  regs_492_clock; // @[RegFile.scala 66:20:@131878.4]
  wire  regs_492_reset; // @[RegFile.scala 66:20:@131878.4]
  wire [63:0] regs_492_io_in; // @[RegFile.scala 66:20:@131878.4]
  wire  regs_492_io_reset; // @[RegFile.scala 66:20:@131878.4]
  wire [63:0] regs_492_io_out; // @[RegFile.scala 66:20:@131878.4]
  wire  regs_492_io_enable; // @[RegFile.scala 66:20:@131878.4]
  wire  regs_493_clock; // @[RegFile.scala 66:20:@131892.4]
  wire  regs_493_reset; // @[RegFile.scala 66:20:@131892.4]
  wire [63:0] regs_493_io_in; // @[RegFile.scala 66:20:@131892.4]
  wire  regs_493_io_reset; // @[RegFile.scala 66:20:@131892.4]
  wire [63:0] regs_493_io_out; // @[RegFile.scala 66:20:@131892.4]
  wire  regs_493_io_enable; // @[RegFile.scala 66:20:@131892.4]
  wire  regs_494_clock; // @[RegFile.scala 66:20:@131906.4]
  wire  regs_494_reset; // @[RegFile.scala 66:20:@131906.4]
  wire [63:0] regs_494_io_in; // @[RegFile.scala 66:20:@131906.4]
  wire  regs_494_io_reset; // @[RegFile.scala 66:20:@131906.4]
  wire [63:0] regs_494_io_out; // @[RegFile.scala 66:20:@131906.4]
  wire  regs_494_io_enable; // @[RegFile.scala 66:20:@131906.4]
  wire  regs_495_clock; // @[RegFile.scala 66:20:@131920.4]
  wire  regs_495_reset; // @[RegFile.scala 66:20:@131920.4]
  wire [63:0] regs_495_io_in; // @[RegFile.scala 66:20:@131920.4]
  wire  regs_495_io_reset; // @[RegFile.scala 66:20:@131920.4]
  wire [63:0] regs_495_io_out; // @[RegFile.scala 66:20:@131920.4]
  wire  regs_495_io_enable; // @[RegFile.scala 66:20:@131920.4]
  wire  regs_496_clock; // @[RegFile.scala 66:20:@131934.4]
  wire  regs_496_reset; // @[RegFile.scala 66:20:@131934.4]
  wire [63:0] regs_496_io_in; // @[RegFile.scala 66:20:@131934.4]
  wire  regs_496_io_reset; // @[RegFile.scala 66:20:@131934.4]
  wire [63:0] regs_496_io_out; // @[RegFile.scala 66:20:@131934.4]
  wire  regs_496_io_enable; // @[RegFile.scala 66:20:@131934.4]
  wire  regs_497_clock; // @[RegFile.scala 66:20:@131948.4]
  wire  regs_497_reset; // @[RegFile.scala 66:20:@131948.4]
  wire [63:0] regs_497_io_in; // @[RegFile.scala 66:20:@131948.4]
  wire  regs_497_io_reset; // @[RegFile.scala 66:20:@131948.4]
  wire [63:0] regs_497_io_out; // @[RegFile.scala 66:20:@131948.4]
  wire  regs_497_io_enable; // @[RegFile.scala 66:20:@131948.4]
  wire  regs_498_clock; // @[RegFile.scala 66:20:@131962.4]
  wire  regs_498_reset; // @[RegFile.scala 66:20:@131962.4]
  wire [63:0] regs_498_io_in; // @[RegFile.scala 66:20:@131962.4]
  wire  regs_498_io_reset; // @[RegFile.scala 66:20:@131962.4]
  wire [63:0] regs_498_io_out; // @[RegFile.scala 66:20:@131962.4]
  wire  regs_498_io_enable; // @[RegFile.scala 66:20:@131962.4]
  wire  regs_499_clock; // @[RegFile.scala 66:20:@131976.4]
  wire  regs_499_reset; // @[RegFile.scala 66:20:@131976.4]
  wire [63:0] regs_499_io_in; // @[RegFile.scala 66:20:@131976.4]
  wire  regs_499_io_reset; // @[RegFile.scala 66:20:@131976.4]
  wire [63:0] regs_499_io_out; // @[RegFile.scala 66:20:@131976.4]
  wire  regs_499_io_enable; // @[RegFile.scala 66:20:@131976.4]
  wire  regs_500_clock; // @[RegFile.scala 66:20:@131990.4]
  wire  regs_500_reset; // @[RegFile.scala 66:20:@131990.4]
  wire [63:0] regs_500_io_in; // @[RegFile.scala 66:20:@131990.4]
  wire  regs_500_io_reset; // @[RegFile.scala 66:20:@131990.4]
  wire [63:0] regs_500_io_out; // @[RegFile.scala 66:20:@131990.4]
  wire  regs_500_io_enable; // @[RegFile.scala 66:20:@131990.4]
  wire  regs_501_clock; // @[RegFile.scala 66:20:@132004.4]
  wire  regs_501_reset; // @[RegFile.scala 66:20:@132004.4]
  wire [63:0] regs_501_io_in; // @[RegFile.scala 66:20:@132004.4]
  wire  regs_501_io_reset; // @[RegFile.scala 66:20:@132004.4]
  wire [63:0] regs_501_io_out; // @[RegFile.scala 66:20:@132004.4]
  wire  regs_501_io_enable; // @[RegFile.scala 66:20:@132004.4]
  wire  regs_502_clock; // @[RegFile.scala 66:20:@132018.4]
  wire  regs_502_reset; // @[RegFile.scala 66:20:@132018.4]
  wire [63:0] regs_502_io_in; // @[RegFile.scala 66:20:@132018.4]
  wire  regs_502_io_reset; // @[RegFile.scala 66:20:@132018.4]
  wire [63:0] regs_502_io_out; // @[RegFile.scala 66:20:@132018.4]
  wire  regs_502_io_enable; // @[RegFile.scala 66:20:@132018.4]
  wire [63:0] rport_io_ins_0; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_1; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_2; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_3; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_4; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_5; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_6; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_7; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_8; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_9; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_10; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_11; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_12; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_13; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_14; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_15; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_16; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_17; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_18; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_19; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_20; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_21; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_22; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_23; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_24; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_25; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_26; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_27; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_28; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_29; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_30; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_31; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_32; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_33; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_34; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_35; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_36; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_37; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_38; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_39; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_40; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_41; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_42; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_43; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_44; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_45; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_46; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_47; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_48; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_49; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_50; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_51; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_52; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_53; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_54; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_55; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_56; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_57; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_58; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_59; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_60; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_61; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_62; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_63; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_64; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_65; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_66; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_67; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_68; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_69; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_70; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_71; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_72; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_73; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_74; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_75; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_76; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_77; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_78; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_79; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_80; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_81; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_82; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_83; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_84; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_85; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_86; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_87; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_88; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_89; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_90; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_91; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_92; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_93; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_94; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_95; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_96; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_97; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_98; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_99; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_100; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_101; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_102; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_103; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_104; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_105; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_106; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_107; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_108; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_109; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_110; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_111; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_112; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_113; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_114; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_115; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_116; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_117; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_118; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_119; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_120; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_121; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_122; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_123; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_124; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_125; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_126; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_127; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_128; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_129; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_130; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_131; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_132; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_133; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_134; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_135; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_136; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_137; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_138; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_139; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_140; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_141; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_142; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_143; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_144; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_145; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_146; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_147; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_148; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_149; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_150; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_151; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_152; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_153; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_154; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_155; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_156; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_157; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_158; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_159; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_160; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_161; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_162; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_163; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_164; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_165; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_166; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_167; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_168; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_169; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_170; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_171; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_172; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_173; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_174; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_175; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_176; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_177; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_178; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_179; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_180; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_181; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_182; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_183; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_184; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_185; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_186; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_187; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_188; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_189; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_190; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_191; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_192; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_193; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_194; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_195; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_196; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_197; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_198; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_199; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_200; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_201; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_202; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_203; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_204; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_205; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_206; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_207; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_208; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_209; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_210; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_211; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_212; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_213; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_214; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_215; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_216; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_217; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_218; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_219; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_220; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_221; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_222; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_223; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_224; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_225; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_226; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_227; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_228; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_229; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_230; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_231; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_232; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_233; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_234; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_235; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_236; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_237; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_238; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_239; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_240; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_241; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_242; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_243; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_244; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_245; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_246; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_247; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_248; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_249; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_250; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_251; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_252; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_253; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_254; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_255; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_256; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_257; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_258; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_259; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_260; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_261; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_262; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_263; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_264; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_265; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_266; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_267; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_268; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_269; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_270; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_271; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_272; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_273; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_274; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_275; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_276; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_277; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_278; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_279; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_280; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_281; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_282; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_283; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_284; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_285; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_286; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_287; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_288; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_289; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_290; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_291; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_292; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_293; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_294; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_295; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_296; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_297; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_298; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_299; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_300; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_301; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_302; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_303; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_304; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_305; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_306; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_307; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_308; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_309; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_310; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_311; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_312; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_313; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_314; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_315; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_316; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_317; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_318; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_319; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_320; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_321; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_322; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_323; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_324; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_325; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_326; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_327; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_328; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_329; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_330; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_331; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_332; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_333; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_334; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_335; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_336; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_337; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_338; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_339; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_340; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_341; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_342; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_343; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_344; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_345; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_346; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_347; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_348; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_349; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_350; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_351; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_352; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_353; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_354; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_355; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_356; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_357; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_358; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_359; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_360; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_361; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_362; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_363; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_364; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_365; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_366; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_367; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_368; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_369; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_370; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_371; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_372; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_373; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_374; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_375; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_376; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_377; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_378; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_379; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_380; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_381; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_382; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_383; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_384; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_385; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_386; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_387; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_388; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_389; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_390; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_391; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_392; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_393; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_394; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_395; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_396; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_397; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_398; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_399; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_400; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_401; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_402; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_403; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_404; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_405; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_406; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_407; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_408; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_409; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_410; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_411; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_412; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_413; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_414; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_415; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_416; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_417; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_418; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_419; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_420; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_421; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_422; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_423; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_424; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_425; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_426; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_427; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_428; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_429; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_430; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_431; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_432; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_433; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_434; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_435; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_436; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_437; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_438; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_439; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_440; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_441; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_442; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_443; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_444; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_445; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_446; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_447; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_448; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_449; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_450; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_451; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_452; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_453; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_454; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_455; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_456; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_457; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_458; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_459; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_460; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_461; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_462; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_463; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_464; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_465; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_466; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_467; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_468; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_469; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_470; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_471; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_472; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_473; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_474; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_475; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_476; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_477; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_478; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_479; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_480; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_481; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_482; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_483; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_484; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_485; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_486; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_487; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_488; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_489; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_490; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_491; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_492; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_493; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_494; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_495; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_496; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_497; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_498; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_499; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_500; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_501; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_ins_502; // @[RegFile.scala 95:21:@132032.4]
  wire [8:0] rport_io_sel; // @[RegFile.scala 95:21:@132032.4]
  wire [63:0] rport_io_out; // @[RegFile.scala 95:21:@132032.4]
  wire  _T_3078; // @[RegFile.scala 80:42:@124994.4]
  wire  _T_3084; // @[RegFile.scala 68:46:@125006.4]
  wire  _T_3085; // @[RegFile.scala 68:34:@125007.4]
  wire  _T_3098; // @[RegFile.scala 80:42:@125025.4]
  wire  _T_3104; // @[RegFile.scala 80:42:@125037.4]
  wire  _T_3110; // @[RegFile.scala 74:80:@125049.4]
  wire  _T_3111; // @[RegFile.scala 74:68:@125050.4]
  FringeFF regs_0 ( // @[RegFile.scala 66:20:@124991.4]
    .clock(regs_0_clock),
    .reset(regs_0_reset),
    .io_in(regs_0_io_in),
    .io_reset(regs_0_io_reset),
    .io_out(regs_0_io_out),
    .io_enable(regs_0_io_enable)
  );
  FringeFF regs_1 ( // @[RegFile.scala 66:20:@125003.4]
    .clock(regs_1_clock),
    .reset(regs_1_reset),
    .io_in(regs_1_io_in),
    .io_reset(regs_1_io_reset),
    .io_out(regs_1_io_out),
    .io_enable(regs_1_io_enable)
  );
  FringeFF regs_2 ( // @[RegFile.scala 66:20:@125022.4]
    .clock(regs_2_clock),
    .reset(regs_2_reset),
    .io_in(regs_2_io_in),
    .io_reset(regs_2_io_reset),
    .io_out(regs_2_io_out),
    .io_enable(regs_2_io_enable)
  );
  FringeFF regs_3 ( // @[RegFile.scala 66:20:@125034.4]
    .clock(regs_3_clock),
    .reset(regs_3_reset),
    .io_in(regs_3_io_in),
    .io_reset(regs_3_io_reset),
    .io_out(regs_3_io_out),
    .io_enable(regs_3_io_enable)
  );
  FringeFF regs_4 ( // @[RegFile.scala 66:20:@125046.4]
    .clock(regs_4_clock),
    .reset(regs_4_reset),
    .io_in(regs_4_io_in),
    .io_reset(regs_4_io_reset),
    .io_out(regs_4_io_out),
    .io_enable(regs_4_io_enable)
  );
  FringeFF regs_5 ( // @[RegFile.scala 66:20:@125060.4]
    .clock(regs_5_clock),
    .reset(regs_5_reset),
    .io_in(regs_5_io_in),
    .io_reset(regs_5_io_reset),
    .io_out(regs_5_io_out),
    .io_enable(regs_5_io_enable)
  );
  FringeFF regs_6 ( // @[RegFile.scala 66:20:@125074.4]
    .clock(regs_6_clock),
    .reset(regs_6_reset),
    .io_in(regs_6_io_in),
    .io_reset(regs_6_io_reset),
    .io_out(regs_6_io_out),
    .io_enable(regs_6_io_enable)
  );
  FringeFF regs_7 ( // @[RegFile.scala 66:20:@125088.4]
    .clock(regs_7_clock),
    .reset(regs_7_reset),
    .io_in(regs_7_io_in),
    .io_reset(regs_7_io_reset),
    .io_out(regs_7_io_out),
    .io_enable(regs_7_io_enable)
  );
  FringeFF regs_8 ( // @[RegFile.scala 66:20:@125102.4]
    .clock(regs_8_clock),
    .reset(regs_8_reset),
    .io_in(regs_8_io_in),
    .io_reset(regs_8_io_reset),
    .io_out(regs_8_io_out),
    .io_enable(regs_8_io_enable)
  );
  FringeFF regs_9 ( // @[RegFile.scala 66:20:@125116.4]
    .clock(regs_9_clock),
    .reset(regs_9_reset),
    .io_in(regs_9_io_in),
    .io_reset(regs_9_io_reset),
    .io_out(regs_9_io_out),
    .io_enable(regs_9_io_enable)
  );
  FringeFF regs_10 ( // @[RegFile.scala 66:20:@125130.4]
    .clock(regs_10_clock),
    .reset(regs_10_reset),
    .io_in(regs_10_io_in),
    .io_reset(regs_10_io_reset),
    .io_out(regs_10_io_out),
    .io_enable(regs_10_io_enable)
  );
  FringeFF regs_11 ( // @[RegFile.scala 66:20:@125144.4]
    .clock(regs_11_clock),
    .reset(regs_11_reset),
    .io_in(regs_11_io_in),
    .io_reset(regs_11_io_reset),
    .io_out(regs_11_io_out),
    .io_enable(regs_11_io_enable)
  );
  FringeFF regs_12 ( // @[RegFile.scala 66:20:@125158.4]
    .clock(regs_12_clock),
    .reset(regs_12_reset),
    .io_in(regs_12_io_in),
    .io_reset(regs_12_io_reset),
    .io_out(regs_12_io_out),
    .io_enable(regs_12_io_enable)
  );
  FringeFF regs_13 ( // @[RegFile.scala 66:20:@125172.4]
    .clock(regs_13_clock),
    .reset(regs_13_reset),
    .io_in(regs_13_io_in),
    .io_reset(regs_13_io_reset),
    .io_out(regs_13_io_out),
    .io_enable(regs_13_io_enable)
  );
  FringeFF regs_14 ( // @[RegFile.scala 66:20:@125186.4]
    .clock(regs_14_clock),
    .reset(regs_14_reset),
    .io_in(regs_14_io_in),
    .io_reset(regs_14_io_reset),
    .io_out(regs_14_io_out),
    .io_enable(regs_14_io_enable)
  );
  FringeFF regs_15 ( // @[RegFile.scala 66:20:@125200.4]
    .clock(regs_15_clock),
    .reset(regs_15_reset),
    .io_in(regs_15_io_in),
    .io_reset(regs_15_io_reset),
    .io_out(regs_15_io_out),
    .io_enable(regs_15_io_enable)
  );
  FringeFF regs_16 ( // @[RegFile.scala 66:20:@125214.4]
    .clock(regs_16_clock),
    .reset(regs_16_reset),
    .io_in(regs_16_io_in),
    .io_reset(regs_16_io_reset),
    .io_out(regs_16_io_out),
    .io_enable(regs_16_io_enable)
  );
  FringeFF regs_17 ( // @[RegFile.scala 66:20:@125228.4]
    .clock(regs_17_clock),
    .reset(regs_17_reset),
    .io_in(regs_17_io_in),
    .io_reset(regs_17_io_reset),
    .io_out(regs_17_io_out),
    .io_enable(regs_17_io_enable)
  );
  FringeFF regs_18 ( // @[RegFile.scala 66:20:@125242.4]
    .clock(regs_18_clock),
    .reset(regs_18_reset),
    .io_in(regs_18_io_in),
    .io_reset(regs_18_io_reset),
    .io_out(regs_18_io_out),
    .io_enable(regs_18_io_enable)
  );
  FringeFF regs_19 ( // @[RegFile.scala 66:20:@125256.4]
    .clock(regs_19_clock),
    .reset(regs_19_reset),
    .io_in(regs_19_io_in),
    .io_reset(regs_19_io_reset),
    .io_out(regs_19_io_out),
    .io_enable(regs_19_io_enable)
  );
  FringeFF regs_20 ( // @[RegFile.scala 66:20:@125270.4]
    .clock(regs_20_clock),
    .reset(regs_20_reset),
    .io_in(regs_20_io_in),
    .io_reset(regs_20_io_reset),
    .io_out(regs_20_io_out),
    .io_enable(regs_20_io_enable)
  );
  FringeFF regs_21 ( // @[RegFile.scala 66:20:@125284.4]
    .clock(regs_21_clock),
    .reset(regs_21_reset),
    .io_in(regs_21_io_in),
    .io_reset(regs_21_io_reset),
    .io_out(regs_21_io_out),
    .io_enable(regs_21_io_enable)
  );
  FringeFF regs_22 ( // @[RegFile.scala 66:20:@125298.4]
    .clock(regs_22_clock),
    .reset(regs_22_reset),
    .io_in(regs_22_io_in),
    .io_reset(regs_22_io_reset),
    .io_out(regs_22_io_out),
    .io_enable(regs_22_io_enable)
  );
  FringeFF regs_23 ( // @[RegFile.scala 66:20:@125312.4]
    .clock(regs_23_clock),
    .reset(regs_23_reset),
    .io_in(regs_23_io_in),
    .io_reset(regs_23_io_reset),
    .io_out(regs_23_io_out),
    .io_enable(regs_23_io_enable)
  );
  FringeFF regs_24 ( // @[RegFile.scala 66:20:@125326.4]
    .clock(regs_24_clock),
    .reset(regs_24_reset),
    .io_in(regs_24_io_in),
    .io_reset(regs_24_io_reset),
    .io_out(regs_24_io_out),
    .io_enable(regs_24_io_enable)
  );
  FringeFF regs_25 ( // @[RegFile.scala 66:20:@125340.4]
    .clock(regs_25_clock),
    .reset(regs_25_reset),
    .io_in(regs_25_io_in),
    .io_reset(regs_25_io_reset),
    .io_out(regs_25_io_out),
    .io_enable(regs_25_io_enable)
  );
  FringeFF regs_26 ( // @[RegFile.scala 66:20:@125354.4]
    .clock(regs_26_clock),
    .reset(regs_26_reset),
    .io_in(regs_26_io_in),
    .io_reset(regs_26_io_reset),
    .io_out(regs_26_io_out),
    .io_enable(regs_26_io_enable)
  );
  FringeFF regs_27 ( // @[RegFile.scala 66:20:@125368.4]
    .clock(regs_27_clock),
    .reset(regs_27_reset),
    .io_in(regs_27_io_in),
    .io_reset(regs_27_io_reset),
    .io_out(regs_27_io_out),
    .io_enable(regs_27_io_enable)
  );
  FringeFF regs_28 ( // @[RegFile.scala 66:20:@125382.4]
    .clock(regs_28_clock),
    .reset(regs_28_reset),
    .io_in(regs_28_io_in),
    .io_reset(regs_28_io_reset),
    .io_out(regs_28_io_out),
    .io_enable(regs_28_io_enable)
  );
  FringeFF regs_29 ( // @[RegFile.scala 66:20:@125396.4]
    .clock(regs_29_clock),
    .reset(regs_29_reset),
    .io_in(regs_29_io_in),
    .io_reset(regs_29_io_reset),
    .io_out(regs_29_io_out),
    .io_enable(regs_29_io_enable)
  );
  FringeFF regs_30 ( // @[RegFile.scala 66:20:@125410.4]
    .clock(regs_30_clock),
    .reset(regs_30_reset),
    .io_in(regs_30_io_in),
    .io_reset(regs_30_io_reset),
    .io_out(regs_30_io_out),
    .io_enable(regs_30_io_enable)
  );
  FringeFF regs_31 ( // @[RegFile.scala 66:20:@125424.4]
    .clock(regs_31_clock),
    .reset(regs_31_reset),
    .io_in(regs_31_io_in),
    .io_reset(regs_31_io_reset),
    .io_out(regs_31_io_out),
    .io_enable(regs_31_io_enable)
  );
  FringeFF regs_32 ( // @[RegFile.scala 66:20:@125438.4]
    .clock(regs_32_clock),
    .reset(regs_32_reset),
    .io_in(regs_32_io_in),
    .io_reset(regs_32_io_reset),
    .io_out(regs_32_io_out),
    .io_enable(regs_32_io_enable)
  );
  FringeFF regs_33 ( // @[RegFile.scala 66:20:@125452.4]
    .clock(regs_33_clock),
    .reset(regs_33_reset),
    .io_in(regs_33_io_in),
    .io_reset(regs_33_io_reset),
    .io_out(regs_33_io_out),
    .io_enable(regs_33_io_enable)
  );
  FringeFF regs_34 ( // @[RegFile.scala 66:20:@125466.4]
    .clock(regs_34_clock),
    .reset(regs_34_reset),
    .io_in(regs_34_io_in),
    .io_reset(regs_34_io_reset),
    .io_out(regs_34_io_out),
    .io_enable(regs_34_io_enable)
  );
  FringeFF regs_35 ( // @[RegFile.scala 66:20:@125480.4]
    .clock(regs_35_clock),
    .reset(regs_35_reset),
    .io_in(regs_35_io_in),
    .io_reset(regs_35_io_reset),
    .io_out(regs_35_io_out),
    .io_enable(regs_35_io_enable)
  );
  FringeFF regs_36 ( // @[RegFile.scala 66:20:@125494.4]
    .clock(regs_36_clock),
    .reset(regs_36_reset),
    .io_in(regs_36_io_in),
    .io_reset(regs_36_io_reset),
    .io_out(regs_36_io_out),
    .io_enable(regs_36_io_enable)
  );
  FringeFF regs_37 ( // @[RegFile.scala 66:20:@125508.4]
    .clock(regs_37_clock),
    .reset(regs_37_reset),
    .io_in(regs_37_io_in),
    .io_reset(regs_37_io_reset),
    .io_out(regs_37_io_out),
    .io_enable(regs_37_io_enable)
  );
  FringeFF regs_38 ( // @[RegFile.scala 66:20:@125522.4]
    .clock(regs_38_clock),
    .reset(regs_38_reset),
    .io_in(regs_38_io_in),
    .io_reset(regs_38_io_reset),
    .io_out(regs_38_io_out),
    .io_enable(regs_38_io_enable)
  );
  FringeFF regs_39 ( // @[RegFile.scala 66:20:@125536.4]
    .clock(regs_39_clock),
    .reset(regs_39_reset),
    .io_in(regs_39_io_in),
    .io_reset(regs_39_io_reset),
    .io_out(regs_39_io_out),
    .io_enable(regs_39_io_enable)
  );
  FringeFF regs_40 ( // @[RegFile.scala 66:20:@125550.4]
    .clock(regs_40_clock),
    .reset(regs_40_reset),
    .io_in(regs_40_io_in),
    .io_reset(regs_40_io_reset),
    .io_out(regs_40_io_out),
    .io_enable(regs_40_io_enable)
  );
  FringeFF regs_41 ( // @[RegFile.scala 66:20:@125564.4]
    .clock(regs_41_clock),
    .reset(regs_41_reset),
    .io_in(regs_41_io_in),
    .io_reset(regs_41_io_reset),
    .io_out(regs_41_io_out),
    .io_enable(regs_41_io_enable)
  );
  FringeFF regs_42 ( // @[RegFile.scala 66:20:@125578.4]
    .clock(regs_42_clock),
    .reset(regs_42_reset),
    .io_in(regs_42_io_in),
    .io_reset(regs_42_io_reset),
    .io_out(regs_42_io_out),
    .io_enable(regs_42_io_enable)
  );
  FringeFF regs_43 ( // @[RegFile.scala 66:20:@125592.4]
    .clock(regs_43_clock),
    .reset(regs_43_reset),
    .io_in(regs_43_io_in),
    .io_reset(regs_43_io_reset),
    .io_out(regs_43_io_out),
    .io_enable(regs_43_io_enable)
  );
  FringeFF regs_44 ( // @[RegFile.scala 66:20:@125606.4]
    .clock(regs_44_clock),
    .reset(regs_44_reset),
    .io_in(regs_44_io_in),
    .io_reset(regs_44_io_reset),
    .io_out(regs_44_io_out),
    .io_enable(regs_44_io_enable)
  );
  FringeFF regs_45 ( // @[RegFile.scala 66:20:@125620.4]
    .clock(regs_45_clock),
    .reset(regs_45_reset),
    .io_in(regs_45_io_in),
    .io_reset(regs_45_io_reset),
    .io_out(regs_45_io_out),
    .io_enable(regs_45_io_enable)
  );
  FringeFF regs_46 ( // @[RegFile.scala 66:20:@125634.4]
    .clock(regs_46_clock),
    .reset(regs_46_reset),
    .io_in(regs_46_io_in),
    .io_reset(regs_46_io_reset),
    .io_out(regs_46_io_out),
    .io_enable(regs_46_io_enable)
  );
  FringeFF regs_47 ( // @[RegFile.scala 66:20:@125648.4]
    .clock(regs_47_clock),
    .reset(regs_47_reset),
    .io_in(regs_47_io_in),
    .io_reset(regs_47_io_reset),
    .io_out(regs_47_io_out),
    .io_enable(regs_47_io_enable)
  );
  FringeFF regs_48 ( // @[RegFile.scala 66:20:@125662.4]
    .clock(regs_48_clock),
    .reset(regs_48_reset),
    .io_in(regs_48_io_in),
    .io_reset(regs_48_io_reset),
    .io_out(regs_48_io_out),
    .io_enable(regs_48_io_enable)
  );
  FringeFF regs_49 ( // @[RegFile.scala 66:20:@125676.4]
    .clock(regs_49_clock),
    .reset(regs_49_reset),
    .io_in(regs_49_io_in),
    .io_reset(regs_49_io_reset),
    .io_out(regs_49_io_out),
    .io_enable(regs_49_io_enable)
  );
  FringeFF regs_50 ( // @[RegFile.scala 66:20:@125690.4]
    .clock(regs_50_clock),
    .reset(regs_50_reset),
    .io_in(regs_50_io_in),
    .io_reset(regs_50_io_reset),
    .io_out(regs_50_io_out),
    .io_enable(regs_50_io_enable)
  );
  FringeFF regs_51 ( // @[RegFile.scala 66:20:@125704.4]
    .clock(regs_51_clock),
    .reset(regs_51_reset),
    .io_in(regs_51_io_in),
    .io_reset(regs_51_io_reset),
    .io_out(regs_51_io_out),
    .io_enable(regs_51_io_enable)
  );
  FringeFF regs_52 ( // @[RegFile.scala 66:20:@125718.4]
    .clock(regs_52_clock),
    .reset(regs_52_reset),
    .io_in(regs_52_io_in),
    .io_reset(regs_52_io_reset),
    .io_out(regs_52_io_out),
    .io_enable(regs_52_io_enable)
  );
  FringeFF regs_53 ( // @[RegFile.scala 66:20:@125732.4]
    .clock(regs_53_clock),
    .reset(regs_53_reset),
    .io_in(regs_53_io_in),
    .io_reset(regs_53_io_reset),
    .io_out(regs_53_io_out),
    .io_enable(regs_53_io_enable)
  );
  FringeFF regs_54 ( // @[RegFile.scala 66:20:@125746.4]
    .clock(regs_54_clock),
    .reset(regs_54_reset),
    .io_in(regs_54_io_in),
    .io_reset(regs_54_io_reset),
    .io_out(regs_54_io_out),
    .io_enable(regs_54_io_enable)
  );
  FringeFF regs_55 ( // @[RegFile.scala 66:20:@125760.4]
    .clock(regs_55_clock),
    .reset(regs_55_reset),
    .io_in(regs_55_io_in),
    .io_reset(regs_55_io_reset),
    .io_out(regs_55_io_out),
    .io_enable(regs_55_io_enable)
  );
  FringeFF regs_56 ( // @[RegFile.scala 66:20:@125774.4]
    .clock(regs_56_clock),
    .reset(regs_56_reset),
    .io_in(regs_56_io_in),
    .io_reset(regs_56_io_reset),
    .io_out(regs_56_io_out),
    .io_enable(regs_56_io_enable)
  );
  FringeFF regs_57 ( // @[RegFile.scala 66:20:@125788.4]
    .clock(regs_57_clock),
    .reset(regs_57_reset),
    .io_in(regs_57_io_in),
    .io_reset(regs_57_io_reset),
    .io_out(regs_57_io_out),
    .io_enable(regs_57_io_enable)
  );
  FringeFF regs_58 ( // @[RegFile.scala 66:20:@125802.4]
    .clock(regs_58_clock),
    .reset(regs_58_reset),
    .io_in(regs_58_io_in),
    .io_reset(regs_58_io_reset),
    .io_out(regs_58_io_out),
    .io_enable(regs_58_io_enable)
  );
  FringeFF regs_59 ( // @[RegFile.scala 66:20:@125816.4]
    .clock(regs_59_clock),
    .reset(regs_59_reset),
    .io_in(regs_59_io_in),
    .io_reset(regs_59_io_reset),
    .io_out(regs_59_io_out),
    .io_enable(regs_59_io_enable)
  );
  FringeFF regs_60 ( // @[RegFile.scala 66:20:@125830.4]
    .clock(regs_60_clock),
    .reset(regs_60_reset),
    .io_in(regs_60_io_in),
    .io_reset(regs_60_io_reset),
    .io_out(regs_60_io_out),
    .io_enable(regs_60_io_enable)
  );
  FringeFF regs_61 ( // @[RegFile.scala 66:20:@125844.4]
    .clock(regs_61_clock),
    .reset(regs_61_reset),
    .io_in(regs_61_io_in),
    .io_reset(regs_61_io_reset),
    .io_out(regs_61_io_out),
    .io_enable(regs_61_io_enable)
  );
  FringeFF regs_62 ( // @[RegFile.scala 66:20:@125858.4]
    .clock(regs_62_clock),
    .reset(regs_62_reset),
    .io_in(regs_62_io_in),
    .io_reset(regs_62_io_reset),
    .io_out(regs_62_io_out),
    .io_enable(regs_62_io_enable)
  );
  FringeFF regs_63 ( // @[RegFile.scala 66:20:@125872.4]
    .clock(regs_63_clock),
    .reset(regs_63_reset),
    .io_in(regs_63_io_in),
    .io_reset(regs_63_io_reset),
    .io_out(regs_63_io_out),
    .io_enable(regs_63_io_enable)
  );
  FringeFF regs_64 ( // @[RegFile.scala 66:20:@125886.4]
    .clock(regs_64_clock),
    .reset(regs_64_reset),
    .io_in(regs_64_io_in),
    .io_reset(regs_64_io_reset),
    .io_out(regs_64_io_out),
    .io_enable(regs_64_io_enable)
  );
  FringeFF regs_65 ( // @[RegFile.scala 66:20:@125900.4]
    .clock(regs_65_clock),
    .reset(regs_65_reset),
    .io_in(regs_65_io_in),
    .io_reset(regs_65_io_reset),
    .io_out(regs_65_io_out),
    .io_enable(regs_65_io_enable)
  );
  FringeFF regs_66 ( // @[RegFile.scala 66:20:@125914.4]
    .clock(regs_66_clock),
    .reset(regs_66_reset),
    .io_in(regs_66_io_in),
    .io_reset(regs_66_io_reset),
    .io_out(regs_66_io_out),
    .io_enable(regs_66_io_enable)
  );
  FringeFF regs_67 ( // @[RegFile.scala 66:20:@125928.4]
    .clock(regs_67_clock),
    .reset(regs_67_reset),
    .io_in(regs_67_io_in),
    .io_reset(regs_67_io_reset),
    .io_out(regs_67_io_out),
    .io_enable(regs_67_io_enable)
  );
  FringeFF regs_68 ( // @[RegFile.scala 66:20:@125942.4]
    .clock(regs_68_clock),
    .reset(regs_68_reset),
    .io_in(regs_68_io_in),
    .io_reset(regs_68_io_reset),
    .io_out(regs_68_io_out),
    .io_enable(regs_68_io_enable)
  );
  FringeFF regs_69 ( // @[RegFile.scala 66:20:@125956.4]
    .clock(regs_69_clock),
    .reset(regs_69_reset),
    .io_in(regs_69_io_in),
    .io_reset(regs_69_io_reset),
    .io_out(regs_69_io_out),
    .io_enable(regs_69_io_enable)
  );
  FringeFF regs_70 ( // @[RegFile.scala 66:20:@125970.4]
    .clock(regs_70_clock),
    .reset(regs_70_reset),
    .io_in(regs_70_io_in),
    .io_reset(regs_70_io_reset),
    .io_out(regs_70_io_out),
    .io_enable(regs_70_io_enable)
  );
  FringeFF regs_71 ( // @[RegFile.scala 66:20:@125984.4]
    .clock(regs_71_clock),
    .reset(regs_71_reset),
    .io_in(regs_71_io_in),
    .io_reset(regs_71_io_reset),
    .io_out(regs_71_io_out),
    .io_enable(regs_71_io_enable)
  );
  FringeFF regs_72 ( // @[RegFile.scala 66:20:@125998.4]
    .clock(regs_72_clock),
    .reset(regs_72_reset),
    .io_in(regs_72_io_in),
    .io_reset(regs_72_io_reset),
    .io_out(regs_72_io_out),
    .io_enable(regs_72_io_enable)
  );
  FringeFF regs_73 ( // @[RegFile.scala 66:20:@126012.4]
    .clock(regs_73_clock),
    .reset(regs_73_reset),
    .io_in(regs_73_io_in),
    .io_reset(regs_73_io_reset),
    .io_out(regs_73_io_out),
    .io_enable(regs_73_io_enable)
  );
  FringeFF regs_74 ( // @[RegFile.scala 66:20:@126026.4]
    .clock(regs_74_clock),
    .reset(regs_74_reset),
    .io_in(regs_74_io_in),
    .io_reset(regs_74_io_reset),
    .io_out(regs_74_io_out),
    .io_enable(regs_74_io_enable)
  );
  FringeFF regs_75 ( // @[RegFile.scala 66:20:@126040.4]
    .clock(regs_75_clock),
    .reset(regs_75_reset),
    .io_in(regs_75_io_in),
    .io_reset(regs_75_io_reset),
    .io_out(regs_75_io_out),
    .io_enable(regs_75_io_enable)
  );
  FringeFF regs_76 ( // @[RegFile.scala 66:20:@126054.4]
    .clock(regs_76_clock),
    .reset(regs_76_reset),
    .io_in(regs_76_io_in),
    .io_reset(regs_76_io_reset),
    .io_out(regs_76_io_out),
    .io_enable(regs_76_io_enable)
  );
  FringeFF regs_77 ( // @[RegFile.scala 66:20:@126068.4]
    .clock(regs_77_clock),
    .reset(regs_77_reset),
    .io_in(regs_77_io_in),
    .io_reset(regs_77_io_reset),
    .io_out(regs_77_io_out),
    .io_enable(regs_77_io_enable)
  );
  FringeFF regs_78 ( // @[RegFile.scala 66:20:@126082.4]
    .clock(regs_78_clock),
    .reset(regs_78_reset),
    .io_in(regs_78_io_in),
    .io_reset(regs_78_io_reset),
    .io_out(regs_78_io_out),
    .io_enable(regs_78_io_enable)
  );
  FringeFF regs_79 ( // @[RegFile.scala 66:20:@126096.4]
    .clock(regs_79_clock),
    .reset(regs_79_reset),
    .io_in(regs_79_io_in),
    .io_reset(regs_79_io_reset),
    .io_out(regs_79_io_out),
    .io_enable(regs_79_io_enable)
  );
  FringeFF regs_80 ( // @[RegFile.scala 66:20:@126110.4]
    .clock(regs_80_clock),
    .reset(regs_80_reset),
    .io_in(regs_80_io_in),
    .io_reset(regs_80_io_reset),
    .io_out(regs_80_io_out),
    .io_enable(regs_80_io_enable)
  );
  FringeFF regs_81 ( // @[RegFile.scala 66:20:@126124.4]
    .clock(regs_81_clock),
    .reset(regs_81_reset),
    .io_in(regs_81_io_in),
    .io_reset(regs_81_io_reset),
    .io_out(regs_81_io_out),
    .io_enable(regs_81_io_enable)
  );
  FringeFF regs_82 ( // @[RegFile.scala 66:20:@126138.4]
    .clock(regs_82_clock),
    .reset(regs_82_reset),
    .io_in(regs_82_io_in),
    .io_reset(regs_82_io_reset),
    .io_out(regs_82_io_out),
    .io_enable(regs_82_io_enable)
  );
  FringeFF regs_83 ( // @[RegFile.scala 66:20:@126152.4]
    .clock(regs_83_clock),
    .reset(regs_83_reset),
    .io_in(regs_83_io_in),
    .io_reset(regs_83_io_reset),
    .io_out(regs_83_io_out),
    .io_enable(regs_83_io_enable)
  );
  FringeFF regs_84 ( // @[RegFile.scala 66:20:@126166.4]
    .clock(regs_84_clock),
    .reset(regs_84_reset),
    .io_in(regs_84_io_in),
    .io_reset(regs_84_io_reset),
    .io_out(regs_84_io_out),
    .io_enable(regs_84_io_enable)
  );
  FringeFF regs_85 ( // @[RegFile.scala 66:20:@126180.4]
    .clock(regs_85_clock),
    .reset(regs_85_reset),
    .io_in(regs_85_io_in),
    .io_reset(regs_85_io_reset),
    .io_out(regs_85_io_out),
    .io_enable(regs_85_io_enable)
  );
  FringeFF regs_86 ( // @[RegFile.scala 66:20:@126194.4]
    .clock(regs_86_clock),
    .reset(regs_86_reset),
    .io_in(regs_86_io_in),
    .io_reset(regs_86_io_reset),
    .io_out(regs_86_io_out),
    .io_enable(regs_86_io_enable)
  );
  FringeFF regs_87 ( // @[RegFile.scala 66:20:@126208.4]
    .clock(regs_87_clock),
    .reset(regs_87_reset),
    .io_in(regs_87_io_in),
    .io_reset(regs_87_io_reset),
    .io_out(regs_87_io_out),
    .io_enable(regs_87_io_enable)
  );
  FringeFF regs_88 ( // @[RegFile.scala 66:20:@126222.4]
    .clock(regs_88_clock),
    .reset(regs_88_reset),
    .io_in(regs_88_io_in),
    .io_reset(regs_88_io_reset),
    .io_out(regs_88_io_out),
    .io_enable(regs_88_io_enable)
  );
  FringeFF regs_89 ( // @[RegFile.scala 66:20:@126236.4]
    .clock(regs_89_clock),
    .reset(regs_89_reset),
    .io_in(regs_89_io_in),
    .io_reset(regs_89_io_reset),
    .io_out(regs_89_io_out),
    .io_enable(regs_89_io_enable)
  );
  FringeFF regs_90 ( // @[RegFile.scala 66:20:@126250.4]
    .clock(regs_90_clock),
    .reset(regs_90_reset),
    .io_in(regs_90_io_in),
    .io_reset(regs_90_io_reset),
    .io_out(regs_90_io_out),
    .io_enable(regs_90_io_enable)
  );
  FringeFF regs_91 ( // @[RegFile.scala 66:20:@126264.4]
    .clock(regs_91_clock),
    .reset(regs_91_reset),
    .io_in(regs_91_io_in),
    .io_reset(regs_91_io_reset),
    .io_out(regs_91_io_out),
    .io_enable(regs_91_io_enable)
  );
  FringeFF regs_92 ( // @[RegFile.scala 66:20:@126278.4]
    .clock(regs_92_clock),
    .reset(regs_92_reset),
    .io_in(regs_92_io_in),
    .io_reset(regs_92_io_reset),
    .io_out(regs_92_io_out),
    .io_enable(regs_92_io_enable)
  );
  FringeFF regs_93 ( // @[RegFile.scala 66:20:@126292.4]
    .clock(regs_93_clock),
    .reset(regs_93_reset),
    .io_in(regs_93_io_in),
    .io_reset(regs_93_io_reset),
    .io_out(regs_93_io_out),
    .io_enable(regs_93_io_enable)
  );
  FringeFF regs_94 ( // @[RegFile.scala 66:20:@126306.4]
    .clock(regs_94_clock),
    .reset(regs_94_reset),
    .io_in(regs_94_io_in),
    .io_reset(regs_94_io_reset),
    .io_out(regs_94_io_out),
    .io_enable(regs_94_io_enable)
  );
  FringeFF regs_95 ( // @[RegFile.scala 66:20:@126320.4]
    .clock(regs_95_clock),
    .reset(regs_95_reset),
    .io_in(regs_95_io_in),
    .io_reset(regs_95_io_reset),
    .io_out(regs_95_io_out),
    .io_enable(regs_95_io_enable)
  );
  FringeFF regs_96 ( // @[RegFile.scala 66:20:@126334.4]
    .clock(regs_96_clock),
    .reset(regs_96_reset),
    .io_in(regs_96_io_in),
    .io_reset(regs_96_io_reset),
    .io_out(regs_96_io_out),
    .io_enable(regs_96_io_enable)
  );
  FringeFF regs_97 ( // @[RegFile.scala 66:20:@126348.4]
    .clock(regs_97_clock),
    .reset(regs_97_reset),
    .io_in(regs_97_io_in),
    .io_reset(regs_97_io_reset),
    .io_out(regs_97_io_out),
    .io_enable(regs_97_io_enable)
  );
  FringeFF regs_98 ( // @[RegFile.scala 66:20:@126362.4]
    .clock(regs_98_clock),
    .reset(regs_98_reset),
    .io_in(regs_98_io_in),
    .io_reset(regs_98_io_reset),
    .io_out(regs_98_io_out),
    .io_enable(regs_98_io_enable)
  );
  FringeFF regs_99 ( // @[RegFile.scala 66:20:@126376.4]
    .clock(regs_99_clock),
    .reset(regs_99_reset),
    .io_in(regs_99_io_in),
    .io_reset(regs_99_io_reset),
    .io_out(regs_99_io_out),
    .io_enable(regs_99_io_enable)
  );
  FringeFF regs_100 ( // @[RegFile.scala 66:20:@126390.4]
    .clock(regs_100_clock),
    .reset(regs_100_reset),
    .io_in(regs_100_io_in),
    .io_reset(regs_100_io_reset),
    .io_out(regs_100_io_out),
    .io_enable(regs_100_io_enable)
  );
  FringeFF regs_101 ( // @[RegFile.scala 66:20:@126404.4]
    .clock(regs_101_clock),
    .reset(regs_101_reset),
    .io_in(regs_101_io_in),
    .io_reset(regs_101_io_reset),
    .io_out(regs_101_io_out),
    .io_enable(regs_101_io_enable)
  );
  FringeFF regs_102 ( // @[RegFile.scala 66:20:@126418.4]
    .clock(regs_102_clock),
    .reset(regs_102_reset),
    .io_in(regs_102_io_in),
    .io_reset(regs_102_io_reset),
    .io_out(regs_102_io_out),
    .io_enable(regs_102_io_enable)
  );
  FringeFF regs_103 ( // @[RegFile.scala 66:20:@126432.4]
    .clock(regs_103_clock),
    .reset(regs_103_reset),
    .io_in(regs_103_io_in),
    .io_reset(regs_103_io_reset),
    .io_out(regs_103_io_out),
    .io_enable(regs_103_io_enable)
  );
  FringeFF regs_104 ( // @[RegFile.scala 66:20:@126446.4]
    .clock(regs_104_clock),
    .reset(regs_104_reset),
    .io_in(regs_104_io_in),
    .io_reset(regs_104_io_reset),
    .io_out(regs_104_io_out),
    .io_enable(regs_104_io_enable)
  );
  FringeFF regs_105 ( // @[RegFile.scala 66:20:@126460.4]
    .clock(regs_105_clock),
    .reset(regs_105_reset),
    .io_in(regs_105_io_in),
    .io_reset(regs_105_io_reset),
    .io_out(regs_105_io_out),
    .io_enable(regs_105_io_enable)
  );
  FringeFF regs_106 ( // @[RegFile.scala 66:20:@126474.4]
    .clock(regs_106_clock),
    .reset(regs_106_reset),
    .io_in(regs_106_io_in),
    .io_reset(regs_106_io_reset),
    .io_out(regs_106_io_out),
    .io_enable(regs_106_io_enable)
  );
  FringeFF regs_107 ( // @[RegFile.scala 66:20:@126488.4]
    .clock(regs_107_clock),
    .reset(regs_107_reset),
    .io_in(regs_107_io_in),
    .io_reset(regs_107_io_reset),
    .io_out(regs_107_io_out),
    .io_enable(regs_107_io_enable)
  );
  FringeFF regs_108 ( // @[RegFile.scala 66:20:@126502.4]
    .clock(regs_108_clock),
    .reset(regs_108_reset),
    .io_in(regs_108_io_in),
    .io_reset(regs_108_io_reset),
    .io_out(regs_108_io_out),
    .io_enable(regs_108_io_enable)
  );
  FringeFF regs_109 ( // @[RegFile.scala 66:20:@126516.4]
    .clock(regs_109_clock),
    .reset(regs_109_reset),
    .io_in(regs_109_io_in),
    .io_reset(regs_109_io_reset),
    .io_out(regs_109_io_out),
    .io_enable(regs_109_io_enable)
  );
  FringeFF regs_110 ( // @[RegFile.scala 66:20:@126530.4]
    .clock(regs_110_clock),
    .reset(regs_110_reset),
    .io_in(regs_110_io_in),
    .io_reset(regs_110_io_reset),
    .io_out(regs_110_io_out),
    .io_enable(regs_110_io_enable)
  );
  FringeFF regs_111 ( // @[RegFile.scala 66:20:@126544.4]
    .clock(regs_111_clock),
    .reset(regs_111_reset),
    .io_in(regs_111_io_in),
    .io_reset(regs_111_io_reset),
    .io_out(regs_111_io_out),
    .io_enable(regs_111_io_enable)
  );
  FringeFF regs_112 ( // @[RegFile.scala 66:20:@126558.4]
    .clock(regs_112_clock),
    .reset(regs_112_reset),
    .io_in(regs_112_io_in),
    .io_reset(regs_112_io_reset),
    .io_out(regs_112_io_out),
    .io_enable(regs_112_io_enable)
  );
  FringeFF regs_113 ( // @[RegFile.scala 66:20:@126572.4]
    .clock(regs_113_clock),
    .reset(regs_113_reset),
    .io_in(regs_113_io_in),
    .io_reset(regs_113_io_reset),
    .io_out(regs_113_io_out),
    .io_enable(regs_113_io_enable)
  );
  FringeFF regs_114 ( // @[RegFile.scala 66:20:@126586.4]
    .clock(regs_114_clock),
    .reset(regs_114_reset),
    .io_in(regs_114_io_in),
    .io_reset(regs_114_io_reset),
    .io_out(regs_114_io_out),
    .io_enable(regs_114_io_enable)
  );
  FringeFF regs_115 ( // @[RegFile.scala 66:20:@126600.4]
    .clock(regs_115_clock),
    .reset(regs_115_reset),
    .io_in(regs_115_io_in),
    .io_reset(regs_115_io_reset),
    .io_out(regs_115_io_out),
    .io_enable(regs_115_io_enable)
  );
  FringeFF regs_116 ( // @[RegFile.scala 66:20:@126614.4]
    .clock(regs_116_clock),
    .reset(regs_116_reset),
    .io_in(regs_116_io_in),
    .io_reset(regs_116_io_reset),
    .io_out(regs_116_io_out),
    .io_enable(regs_116_io_enable)
  );
  FringeFF regs_117 ( // @[RegFile.scala 66:20:@126628.4]
    .clock(regs_117_clock),
    .reset(regs_117_reset),
    .io_in(regs_117_io_in),
    .io_reset(regs_117_io_reset),
    .io_out(regs_117_io_out),
    .io_enable(regs_117_io_enable)
  );
  FringeFF regs_118 ( // @[RegFile.scala 66:20:@126642.4]
    .clock(regs_118_clock),
    .reset(regs_118_reset),
    .io_in(regs_118_io_in),
    .io_reset(regs_118_io_reset),
    .io_out(regs_118_io_out),
    .io_enable(regs_118_io_enable)
  );
  FringeFF regs_119 ( // @[RegFile.scala 66:20:@126656.4]
    .clock(regs_119_clock),
    .reset(regs_119_reset),
    .io_in(regs_119_io_in),
    .io_reset(regs_119_io_reset),
    .io_out(regs_119_io_out),
    .io_enable(regs_119_io_enable)
  );
  FringeFF regs_120 ( // @[RegFile.scala 66:20:@126670.4]
    .clock(regs_120_clock),
    .reset(regs_120_reset),
    .io_in(regs_120_io_in),
    .io_reset(regs_120_io_reset),
    .io_out(regs_120_io_out),
    .io_enable(regs_120_io_enable)
  );
  FringeFF regs_121 ( // @[RegFile.scala 66:20:@126684.4]
    .clock(regs_121_clock),
    .reset(regs_121_reset),
    .io_in(regs_121_io_in),
    .io_reset(regs_121_io_reset),
    .io_out(regs_121_io_out),
    .io_enable(regs_121_io_enable)
  );
  FringeFF regs_122 ( // @[RegFile.scala 66:20:@126698.4]
    .clock(regs_122_clock),
    .reset(regs_122_reset),
    .io_in(regs_122_io_in),
    .io_reset(regs_122_io_reset),
    .io_out(regs_122_io_out),
    .io_enable(regs_122_io_enable)
  );
  FringeFF regs_123 ( // @[RegFile.scala 66:20:@126712.4]
    .clock(regs_123_clock),
    .reset(regs_123_reset),
    .io_in(regs_123_io_in),
    .io_reset(regs_123_io_reset),
    .io_out(regs_123_io_out),
    .io_enable(regs_123_io_enable)
  );
  FringeFF regs_124 ( // @[RegFile.scala 66:20:@126726.4]
    .clock(regs_124_clock),
    .reset(regs_124_reset),
    .io_in(regs_124_io_in),
    .io_reset(regs_124_io_reset),
    .io_out(regs_124_io_out),
    .io_enable(regs_124_io_enable)
  );
  FringeFF regs_125 ( // @[RegFile.scala 66:20:@126740.4]
    .clock(regs_125_clock),
    .reset(regs_125_reset),
    .io_in(regs_125_io_in),
    .io_reset(regs_125_io_reset),
    .io_out(regs_125_io_out),
    .io_enable(regs_125_io_enable)
  );
  FringeFF regs_126 ( // @[RegFile.scala 66:20:@126754.4]
    .clock(regs_126_clock),
    .reset(regs_126_reset),
    .io_in(regs_126_io_in),
    .io_reset(regs_126_io_reset),
    .io_out(regs_126_io_out),
    .io_enable(regs_126_io_enable)
  );
  FringeFF regs_127 ( // @[RegFile.scala 66:20:@126768.4]
    .clock(regs_127_clock),
    .reset(regs_127_reset),
    .io_in(regs_127_io_in),
    .io_reset(regs_127_io_reset),
    .io_out(regs_127_io_out),
    .io_enable(regs_127_io_enable)
  );
  FringeFF regs_128 ( // @[RegFile.scala 66:20:@126782.4]
    .clock(regs_128_clock),
    .reset(regs_128_reset),
    .io_in(regs_128_io_in),
    .io_reset(regs_128_io_reset),
    .io_out(regs_128_io_out),
    .io_enable(regs_128_io_enable)
  );
  FringeFF regs_129 ( // @[RegFile.scala 66:20:@126796.4]
    .clock(regs_129_clock),
    .reset(regs_129_reset),
    .io_in(regs_129_io_in),
    .io_reset(regs_129_io_reset),
    .io_out(regs_129_io_out),
    .io_enable(regs_129_io_enable)
  );
  FringeFF regs_130 ( // @[RegFile.scala 66:20:@126810.4]
    .clock(regs_130_clock),
    .reset(regs_130_reset),
    .io_in(regs_130_io_in),
    .io_reset(regs_130_io_reset),
    .io_out(regs_130_io_out),
    .io_enable(regs_130_io_enable)
  );
  FringeFF regs_131 ( // @[RegFile.scala 66:20:@126824.4]
    .clock(regs_131_clock),
    .reset(regs_131_reset),
    .io_in(regs_131_io_in),
    .io_reset(regs_131_io_reset),
    .io_out(regs_131_io_out),
    .io_enable(regs_131_io_enable)
  );
  FringeFF regs_132 ( // @[RegFile.scala 66:20:@126838.4]
    .clock(regs_132_clock),
    .reset(regs_132_reset),
    .io_in(regs_132_io_in),
    .io_reset(regs_132_io_reset),
    .io_out(regs_132_io_out),
    .io_enable(regs_132_io_enable)
  );
  FringeFF regs_133 ( // @[RegFile.scala 66:20:@126852.4]
    .clock(regs_133_clock),
    .reset(regs_133_reset),
    .io_in(regs_133_io_in),
    .io_reset(regs_133_io_reset),
    .io_out(regs_133_io_out),
    .io_enable(regs_133_io_enable)
  );
  FringeFF regs_134 ( // @[RegFile.scala 66:20:@126866.4]
    .clock(regs_134_clock),
    .reset(regs_134_reset),
    .io_in(regs_134_io_in),
    .io_reset(regs_134_io_reset),
    .io_out(regs_134_io_out),
    .io_enable(regs_134_io_enable)
  );
  FringeFF regs_135 ( // @[RegFile.scala 66:20:@126880.4]
    .clock(regs_135_clock),
    .reset(regs_135_reset),
    .io_in(regs_135_io_in),
    .io_reset(regs_135_io_reset),
    .io_out(regs_135_io_out),
    .io_enable(regs_135_io_enable)
  );
  FringeFF regs_136 ( // @[RegFile.scala 66:20:@126894.4]
    .clock(regs_136_clock),
    .reset(regs_136_reset),
    .io_in(regs_136_io_in),
    .io_reset(regs_136_io_reset),
    .io_out(regs_136_io_out),
    .io_enable(regs_136_io_enable)
  );
  FringeFF regs_137 ( // @[RegFile.scala 66:20:@126908.4]
    .clock(regs_137_clock),
    .reset(regs_137_reset),
    .io_in(regs_137_io_in),
    .io_reset(regs_137_io_reset),
    .io_out(regs_137_io_out),
    .io_enable(regs_137_io_enable)
  );
  FringeFF regs_138 ( // @[RegFile.scala 66:20:@126922.4]
    .clock(regs_138_clock),
    .reset(regs_138_reset),
    .io_in(regs_138_io_in),
    .io_reset(regs_138_io_reset),
    .io_out(regs_138_io_out),
    .io_enable(regs_138_io_enable)
  );
  FringeFF regs_139 ( // @[RegFile.scala 66:20:@126936.4]
    .clock(regs_139_clock),
    .reset(regs_139_reset),
    .io_in(regs_139_io_in),
    .io_reset(regs_139_io_reset),
    .io_out(regs_139_io_out),
    .io_enable(regs_139_io_enable)
  );
  FringeFF regs_140 ( // @[RegFile.scala 66:20:@126950.4]
    .clock(regs_140_clock),
    .reset(regs_140_reset),
    .io_in(regs_140_io_in),
    .io_reset(regs_140_io_reset),
    .io_out(regs_140_io_out),
    .io_enable(regs_140_io_enable)
  );
  FringeFF regs_141 ( // @[RegFile.scala 66:20:@126964.4]
    .clock(regs_141_clock),
    .reset(regs_141_reset),
    .io_in(regs_141_io_in),
    .io_reset(regs_141_io_reset),
    .io_out(regs_141_io_out),
    .io_enable(regs_141_io_enable)
  );
  FringeFF regs_142 ( // @[RegFile.scala 66:20:@126978.4]
    .clock(regs_142_clock),
    .reset(regs_142_reset),
    .io_in(regs_142_io_in),
    .io_reset(regs_142_io_reset),
    .io_out(regs_142_io_out),
    .io_enable(regs_142_io_enable)
  );
  FringeFF regs_143 ( // @[RegFile.scala 66:20:@126992.4]
    .clock(regs_143_clock),
    .reset(regs_143_reset),
    .io_in(regs_143_io_in),
    .io_reset(regs_143_io_reset),
    .io_out(regs_143_io_out),
    .io_enable(regs_143_io_enable)
  );
  FringeFF regs_144 ( // @[RegFile.scala 66:20:@127006.4]
    .clock(regs_144_clock),
    .reset(regs_144_reset),
    .io_in(regs_144_io_in),
    .io_reset(regs_144_io_reset),
    .io_out(regs_144_io_out),
    .io_enable(regs_144_io_enable)
  );
  FringeFF regs_145 ( // @[RegFile.scala 66:20:@127020.4]
    .clock(regs_145_clock),
    .reset(regs_145_reset),
    .io_in(regs_145_io_in),
    .io_reset(regs_145_io_reset),
    .io_out(regs_145_io_out),
    .io_enable(regs_145_io_enable)
  );
  FringeFF regs_146 ( // @[RegFile.scala 66:20:@127034.4]
    .clock(regs_146_clock),
    .reset(regs_146_reset),
    .io_in(regs_146_io_in),
    .io_reset(regs_146_io_reset),
    .io_out(regs_146_io_out),
    .io_enable(regs_146_io_enable)
  );
  FringeFF regs_147 ( // @[RegFile.scala 66:20:@127048.4]
    .clock(regs_147_clock),
    .reset(regs_147_reset),
    .io_in(regs_147_io_in),
    .io_reset(regs_147_io_reset),
    .io_out(regs_147_io_out),
    .io_enable(regs_147_io_enable)
  );
  FringeFF regs_148 ( // @[RegFile.scala 66:20:@127062.4]
    .clock(regs_148_clock),
    .reset(regs_148_reset),
    .io_in(regs_148_io_in),
    .io_reset(regs_148_io_reset),
    .io_out(regs_148_io_out),
    .io_enable(regs_148_io_enable)
  );
  FringeFF regs_149 ( // @[RegFile.scala 66:20:@127076.4]
    .clock(regs_149_clock),
    .reset(regs_149_reset),
    .io_in(regs_149_io_in),
    .io_reset(regs_149_io_reset),
    .io_out(regs_149_io_out),
    .io_enable(regs_149_io_enable)
  );
  FringeFF regs_150 ( // @[RegFile.scala 66:20:@127090.4]
    .clock(regs_150_clock),
    .reset(regs_150_reset),
    .io_in(regs_150_io_in),
    .io_reset(regs_150_io_reset),
    .io_out(regs_150_io_out),
    .io_enable(regs_150_io_enable)
  );
  FringeFF regs_151 ( // @[RegFile.scala 66:20:@127104.4]
    .clock(regs_151_clock),
    .reset(regs_151_reset),
    .io_in(regs_151_io_in),
    .io_reset(regs_151_io_reset),
    .io_out(regs_151_io_out),
    .io_enable(regs_151_io_enable)
  );
  FringeFF regs_152 ( // @[RegFile.scala 66:20:@127118.4]
    .clock(regs_152_clock),
    .reset(regs_152_reset),
    .io_in(regs_152_io_in),
    .io_reset(regs_152_io_reset),
    .io_out(regs_152_io_out),
    .io_enable(regs_152_io_enable)
  );
  FringeFF regs_153 ( // @[RegFile.scala 66:20:@127132.4]
    .clock(regs_153_clock),
    .reset(regs_153_reset),
    .io_in(regs_153_io_in),
    .io_reset(regs_153_io_reset),
    .io_out(regs_153_io_out),
    .io_enable(regs_153_io_enable)
  );
  FringeFF regs_154 ( // @[RegFile.scala 66:20:@127146.4]
    .clock(regs_154_clock),
    .reset(regs_154_reset),
    .io_in(regs_154_io_in),
    .io_reset(regs_154_io_reset),
    .io_out(regs_154_io_out),
    .io_enable(regs_154_io_enable)
  );
  FringeFF regs_155 ( // @[RegFile.scala 66:20:@127160.4]
    .clock(regs_155_clock),
    .reset(regs_155_reset),
    .io_in(regs_155_io_in),
    .io_reset(regs_155_io_reset),
    .io_out(regs_155_io_out),
    .io_enable(regs_155_io_enable)
  );
  FringeFF regs_156 ( // @[RegFile.scala 66:20:@127174.4]
    .clock(regs_156_clock),
    .reset(regs_156_reset),
    .io_in(regs_156_io_in),
    .io_reset(regs_156_io_reset),
    .io_out(regs_156_io_out),
    .io_enable(regs_156_io_enable)
  );
  FringeFF regs_157 ( // @[RegFile.scala 66:20:@127188.4]
    .clock(regs_157_clock),
    .reset(regs_157_reset),
    .io_in(regs_157_io_in),
    .io_reset(regs_157_io_reset),
    .io_out(regs_157_io_out),
    .io_enable(regs_157_io_enable)
  );
  FringeFF regs_158 ( // @[RegFile.scala 66:20:@127202.4]
    .clock(regs_158_clock),
    .reset(regs_158_reset),
    .io_in(regs_158_io_in),
    .io_reset(regs_158_io_reset),
    .io_out(regs_158_io_out),
    .io_enable(regs_158_io_enable)
  );
  FringeFF regs_159 ( // @[RegFile.scala 66:20:@127216.4]
    .clock(regs_159_clock),
    .reset(regs_159_reset),
    .io_in(regs_159_io_in),
    .io_reset(regs_159_io_reset),
    .io_out(regs_159_io_out),
    .io_enable(regs_159_io_enable)
  );
  FringeFF regs_160 ( // @[RegFile.scala 66:20:@127230.4]
    .clock(regs_160_clock),
    .reset(regs_160_reset),
    .io_in(regs_160_io_in),
    .io_reset(regs_160_io_reset),
    .io_out(regs_160_io_out),
    .io_enable(regs_160_io_enable)
  );
  FringeFF regs_161 ( // @[RegFile.scala 66:20:@127244.4]
    .clock(regs_161_clock),
    .reset(regs_161_reset),
    .io_in(regs_161_io_in),
    .io_reset(regs_161_io_reset),
    .io_out(regs_161_io_out),
    .io_enable(regs_161_io_enable)
  );
  FringeFF regs_162 ( // @[RegFile.scala 66:20:@127258.4]
    .clock(regs_162_clock),
    .reset(regs_162_reset),
    .io_in(regs_162_io_in),
    .io_reset(regs_162_io_reset),
    .io_out(regs_162_io_out),
    .io_enable(regs_162_io_enable)
  );
  FringeFF regs_163 ( // @[RegFile.scala 66:20:@127272.4]
    .clock(regs_163_clock),
    .reset(regs_163_reset),
    .io_in(regs_163_io_in),
    .io_reset(regs_163_io_reset),
    .io_out(regs_163_io_out),
    .io_enable(regs_163_io_enable)
  );
  FringeFF regs_164 ( // @[RegFile.scala 66:20:@127286.4]
    .clock(regs_164_clock),
    .reset(regs_164_reset),
    .io_in(regs_164_io_in),
    .io_reset(regs_164_io_reset),
    .io_out(regs_164_io_out),
    .io_enable(regs_164_io_enable)
  );
  FringeFF regs_165 ( // @[RegFile.scala 66:20:@127300.4]
    .clock(regs_165_clock),
    .reset(regs_165_reset),
    .io_in(regs_165_io_in),
    .io_reset(regs_165_io_reset),
    .io_out(regs_165_io_out),
    .io_enable(regs_165_io_enable)
  );
  FringeFF regs_166 ( // @[RegFile.scala 66:20:@127314.4]
    .clock(regs_166_clock),
    .reset(regs_166_reset),
    .io_in(regs_166_io_in),
    .io_reset(regs_166_io_reset),
    .io_out(regs_166_io_out),
    .io_enable(regs_166_io_enable)
  );
  FringeFF regs_167 ( // @[RegFile.scala 66:20:@127328.4]
    .clock(regs_167_clock),
    .reset(regs_167_reset),
    .io_in(regs_167_io_in),
    .io_reset(regs_167_io_reset),
    .io_out(regs_167_io_out),
    .io_enable(regs_167_io_enable)
  );
  FringeFF regs_168 ( // @[RegFile.scala 66:20:@127342.4]
    .clock(regs_168_clock),
    .reset(regs_168_reset),
    .io_in(regs_168_io_in),
    .io_reset(regs_168_io_reset),
    .io_out(regs_168_io_out),
    .io_enable(regs_168_io_enable)
  );
  FringeFF regs_169 ( // @[RegFile.scala 66:20:@127356.4]
    .clock(regs_169_clock),
    .reset(regs_169_reset),
    .io_in(regs_169_io_in),
    .io_reset(regs_169_io_reset),
    .io_out(regs_169_io_out),
    .io_enable(regs_169_io_enable)
  );
  FringeFF regs_170 ( // @[RegFile.scala 66:20:@127370.4]
    .clock(regs_170_clock),
    .reset(regs_170_reset),
    .io_in(regs_170_io_in),
    .io_reset(regs_170_io_reset),
    .io_out(regs_170_io_out),
    .io_enable(regs_170_io_enable)
  );
  FringeFF regs_171 ( // @[RegFile.scala 66:20:@127384.4]
    .clock(regs_171_clock),
    .reset(regs_171_reset),
    .io_in(regs_171_io_in),
    .io_reset(regs_171_io_reset),
    .io_out(regs_171_io_out),
    .io_enable(regs_171_io_enable)
  );
  FringeFF regs_172 ( // @[RegFile.scala 66:20:@127398.4]
    .clock(regs_172_clock),
    .reset(regs_172_reset),
    .io_in(regs_172_io_in),
    .io_reset(regs_172_io_reset),
    .io_out(regs_172_io_out),
    .io_enable(regs_172_io_enable)
  );
  FringeFF regs_173 ( // @[RegFile.scala 66:20:@127412.4]
    .clock(regs_173_clock),
    .reset(regs_173_reset),
    .io_in(regs_173_io_in),
    .io_reset(regs_173_io_reset),
    .io_out(regs_173_io_out),
    .io_enable(regs_173_io_enable)
  );
  FringeFF regs_174 ( // @[RegFile.scala 66:20:@127426.4]
    .clock(regs_174_clock),
    .reset(regs_174_reset),
    .io_in(regs_174_io_in),
    .io_reset(regs_174_io_reset),
    .io_out(regs_174_io_out),
    .io_enable(regs_174_io_enable)
  );
  FringeFF regs_175 ( // @[RegFile.scala 66:20:@127440.4]
    .clock(regs_175_clock),
    .reset(regs_175_reset),
    .io_in(regs_175_io_in),
    .io_reset(regs_175_io_reset),
    .io_out(regs_175_io_out),
    .io_enable(regs_175_io_enable)
  );
  FringeFF regs_176 ( // @[RegFile.scala 66:20:@127454.4]
    .clock(regs_176_clock),
    .reset(regs_176_reset),
    .io_in(regs_176_io_in),
    .io_reset(regs_176_io_reset),
    .io_out(regs_176_io_out),
    .io_enable(regs_176_io_enable)
  );
  FringeFF regs_177 ( // @[RegFile.scala 66:20:@127468.4]
    .clock(regs_177_clock),
    .reset(regs_177_reset),
    .io_in(regs_177_io_in),
    .io_reset(regs_177_io_reset),
    .io_out(regs_177_io_out),
    .io_enable(regs_177_io_enable)
  );
  FringeFF regs_178 ( // @[RegFile.scala 66:20:@127482.4]
    .clock(regs_178_clock),
    .reset(regs_178_reset),
    .io_in(regs_178_io_in),
    .io_reset(regs_178_io_reset),
    .io_out(regs_178_io_out),
    .io_enable(regs_178_io_enable)
  );
  FringeFF regs_179 ( // @[RegFile.scala 66:20:@127496.4]
    .clock(regs_179_clock),
    .reset(regs_179_reset),
    .io_in(regs_179_io_in),
    .io_reset(regs_179_io_reset),
    .io_out(regs_179_io_out),
    .io_enable(regs_179_io_enable)
  );
  FringeFF regs_180 ( // @[RegFile.scala 66:20:@127510.4]
    .clock(regs_180_clock),
    .reset(regs_180_reset),
    .io_in(regs_180_io_in),
    .io_reset(regs_180_io_reset),
    .io_out(regs_180_io_out),
    .io_enable(regs_180_io_enable)
  );
  FringeFF regs_181 ( // @[RegFile.scala 66:20:@127524.4]
    .clock(regs_181_clock),
    .reset(regs_181_reset),
    .io_in(regs_181_io_in),
    .io_reset(regs_181_io_reset),
    .io_out(regs_181_io_out),
    .io_enable(regs_181_io_enable)
  );
  FringeFF regs_182 ( // @[RegFile.scala 66:20:@127538.4]
    .clock(regs_182_clock),
    .reset(regs_182_reset),
    .io_in(regs_182_io_in),
    .io_reset(regs_182_io_reset),
    .io_out(regs_182_io_out),
    .io_enable(regs_182_io_enable)
  );
  FringeFF regs_183 ( // @[RegFile.scala 66:20:@127552.4]
    .clock(regs_183_clock),
    .reset(regs_183_reset),
    .io_in(regs_183_io_in),
    .io_reset(regs_183_io_reset),
    .io_out(regs_183_io_out),
    .io_enable(regs_183_io_enable)
  );
  FringeFF regs_184 ( // @[RegFile.scala 66:20:@127566.4]
    .clock(regs_184_clock),
    .reset(regs_184_reset),
    .io_in(regs_184_io_in),
    .io_reset(regs_184_io_reset),
    .io_out(regs_184_io_out),
    .io_enable(regs_184_io_enable)
  );
  FringeFF regs_185 ( // @[RegFile.scala 66:20:@127580.4]
    .clock(regs_185_clock),
    .reset(regs_185_reset),
    .io_in(regs_185_io_in),
    .io_reset(regs_185_io_reset),
    .io_out(regs_185_io_out),
    .io_enable(regs_185_io_enable)
  );
  FringeFF regs_186 ( // @[RegFile.scala 66:20:@127594.4]
    .clock(regs_186_clock),
    .reset(regs_186_reset),
    .io_in(regs_186_io_in),
    .io_reset(regs_186_io_reset),
    .io_out(regs_186_io_out),
    .io_enable(regs_186_io_enable)
  );
  FringeFF regs_187 ( // @[RegFile.scala 66:20:@127608.4]
    .clock(regs_187_clock),
    .reset(regs_187_reset),
    .io_in(regs_187_io_in),
    .io_reset(regs_187_io_reset),
    .io_out(regs_187_io_out),
    .io_enable(regs_187_io_enable)
  );
  FringeFF regs_188 ( // @[RegFile.scala 66:20:@127622.4]
    .clock(regs_188_clock),
    .reset(regs_188_reset),
    .io_in(regs_188_io_in),
    .io_reset(regs_188_io_reset),
    .io_out(regs_188_io_out),
    .io_enable(regs_188_io_enable)
  );
  FringeFF regs_189 ( // @[RegFile.scala 66:20:@127636.4]
    .clock(regs_189_clock),
    .reset(regs_189_reset),
    .io_in(regs_189_io_in),
    .io_reset(regs_189_io_reset),
    .io_out(regs_189_io_out),
    .io_enable(regs_189_io_enable)
  );
  FringeFF regs_190 ( // @[RegFile.scala 66:20:@127650.4]
    .clock(regs_190_clock),
    .reset(regs_190_reset),
    .io_in(regs_190_io_in),
    .io_reset(regs_190_io_reset),
    .io_out(regs_190_io_out),
    .io_enable(regs_190_io_enable)
  );
  FringeFF regs_191 ( // @[RegFile.scala 66:20:@127664.4]
    .clock(regs_191_clock),
    .reset(regs_191_reset),
    .io_in(regs_191_io_in),
    .io_reset(regs_191_io_reset),
    .io_out(regs_191_io_out),
    .io_enable(regs_191_io_enable)
  );
  FringeFF regs_192 ( // @[RegFile.scala 66:20:@127678.4]
    .clock(regs_192_clock),
    .reset(regs_192_reset),
    .io_in(regs_192_io_in),
    .io_reset(regs_192_io_reset),
    .io_out(regs_192_io_out),
    .io_enable(regs_192_io_enable)
  );
  FringeFF regs_193 ( // @[RegFile.scala 66:20:@127692.4]
    .clock(regs_193_clock),
    .reset(regs_193_reset),
    .io_in(regs_193_io_in),
    .io_reset(regs_193_io_reset),
    .io_out(regs_193_io_out),
    .io_enable(regs_193_io_enable)
  );
  FringeFF regs_194 ( // @[RegFile.scala 66:20:@127706.4]
    .clock(regs_194_clock),
    .reset(regs_194_reset),
    .io_in(regs_194_io_in),
    .io_reset(regs_194_io_reset),
    .io_out(regs_194_io_out),
    .io_enable(regs_194_io_enable)
  );
  FringeFF regs_195 ( // @[RegFile.scala 66:20:@127720.4]
    .clock(regs_195_clock),
    .reset(regs_195_reset),
    .io_in(regs_195_io_in),
    .io_reset(regs_195_io_reset),
    .io_out(regs_195_io_out),
    .io_enable(regs_195_io_enable)
  );
  FringeFF regs_196 ( // @[RegFile.scala 66:20:@127734.4]
    .clock(regs_196_clock),
    .reset(regs_196_reset),
    .io_in(regs_196_io_in),
    .io_reset(regs_196_io_reset),
    .io_out(regs_196_io_out),
    .io_enable(regs_196_io_enable)
  );
  FringeFF regs_197 ( // @[RegFile.scala 66:20:@127748.4]
    .clock(regs_197_clock),
    .reset(regs_197_reset),
    .io_in(regs_197_io_in),
    .io_reset(regs_197_io_reset),
    .io_out(regs_197_io_out),
    .io_enable(regs_197_io_enable)
  );
  FringeFF regs_198 ( // @[RegFile.scala 66:20:@127762.4]
    .clock(regs_198_clock),
    .reset(regs_198_reset),
    .io_in(regs_198_io_in),
    .io_reset(regs_198_io_reset),
    .io_out(regs_198_io_out),
    .io_enable(regs_198_io_enable)
  );
  FringeFF regs_199 ( // @[RegFile.scala 66:20:@127776.4]
    .clock(regs_199_clock),
    .reset(regs_199_reset),
    .io_in(regs_199_io_in),
    .io_reset(regs_199_io_reset),
    .io_out(regs_199_io_out),
    .io_enable(regs_199_io_enable)
  );
  FringeFF regs_200 ( // @[RegFile.scala 66:20:@127790.4]
    .clock(regs_200_clock),
    .reset(regs_200_reset),
    .io_in(regs_200_io_in),
    .io_reset(regs_200_io_reset),
    .io_out(regs_200_io_out),
    .io_enable(regs_200_io_enable)
  );
  FringeFF regs_201 ( // @[RegFile.scala 66:20:@127804.4]
    .clock(regs_201_clock),
    .reset(regs_201_reset),
    .io_in(regs_201_io_in),
    .io_reset(regs_201_io_reset),
    .io_out(regs_201_io_out),
    .io_enable(regs_201_io_enable)
  );
  FringeFF regs_202 ( // @[RegFile.scala 66:20:@127818.4]
    .clock(regs_202_clock),
    .reset(regs_202_reset),
    .io_in(regs_202_io_in),
    .io_reset(regs_202_io_reset),
    .io_out(regs_202_io_out),
    .io_enable(regs_202_io_enable)
  );
  FringeFF regs_203 ( // @[RegFile.scala 66:20:@127832.4]
    .clock(regs_203_clock),
    .reset(regs_203_reset),
    .io_in(regs_203_io_in),
    .io_reset(regs_203_io_reset),
    .io_out(regs_203_io_out),
    .io_enable(regs_203_io_enable)
  );
  FringeFF regs_204 ( // @[RegFile.scala 66:20:@127846.4]
    .clock(regs_204_clock),
    .reset(regs_204_reset),
    .io_in(regs_204_io_in),
    .io_reset(regs_204_io_reset),
    .io_out(regs_204_io_out),
    .io_enable(regs_204_io_enable)
  );
  FringeFF regs_205 ( // @[RegFile.scala 66:20:@127860.4]
    .clock(regs_205_clock),
    .reset(regs_205_reset),
    .io_in(regs_205_io_in),
    .io_reset(regs_205_io_reset),
    .io_out(regs_205_io_out),
    .io_enable(regs_205_io_enable)
  );
  FringeFF regs_206 ( // @[RegFile.scala 66:20:@127874.4]
    .clock(regs_206_clock),
    .reset(regs_206_reset),
    .io_in(regs_206_io_in),
    .io_reset(regs_206_io_reset),
    .io_out(regs_206_io_out),
    .io_enable(regs_206_io_enable)
  );
  FringeFF regs_207 ( // @[RegFile.scala 66:20:@127888.4]
    .clock(regs_207_clock),
    .reset(regs_207_reset),
    .io_in(regs_207_io_in),
    .io_reset(regs_207_io_reset),
    .io_out(regs_207_io_out),
    .io_enable(regs_207_io_enable)
  );
  FringeFF regs_208 ( // @[RegFile.scala 66:20:@127902.4]
    .clock(regs_208_clock),
    .reset(regs_208_reset),
    .io_in(regs_208_io_in),
    .io_reset(regs_208_io_reset),
    .io_out(regs_208_io_out),
    .io_enable(regs_208_io_enable)
  );
  FringeFF regs_209 ( // @[RegFile.scala 66:20:@127916.4]
    .clock(regs_209_clock),
    .reset(regs_209_reset),
    .io_in(regs_209_io_in),
    .io_reset(regs_209_io_reset),
    .io_out(regs_209_io_out),
    .io_enable(regs_209_io_enable)
  );
  FringeFF regs_210 ( // @[RegFile.scala 66:20:@127930.4]
    .clock(regs_210_clock),
    .reset(regs_210_reset),
    .io_in(regs_210_io_in),
    .io_reset(regs_210_io_reset),
    .io_out(regs_210_io_out),
    .io_enable(regs_210_io_enable)
  );
  FringeFF regs_211 ( // @[RegFile.scala 66:20:@127944.4]
    .clock(regs_211_clock),
    .reset(regs_211_reset),
    .io_in(regs_211_io_in),
    .io_reset(regs_211_io_reset),
    .io_out(regs_211_io_out),
    .io_enable(regs_211_io_enable)
  );
  FringeFF regs_212 ( // @[RegFile.scala 66:20:@127958.4]
    .clock(regs_212_clock),
    .reset(regs_212_reset),
    .io_in(regs_212_io_in),
    .io_reset(regs_212_io_reset),
    .io_out(regs_212_io_out),
    .io_enable(regs_212_io_enable)
  );
  FringeFF regs_213 ( // @[RegFile.scala 66:20:@127972.4]
    .clock(regs_213_clock),
    .reset(regs_213_reset),
    .io_in(regs_213_io_in),
    .io_reset(regs_213_io_reset),
    .io_out(regs_213_io_out),
    .io_enable(regs_213_io_enable)
  );
  FringeFF regs_214 ( // @[RegFile.scala 66:20:@127986.4]
    .clock(regs_214_clock),
    .reset(regs_214_reset),
    .io_in(regs_214_io_in),
    .io_reset(regs_214_io_reset),
    .io_out(regs_214_io_out),
    .io_enable(regs_214_io_enable)
  );
  FringeFF regs_215 ( // @[RegFile.scala 66:20:@128000.4]
    .clock(regs_215_clock),
    .reset(regs_215_reset),
    .io_in(regs_215_io_in),
    .io_reset(regs_215_io_reset),
    .io_out(regs_215_io_out),
    .io_enable(regs_215_io_enable)
  );
  FringeFF regs_216 ( // @[RegFile.scala 66:20:@128014.4]
    .clock(regs_216_clock),
    .reset(regs_216_reset),
    .io_in(regs_216_io_in),
    .io_reset(regs_216_io_reset),
    .io_out(regs_216_io_out),
    .io_enable(regs_216_io_enable)
  );
  FringeFF regs_217 ( // @[RegFile.scala 66:20:@128028.4]
    .clock(regs_217_clock),
    .reset(regs_217_reset),
    .io_in(regs_217_io_in),
    .io_reset(regs_217_io_reset),
    .io_out(regs_217_io_out),
    .io_enable(regs_217_io_enable)
  );
  FringeFF regs_218 ( // @[RegFile.scala 66:20:@128042.4]
    .clock(regs_218_clock),
    .reset(regs_218_reset),
    .io_in(regs_218_io_in),
    .io_reset(regs_218_io_reset),
    .io_out(regs_218_io_out),
    .io_enable(regs_218_io_enable)
  );
  FringeFF regs_219 ( // @[RegFile.scala 66:20:@128056.4]
    .clock(regs_219_clock),
    .reset(regs_219_reset),
    .io_in(regs_219_io_in),
    .io_reset(regs_219_io_reset),
    .io_out(regs_219_io_out),
    .io_enable(regs_219_io_enable)
  );
  FringeFF regs_220 ( // @[RegFile.scala 66:20:@128070.4]
    .clock(regs_220_clock),
    .reset(regs_220_reset),
    .io_in(regs_220_io_in),
    .io_reset(regs_220_io_reset),
    .io_out(regs_220_io_out),
    .io_enable(regs_220_io_enable)
  );
  FringeFF regs_221 ( // @[RegFile.scala 66:20:@128084.4]
    .clock(regs_221_clock),
    .reset(regs_221_reset),
    .io_in(regs_221_io_in),
    .io_reset(regs_221_io_reset),
    .io_out(regs_221_io_out),
    .io_enable(regs_221_io_enable)
  );
  FringeFF regs_222 ( // @[RegFile.scala 66:20:@128098.4]
    .clock(regs_222_clock),
    .reset(regs_222_reset),
    .io_in(regs_222_io_in),
    .io_reset(regs_222_io_reset),
    .io_out(regs_222_io_out),
    .io_enable(regs_222_io_enable)
  );
  FringeFF regs_223 ( // @[RegFile.scala 66:20:@128112.4]
    .clock(regs_223_clock),
    .reset(regs_223_reset),
    .io_in(regs_223_io_in),
    .io_reset(regs_223_io_reset),
    .io_out(regs_223_io_out),
    .io_enable(regs_223_io_enable)
  );
  FringeFF regs_224 ( // @[RegFile.scala 66:20:@128126.4]
    .clock(regs_224_clock),
    .reset(regs_224_reset),
    .io_in(regs_224_io_in),
    .io_reset(regs_224_io_reset),
    .io_out(regs_224_io_out),
    .io_enable(regs_224_io_enable)
  );
  FringeFF regs_225 ( // @[RegFile.scala 66:20:@128140.4]
    .clock(regs_225_clock),
    .reset(regs_225_reset),
    .io_in(regs_225_io_in),
    .io_reset(regs_225_io_reset),
    .io_out(regs_225_io_out),
    .io_enable(regs_225_io_enable)
  );
  FringeFF regs_226 ( // @[RegFile.scala 66:20:@128154.4]
    .clock(regs_226_clock),
    .reset(regs_226_reset),
    .io_in(regs_226_io_in),
    .io_reset(regs_226_io_reset),
    .io_out(regs_226_io_out),
    .io_enable(regs_226_io_enable)
  );
  FringeFF regs_227 ( // @[RegFile.scala 66:20:@128168.4]
    .clock(regs_227_clock),
    .reset(regs_227_reset),
    .io_in(regs_227_io_in),
    .io_reset(regs_227_io_reset),
    .io_out(regs_227_io_out),
    .io_enable(regs_227_io_enable)
  );
  FringeFF regs_228 ( // @[RegFile.scala 66:20:@128182.4]
    .clock(regs_228_clock),
    .reset(regs_228_reset),
    .io_in(regs_228_io_in),
    .io_reset(regs_228_io_reset),
    .io_out(regs_228_io_out),
    .io_enable(regs_228_io_enable)
  );
  FringeFF regs_229 ( // @[RegFile.scala 66:20:@128196.4]
    .clock(regs_229_clock),
    .reset(regs_229_reset),
    .io_in(regs_229_io_in),
    .io_reset(regs_229_io_reset),
    .io_out(regs_229_io_out),
    .io_enable(regs_229_io_enable)
  );
  FringeFF regs_230 ( // @[RegFile.scala 66:20:@128210.4]
    .clock(regs_230_clock),
    .reset(regs_230_reset),
    .io_in(regs_230_io_in),
    .io_reset(regs_230_io_reset),
    .io_out(regs_230_io_out),
    .io_enable(regs_230_io_enable)
  );
  FringeFF regs_231 ( // @[RegFile.scala 66:20:@128224.4]
    .clock(regs_231_clock),
    .reset(regs_231_reset),
    .io_in(regs_231_io_in),
    .io_reset(regs_231_io_reset),
    .io_out(regs_231_io_out),
    .io_enable(regs_231_io_enable)
  );
  FringeFF regs_232 ( // @[RegFile.scala 66:20:@128238.4]
    .clock(regs_232_clock),
    .reset(regs_232_reset),
    .io_in(regs_232_io_in),
    .io_reset(regs_232_io_reset),
    .io_out(regs_232_io_out),
    .io_enable(regs_232_io_enable)
  );
  FringeFF regs_233 ( // @[RegFile.scala 66:20:@128252.4]
    .clock(regs_233_clock),
    .reset(regs_233_reset),
    .io_in(regs_233_io_in),
    .io_reset(regs_233_io_reset),
    .io_out(regs_233_io_out),
    .io_enable(regs_233_io_enable)
  );
  FringeFF regs_234 ( // @[RegFile.scala 66:20:@128266.4]
    .clock(regs_234_clock),
    .reset(regs_234_reset),
    .io_in(regs_234_io_in),
    .io_reset(regs_234_io_reset),
    .io_out(regs_234_io_out),
    .io_enable(regs_234_io_enable)
  );
  FringeFF regs_235 ( // @[RegFile.scala 66:20:@128280.4]
    .clock(regs_235_clock),
    .reset(regs_235_reset),
    .io_in(regs_235_io_in),
    .io_reset(regs_235_io_reset),
    .io_out(regs_235_io_out),
    .io_enable(regs_235_io_enable)
  );
  FringeFF regs_236 ( // @[RegFile.scala 66:20:@128294.4]
    .clock(regs_236_clock),
    .reset(regs_236_reset),
    .io_in(regs_236_io_in),
    .io_reset(regs_236_io_reset),
    .io_out(regs_236_io_out),
    .io_enable(regs_236_io_enable)
  );
  FringeFF regs_237 ( // @[RegFile.scala 66:20:@128308.4]
    .clock(regs_237_clock),
    .reset(regs_237_reset),
    .io_in(regs_237_io_in),
    .io_reset(regs_237_io_reset),
    .io_out(regs_237_io_out),
    .io_enable(regs_237_io_enable)
  );
  FringeFF regs_238 ( // @[RegFile.scala 66:20:@128322.4]
    .clock(regs_238_clock),
    .reset(regs_238_reset),
    .io_in(regs_238_io_in),
    .io_reset(regs_238_io_reset),
    .io_out(regs_238_io_out),
    .io_enable(regs_238_io_enable)
  );
  FringeFF regs_239 ( // @[RegFile.scala 66:20:@128336.4]
    .clock(regs_239_clock),
    .reset(regs_239_reset),
    .io_in(regs_239_io_in),
    .io_reset(regs_239_io_reset),
    .io_out(regs_239_io_out),
    .io_enable(regs_239_io_enable)
  );
  FringeFF regs_240 ( // @[RegFile.scala 66:20:@128350.4]
    .clock(regs_240_clock),
    .reset(regs_240_reset),
    .io_in(regs_240_io_in),
    .io_reset(regs_240_io_reset),
    .io_out(regs_240_io_out),
    .io_enable(regs_240_io_enable)
  );
  FringeFF regs_241 ( // @[RegFile.scala 66:20:@128364.4]
    .clock(regs_241_clock),
    .reset(regs_241_reset),
    .io_in(regs_241_io_in),
    .io_reset(regs_241_io_reset),
    .io_out(regs_241_io_out),
    .io_enable(regs_241_io_enable)
  );
  FringeFF regs_242 ( // @[RegFile.scala 66:20:@128378.4]
    .clock(regs_242_clock),
    .reset(regs_242_reset),
    .io_in(regs_242_io_in),
    .io_reset(regs_242_io_reset),
    .io_out(regs_242_io_out),
    .io_enable(regs_242_io_enable)
  );
  FringeFF regs_243 ( // @[RegFile.scala 66:20:@128392.4]
    .clock(regs_243_clock),
    .reset(regs_243_reset),
    .io_in(regs_243_io_in),
    .io_reset(regs_243_io_reset),
    .io_out(regs_243_io_out),
    .io_enable(regs_243_io_enable)
  );
  FringeFF regs_244 ( // @[RegFile.scala 66:20:@128406.4]
    .clock(regs_244_clock),
    .reset(regs_244_reset),
    .io_in(regs_244_io_in),
    .io_reset(regs_244_io_reset),
    .io_out(regs_244_io_out),
    .io_enable(regs_244_io_enable)
  );
  FringeFF regs_245 ( // @[RegFile.scala 66:20:@128420.4]
    .clock(regs_245_clock),
    .reset(regs_245_reset),
    .io_in(regs_245_io_in),
    .io_reset(regs_245_io_reset),
    .io_out(regs_245_io_out),
    .io_enable(regs_245_io_enable)
  );
  FringeFF regs_246 ( // @[RegFile.scala 66:20:@128434.4]
    .clock(regs_246_clock),
    .reset(regs_246_reset),
    .io_in(regs_246_io_in),
    .io_reset(regs_246_io_reset),
    .io_out(regs_246_io_out),
    .io_enable(regs_246_io_enable)
  );
  FringeFF regs_247 ( // @[RegFile.scala 66:20:@128448.4]
    .clock(regs_247_clock),
    .reset(regs_247_reset),
    .io_in(regs_247_io_in),
    .io_reset(regs_247_io_reset),
    .io_out(regs_247_io_out),
    .io_enable(regs_247_io_enable)
  );
  FringeFF regs_248 ( // @[RegFile.scala 66:20:@128462.4]
    .clock(regs_248_clock),
    .reset(regs_248_reset),
    .io_in(regs_248_io_in),
    .io_reset(regs_248_io_reset),
    .io_out(regs_248_io_out),
    .io_enable(regs_248_io_enable)
  );
  FringeFF regs_249 ( // @[RegFile.scala 66:20:@128476.4]
    .clock(regs_249_clock),
    .reset(regs_249_reset),
    .io_in(regs_249_io_in),
    .io_reset(regs_249_io_reset),
    .io_out(regs_249_io_out),
    .io_enable(regs_249_io_enable)
  );
  FringeFF regs_250 ( // @[RegFile.scala 66:20:@128490.4]
    .clock(regs_250_clock),
    .reset(regs_250_reset),
    .io_in(regs_250_io_in),
    .io_reset(regs_250_io_reset),
    .io_out(regs_250_io_out),
    .io_enable(regs_250_io_enable)
  );
  FringeFF regs_251 ( // @[RegFile.scala 66:20:@128504.4]
    .clock(regs_251_clock),
    .reset(regs_251_reset),
    .io_in(regs_251_io_in),
    .io_reset(regs_251_io_reset),
    .io_out(regs_251_io_out),
    .io_enable(regs_251_io_enable)
  );
  FringeFF regs_252 ( // @[RegFile.scala 66:20:@128518.4]
    .clock(regs_252_clock),
    .reset(regs_252_reset),
    .io_in(regs_252_io_in),
    .io_reset(regs_252_io_reset),
    .io_out(regs_252_io_out),
    .io_enable(regs_252_io_enable)
  );
  FringeFF regs_253 ( // @[RegFile.scala 66:20:@128532.4]
    .clock(regs_253_clock),
    .reset(regs_253_reset),
    .io_in(regs_253_io_in),
    .io_reset(regs_253_io_reset),
    .io_out(regs_253_io_out),
    .io_enable(regs_253_io_enable)
  );
  FringeFF regs_254 ( // @[RegFile.scala 66:20:@128546.4]
    .clock(regs_254_clock),
    .reset(regs_254_reset),
    .io_in(regs_254_io_in),
    .io_reset(regs_254_io_reset),
    .io_out(regs_254_io_out),
    .io_enable(regs_254_io_enable)
  );
  FringeFF regs_255 ( // @[RegFile.scala 66:20:@128560.4]
    .clock(regs_255_clock),
    .reset(regs_255_reset),
    .io_in(regs_255_io_in),
    .io_reset(regs_255_io_reset),
    .io_out(regs_255_io_out),
    .io_enable(regs_255_io_enable)
  );
  FringeFF regs_256 ( // @[RegFile.scala 66:20:@128574.4]
    .clock(regs_256_clock),
    .reset(regs_256_reset),
    .io_in(regs_256_io_in),
    .io_reset(regs_256_io_reset),
    .io_out(regs_256_io_out),
    .io_enable(regs_256_io_enable)
  );
  FringeFF regs_257 ( // @[RegFile.scala 66:20:@128588.4]
    .clock(regs_257_clock),
    .reset(regs_257_reset),
    .io_in(regs_257_io_in),
    .io_reset(regs_257_io_reset),
    .io_out(regs_257_io_out),
    .io_enable(regs_257_io_enable)
  );
  FringeFF regs_258 ( // @[RegFile.scala 66:20:@128602.4]
    .clock(regs_258_clock),
    .reset(regs_258_reset),
    .io_in(regs_258_io_in),
    .io_reset(regs_258_io_reset),
    .io_out(regs_258_io_out),
    .io_enable(regs_258_io_enable)
  );
  FringeFF regs_259 ( // @[RegFile.scala 66:20:@128616.4]
    .clock(regs_259_clock),
    .reset(regs_259_reset),
    .io_in(regs_259_io_in),
    .io_reset(regs_259_io_reset),
    .io_out(regs_259_io_out),
    .io_enable(regs_259_io_enable)
  );
  FringeFF regs_260 ( // @[RegFile.scala 66:20:@128630.4]
    .clock(regs_260_clock),
    .reset(regs_260_reset),
    .io_in(regs_260_io_in),
    .io_reset(regs_260_io_reset),
    .io_out(regs_260_io_out),
    .io_enable(regs_260_io_enable)
  );
  FringeFF regs_261 ( // @[RegFile.scala 66:20:@128644.4]
    .clock(regs_261_clock),
    .reset(regs_261_reset),
    .io_in(regs_261_io_in),
    .io_reset(regs_261_io_reset),
    .io_out(regs_261_io_out),
    .io_enable(regs_261_io_enable)
  );
  FringeFF regs_262 ( // @[RegFile.scala 66:20:@128658.4]
    .clock(regs_262_clock),
    .reset(regs_262_reset),
    .io_in(regs_262_io_in),
    .io_reset(regs_262_io_reset),
    .io_out(regs_262_io_out),
    .io_enable(regs_262_io_enable)
  );
  FringeFF regs_263 ( // @[RegFile.scala 66:20:@128672.4]
    .clock(regs_263_clock),
    .reset(regs_263_reset),
    .io_in(regs_263_io_in),
    .io_reset(regs_263_io_reset),
    .io_out(regs_263_io_out),
    .io_enable(regs_263_io_enable)
  );
  FringeFF regs_264 ( // @[RegFile.scala 66:20:@128686.4]
    .clock(regs_264_clock),
    .reset(regs_264_reset),
    .io_in(regs_264_io_in),
    .io_reset(regs_264_io_reset),
    .io_out(regs_264_io_out),
    .io_enable(regs_264_io_enable)
  );
  FringeFF regs_265 ( // @[RegFile.scala 66:20:@128700.4]
    .clock(regs_265_clock),
    .reset(regs_265_reset),
    .io_in(regs_265_io_in),
    .io_reset(regs_265_io_reset),
    .io_out(regs_265_io_out),
    .io_enable(regs_265_io_enable)
  );
  FringeFF regs_266 ( // @[RegFile.scala 66:20:@128714.4]
    .clock(regs_266_clock),
    .reset(regs_266_reset),
    .io_in(regs_266_io_in),
    .io_reset(regs_266_io_reset),
    .io_out(regs_266_io_out),
    .io_enable(regs_266_io_enable)
  );
  FringeFF regs_267 ( // @[RegFile.scala 66:20:@128728.4]
    .clock(regs_267_clock),
    .reset(regs_267_reset),
    .io_in(regs_267_io_in),
    .io_reset(regs_267_io_reset),
    .io_out(regs_267_io_out),
    .io_enable(regs_267_io_enable)
  );
  FringeFF regs_268 ( // @[RegFile.scala 66:20:@128742.4]
    .clock(regs_268_clock),
    .reset(regs_268_reset),
    .io_in(regs_268_io_in),
    .io_reset(regs_268_io_reset),
    .io_out(regs_268_io_out),
    .io_enable(regs_268_io_enable)
  );
  FringeFF regs_269 ( // @[RegFile.scala 66:20:@128756.4]
    .clock(regs_269_clock),
    .reset(regs_269_reset),
    .io_in(regs_269_io_in),
    .io_reset(regs_269_io_reset),
    .io_out(regs_269_io_out),
    .io_enable(regs_269_io_enable)
  );
  FringeFF regs_270 ( // @[RegFile.scala 66:20:@128770.4]
    .clock(regs_270_clock),
    .reset(regs_270_reset),
    .io_in(regs_270_io_in),
    .io_reset(regs_270_io_reset),
    .io_out(regs_270_io_out),
    .io_enable(regs_270_io_enable)
  );
  FringeFF regs_271 ( // @[RegFile.scala 66:20:@128784.4]
    .clock(regs_271_clock),
    .reset(regs_271_reset),
    .io_in(regs_271_io_in),
    .io_reset(regs_271_io_reset),
    .io_out(regs_271_io_out),
    .io_enable(regs_271_io_enable)
  );
  FringeFF regs_272 ( // @[RegFile.scala 66:20:@128798.4]
    .clock(regs_272_clock),
    .reset(regs_272_reset),
    .io_in(regs_272_io_in),
    .io_reset(regs_272_io_reset),
    .io_out(regs_272_io_out),
    .io_enable(regs_272_io_enable)
  );
  FringeFF regs_273 ( // @[RegFile.scala 66:20:@128812.4]
    .clock(regs_273_clock),
    .reset(regs_273_reset),
    .io_in(regs_273_io_in),
    .io_reset(regs_273_io_reset),
    .io_out(regs_273_io_out),
    .io_enable(regs_273_io_enable)
  );
  FringeFF regs_274 ( // @[RegFile.scala 66:20:@128826.4]
    .clock(regs_274_clock),
    .reset(regs_274_reset),
    .io_in(regs_274_io_in),
    .io_reset(regs_274_io_reset),
    .io_out(regs_274_io_out),
    .io_enable(regs_274_io_enable)
  );
  FringeFF regs_275 ( // @[RegFile.scala 66:20:@128840.4]
    .clock(regs_275_clock),
    .reset(regs_275_reset),
    .io_in(regs_275_io_in),
    .io_reset(regs_275_io_reset),
    .io_out(regs_275_io_out),
    .io_enable(regs_275_io_enable)
  );
  FringeFF regs_276 ( // @[RegFile.scala 66:20:@128854.4]
    .clock(regs_276_clock),
    .reset(regs_276_reset),
    .io_in(regs_276_io_in),
    .io_reset(regs_276_io_reset),
    .io_out(regs_276_io_out),
    .io_enable(regs_276_io_enable)
  );
  FringeFF regs_277 ( // @[RegFile.scala 66:20:@128868.4]
    .clock(regs_277_clock),
    .reset(regs_277_reset),
    .io_in(regs_277_io_in),
    .io_reset(regs_277_io_reset),
    .io_out(regs_277_io_out),
    .io_enable(regs_277_io_enable)
  );
  FringeFF regs_278 ( // @[RegFile.scala 66:20:@128882.4]
    .clock(regs_278_clock),
    .reset(regs_278_reset),
    .io_in(regs_278_io_in),
    .io_reset(regs_278_io_reset),
    .io_out(regs_278_io_out),
    .io_enable(regs_278_io_enable)
  );
  FringeFF regs_279 ( // @[RegFile.scala 66:20:@128896.4]
    .clock(regs_279_clock),
    .reset(regs_279_reset),
    .io_in(regs_279_io_in),
    .io_reset(regs_279_io_reset),
    .io_out(regs_279_io_out),
    .io_enable(regs_279_io_enable)
  );
  FringeFF regs_280 ( // @[RegFile.scala 66:20:@128910.4]
    .clock(regs_280_clock),
    .reset(regs_280_reset),
    .io_in(regs_280_io_in),
    .io_reset(regs_280_io_reset),
    .io_out(regs_280_io_out),
    .io_enable(regs_280_io_enable)
  );
  FringeFF regs_281 ( // @[RegFile.scala 66:20:@128924.4]
    .clock(regs_281_clock),
    .reset(regs_281_reset),
    .io_in(regs_281_io_in),
    .io_reset(regs_281_io_reset),
    .io_out(regs_281_io_out),
    .io_enable(regs_281_io_enable)
  );
  FringeFF regs_282 ( // @[RegFile.scala 66:20:@128938.4]
    .clock(regs_282_clock),
    .reset(regs_282_reset),
    .io_in(regs_282_io_in),
    .io_reset(regs_282_io_reset),
    .io_out(regs_282_io_out),
    .io_enable(regs_282_io_enable)
  );
  FringeFF regs_283 ( // @[RegFile.scala 66:20:@128952.4]
    .clock(regs_283_clock),
    .reset(regs_283_reset),
    .io_in(regs_283_io_in),
    .io_reset(regs_283_io_reset),
    .io_out(regs_283_io_out),
    .io_enable(regs_283_io_enable)
  );
  FringeFF regs_284 ( // @[RegFile.scala 66:20:@128966.4]
    .clock(regs_284_clock),
    .reset(regs_284_reset),
    .io_in(regs_284_io_in),
    .io_reset(regs_284_io_reset),
    .io_out(regs_284_io_out),
    .io_enable(regs_284_io_enable)
  );
  FringeFF regs_285 ( // @[RegFile.scala 66:20:@128980.4]
    .clock(regs_285_clock),
    .reset(regs_285_reset),
    .io_in(regs_285_io_in),
    .io_reset(regs_285_io_reset),
    .io_out(regs_285_io_out),
    .io_enable(regs_285_io_enable)
  );
  FringeFF regs_286 ( // @[RegFile.scala 66:20:@128994.4]
    .clock(regs_286_clock),
    .reset(regs_286_reset),
    .io_in(regs_286_io_in),
    .io_reset(regs_286_io_reset),
    .io_out(regs_286_io_out),
    .io_enable(regs_286_io_enable)
  );
  FringeFF regs_287 ( // @[RegFile.scala 66:20:@129008.4]
    .clock(regs_287_clock),
    .reset(regs_287_reset),
    .io_in(regs_287_io_in),
    .io_reset(regs_287_io_reset),
    .io_out(regs_287_io_out),
    .io_enable(regs_287_io_enable)
  );
  FringeFF regs_288 ( // @[RegFile.scala 66:20:@129022.4]
    .clock(regs_288_clock),
    .reset(regs_288_reset),
    .io_in(regs_288_io_in),
    .io_reset(regs_288_io_reset),
    .io_out(regs_288_io_out),
    .io_enable(regs_288_io_enable)
  );
  FringeFF regs_289 ( // @[RegFile.scala 66:20:@129036.4]
    .clock(regs_289_clock),
    .reset(regs_289_reset),
    .io_in(regs_289_io_in),
    .io_reset(regs_289_io_reset),
    .io_out(regs_289_io_out),
    .io_enable(regs_289_io_enable)
  );
  FringeFF regs_290 ( // @[RegFile.scala 66:20:@129050.4]
    .clock(regs_290_clock),
    .reset(regs_290_reset),
    .io_in(regs_290_io_in),
    .io_reset(regs_290_io_reset),
    .io_out(regs_290_io_out),
    .io_enable(regs_290_io_enable)
  );
  FringeFF regs_291 ( // @[RegFile.scala 66:20:@129064.4]
    .clock(regs_291_clock),
    .reset(regs_291_reset),
    .io_in(regs_291_io_in),
    .io_reset(regs_291_io_reset),
    .io_out(regs_291_io_out),
    .io_enable(regs_291_io_enable)
  );
  FringeFF regs_292 ( // @[RegFile.scala 66:20:@129078.4]
    .clock(regs_292_clock),
    .reset(regs_292_reset),
    .io_in(regs_292_io_in),
    .io_reset(regs_292_io_reset),
    .io_out(regs_292_io_out),
    .io_enable(regs_292_io_enable)
  );
  FringeFF regs_293 ( // @[RegFile.scala 66:20:@129092.4]
    .clock(regs_293_clock),
    .reset(regs_293_reset),
    .io_in(regs_293_io_in),
    .io_reset(regs_293_io_reset),
    .io_out(regs_293_io_out),
    .io_enable(regs_293_io_enable)
  );
  FringeFF regs_294 ( // @[RegFile.scala 66:20:@129106.4]
    .clock(regs_294_clock),
    .reset(regs_294_reset),
    .io_in(regs_294_io_in),
    .io_reset(regs_294_io_reset),
    .io_out(regs_294_io_out),
    .io_enable(regs_294_io_enable)
  );
  FringeFF regs_295 ( // @[RegFile.scala 66:20:@129120.4]
    .clock(regs_295_clock),
    .reset(regs_295_reset),
    .io_in(regs_295_io_in),
    .io_reset(regs_295_io_reset),
    .io_out(regs_295_io_out),
    .io_enable(regs_295_io_enable)
  );
  FringeFF regs_296 ( // @[RegFile.scala 66:20:@129134.4]
    .clock(regs_296_clock),
    .reset(regs_296_reset),
    .io_in(regs_296_io_in),
    .io_reset(regs_296_io_reset),
    .io_out(regs_296_io_out),
    .io_enable(regs_296_io_enable)
  );
  FringeFF regs_297 ( // @[RegFile.scala 66:20:@129148.4]
    .clock(regs_297_clock),
    .reset(regs_297_reset),
    .io_in(regs_297_io_in),
    .io_reset(regs_297_io_reset),
    .io_out(regs_297_io_out),
    .io_enable(regs_297_io_enable)
  );
  FringeFF regs_298 ( // @[RegFile.scala 66:20:@129162.4]
    .clock(regs_298_clock),
    .reset(regs_298_reset),
    .io_in(regs_298_io_in),
    .io_reset(regs_298_io_reset),
    .io_out(regs_298_io_out),
    .io_enable(regs_298_io_enable)
  );
  FringeFF regs_299 ( // @[RegFile.scala 66:20:@129176.4]
    .clock(regs_299_clock),
    .reset(regs_299_reset),
    .io_in(regs_299_io_in),
    .io_reset(regs_299_io_reset),
    .io_out(regs_299_io_out),
    .io_enable(regs_299_io_enable)
  );
  FringeFF regs_300 ( // @[RegFile.scala 66:20:@129190.4]
    .clock(regs_300_clock),
    .reset(regs_300_reset),
    .io_in(regs_300_io_in),
    .io_reset(regs_300_io_reset),
    .io_out(regs_300_io_out),
    .io_enable(regs_300_io_enable)
  );
  FringeFF regs_301 ( // @[RegFile.scala 66:20:@129204.4]
    .clock(regs_301_clock),
    .reset(regs_301_reset),
    .io_in(regs_301_io_in),
    .io_reset(regs_301_io_reset),
    .io_out(regs_301_io_out),
    .io_enable(regs_301_io_enable)
  );
  FringeFF regs_302 ( // @[RegFile.scala 66:20:@129218.4]
    .clock(regs_302_clock),
    .reset(regs_302_reset),
    .io_in(regs_302_io_in),
    .io_reset(regs_302_io_reset),
    .io_out(regs_302_io_out),
    .io_enable(regs_302_io_enable)
  );
  FringeFF regs_303 ( // @[RegFile.scala 66:20:@129232.4]
    .clock(regs_303_clock),
    .reset(regs_303_reset),
    .io_in(regs_303_io_in),
    .io_reset(regs_303_io_reset),
    .io_out(regs_303_io_out),
    .io_enable(regs_303_io_enable)
  );
  FringeFF regs_304 ( // @[RegFile.scala 66:20:@129246.4]
    .clock(regs_304_clock),
    .reset(regs_304_reset),
    .io_in(regs_304_io_in),
    .io_reset(regs_304_io_reset),
    .io_out(regs_304_io_out),
    .io_enable(regs_304_io_enable)
  );
  FringeFF regs_305 ( // @[RegFile.scala 66:20:@129260.4]
    .clock(regs_305_clock),
    .reset(regs_305_reset),
    .io_in(regs_305_io_in),
    .io_reset(regs_305_io_reset),
    .io_out(regs_305_io_out),
    .io_enable(regs_305_io_enable)
  );
  FringeFF regs_306 ( // @[RegFile.scala 66:20:@129274.4]
    .clock(regs_306_clock),
    .reset(regs_306_reset),
    .io_in(regs_306_io_in),
    .io_reset(regs_306_io_reset),
    .io_out(regs_306_io_out),
    .io_enable(regs_306_io_enable)
  );
  FringeFF regs_307 ( // @[RegFile.scala 66:20:@129288.4]
    .clock(regs_307_clock),
    .reset(regs_307_reset),
    .io_in(regs_307_io_in),
    .io_reset(regs_307_io_reset),
    .io_out(regs_307_io_out),
    .io_enable(regs_307_io_enable)
  );
  FringeFF regs_308 ( // @[RegFile.scala 66:20:@129302.4]
    .clock(regs_308_clock),
    .reset(regs_308_reset),
    .io_in(regs_308_io_in),
    .io_reset(regs_308_io_reset),
    .io_out(regs_308_io_out),
    .io_enable(regs_308_io_enable)
  );
  FringeFF regs_309 ( // @[RegFile.scala 66:20:@129316.4]
    .clock(regs_309_clock),
    .reset(regs_309_reset),
    .io_in(regs_309_io_in),
    .io_reset(regs_309_io_reset),
    .io_out(regs_309_io_out),
    .io_enable(regs_309_io_enable)
  );
  FringeFF regs_310 ( // @[RegFile.scala 66:20:@129330.4]
    .clock(regs_310_clock),
    .reset(regs_310_reset),
    .io_in(regs_310_io_in),
    .io_reset(regs_310_io_reset),
    .io_out(regs_310_io_out),
    .io_enable(regs_310_io_enable)
  );
  FringeFF regs_311 ( // @[RegFile.scala 66:20:@129344.4]
    .clock(regs_311_clock),
    .reset(regs_311_reset),
    .io_in(regs_311_io_in),
    .io_reset(regs_311_io_reset),
    .io_out(regs_311_io_out),
    .io_enable(regs_311_io_enable)
  );
  FringeFF regs_312 ( // @[RegFile.scala 66:20:@129358.4]
    .clock(regs_312_clock),
    .reset(regs_312_reset),
    .io_in(regs_312_io_in),
    .io_reset(regs_312_io_reset),
    .io_out(regs_312_io_out),
    .io_enable(regs_312_io_enable)
  );
  FringeFF regs_313 ( // @[RegFile.scala 66:20:@129372.4]
    .clock(regs_313_clock),
    .reset(regs_313_reset),
    .io_in(regs_313_io_in),
    .io_reset(regs_313_io_reset),
    .io_out(regs_313_io_out),
    .io_enable(regs_313_io_enable)
  );
  FringeFF regs_314 ( // @[RegFile.scala 66:20:@129386.4]
    .clock(regs_314_clock),
    .reset(regs_314_reset),
    .io_in(regs_314_io_in),
    .io_reset(regs_314_io_reset),
    .io_out(regs_314_io_out),
    .io_enable(regs_314_io_enable)
  );
  FringeFF regs_315 ( // @[RegFile.scala 66:20:@129400.4]
    .clock(regs_315_clock),
    .reset(regs_315_reset),
    .io_in(regs_315_io_in),
    .io_reset(regs_315_io_reset),
    .io_out(regs_315_io_out),
    .io_enable(regs_315_io_enable)
  );
  FringeFF regs_316 ( // @[RegFile.scala 66:20:@129414.4]
    .clock(regs_316_clock),
    .reset(regs_316_reset),
    .io_in(regs_316_io_in),
    .io_reset(regs_316_io_reset),
    .io_out(regs_316_io_out),
    .io_enable(regs_316_io_enable)
  );
  FringeFF regs_317 ( // @[RegFile.scala 66:20:@129428.4]
    .clock(regs_317_clock),
    .reset(regs_317_reset),
    .io_in(regs_317_io_in),
    .io_reset(regs_317_io_reset),
    .io_out(regs_317_io_out),
    .io_enable(regs_317_io_enable)
  );
  FringeFF regs_318 ( // @[RegFile.scala 66:20:@129442.4]
    .clock(regs_318_clock),
    .reset(regs_318_reset),
    .io_in(regs_318_io_in),
    .io_reset(regs_318_io_reset),
    .io_out(regs_318_io_out),
    .io_enable(regs_318_io_enable)
  );
  FringeFF regs_319 ( // @[RegFile.scala 66:20:@129456.4]
    .clock(regs_319_clock),
    .reset(regs_319_reset),
    .io_in(regs_319_io_in),
    .io_reset(regs_319_io_reset),
    .io_out(regs_319_io_out),
    .io_enable(regs_319_io_enable)
  );
  FringeFF regs_320 ( // @[RegFile.scala 66:20:@129470.4]
    .clock(regs_320_clock),
    .reset(regs_320_reset),
    .io_in(regs_320_io_in),
    .io_reset(regs_320_io_reset),
    .io_out(regs_320_io_out),
    .io_enable(regs_320_io_enable)
  );
  FringeFF regs_321 ( // @[RegFile.scala 66:20:@129484.4]
    .clock(regs_321_clock),
    .reset(regs_321_reset),
    .io_in(regs_321_io_in),
    .io_reset(regs_321_io_reset),
    .io_out(regs_321_io_out),
    .io_enable(regs_321_io_enable)
  );
  FringeFF regs_322 ( // @[RegFile.scala 66:20:@129498.4]
    .clock(regs_322_clock),
    .reset(regs_322_reset),
    .io_in(regs_322_io_in),
    .io_reset(regs_322_io_reset),
    .io_out(regs_322_io_out),
    .io_enable(regs_322_io_enable)
  );
  FringeFF regs_323 ( // @[RegFile.scala 66:20:@129512.4]
    .clock(regs_323_clock),
    .reset(regs_323_reset),
    .io_in(regs_323_io_in),
    .io_reset(regs_323_io_reset),
    .io_out(regs_323_io_out),
    .io_enable(regs_323_io_enable)
  );
  FringeFF regs_324 ( // @[RegFile.scala 66:20:@129526.4]
    .clock(regs_324_clock),
    .reset(regs_324_reset),
    .io_in(regs_324_io_in),
    .io_reset(regs_324_io_reset),
    .io_out(regs_324_io_out),
    .io_enable(regs_324_io_enable)
  );
  FringeFF regs_325 ( // @[RegFile.scala 66:20:@129540.4]
    .clock(regs_325_clock),
    .reset(regs_325_reset),
    .io_in(regs_325_io_in),
    .io_reset(regs_325_io_reset),
    .io_out(regs_325_io_out),
    .io_enable(regs_325_io_enable)
  );
  FringeFF regs_326 ( // @[RegFile.scala 66:20:@129554.4]
    .clock(regs_326_clock),
    .reset(regs_326_reset),
    .io_in(regs_326_io_in),
    .io_reset(regs_326_io_reset),
    .io_out(regs_326_io_out),
    .io_enable(regs_326_io_enable)
  );
  FringeFF regs_327 ( // @[RegFile.scala 66:20:@129568.4]
    .clock(regs_327_clock),
    .reset(regs_327_reset),
    .io_in(regs_327_io_in),
    .io_reset(regs_327_io_reset),
    .io_out(regs_327_io_out),
    .io_enable(regs_327_io_enable)
  );
  FringeFF regs_328 ( // @[RegFile.scala 66:20:@129582.4]
    .clock(regs_328_clock),
    .reset(regs_328_reset),
    .io_in(regs_328_io_in),
    .io_reset(regs_328_io_reset),
    .io_out(regs_328_io_out),
    .io_enable(regs_328_io_enable)
  );
  FringeFF regs_329 ( // @[RegFile.scala 66:20:@129596.4]
    .clock(regs_329_clock),
    .reset(regs_329_reset),
    .io_in(regs_329_io_in),
    .io_reset(regs_329_io_reset),
    .io_out(regs_329_io_out),
    .io_enable(regs_329_io_enable)
  );
  FringeFF regs_330 ( // @[RegFile.scala 66:20:@129610.4]
    .clock(regs_330_clock),
    .reset(regs_330_reset),
    .io_in(regs_330_io_in),
    .io_reset(regs_330_io_reset),
    .io_out(regs_330_io_out),
    .io_enable(regs_330_io_enable)
  );
  FringeFF regs_331 ( // @[RegFile.scala 66:20:@129624.4]
    .clock(regs_331_clock),
    .reset(regs_331_reset),
    .io_in(regs_331_io_in),
    .io_reset(regs_331_io_reset),
    .io_out(regs_331_io_out),
    .io_enable(regs_331_io_enable)
  );
  FringeFF regs_332 ( // @[RegFile.scala 66:20:@129638.4]
    .clock(regs_332_clock),
    .reset(regs_332_reset),
    .io_in(regs_332_io_in),
    .io_reset(regs_332_io_reset),
    .io_out(regs_332_io_out),
    .io_enable(regs_332_io_enable)
  );
  FringeFF regs_333 ( // @[RegFile.scala 66:20:@129652.4]
    .clock(regs_333_clock),
    .reset(regs_333_reset),
    .io_in(regs_333_io_in),
    .io_reset(regs_333_io_reset),
    .io_out(regs_333_io_out),
    .io_enable(regs_333_io_enable)
  );
  FringeFF regs_334 ( // @[RegFile.scala 66:20:@129666.4]
    .clock(regs_334_clock),
    .reset(regs_334_reset),
    .io_in(regs_334_io_in),
    .io_reset(regs_334_io_reset),
    .io_out(regs_334_io_out),
    .io_enable(regs_334_io_enable)
  );
  FringeFF regs_335 ( // @[RegFile.scala 66:20:@129680.4]
    .clock(regs_335_clock),
    .reset(regs_335_reset),
    .io_in(regs_335_io_in),
    .io_reset(regs_335_io_reset),
    .io_out(regs_335_io_out),
    .io_enable(regs_335_io_enable)
  );
  FringeFF regs_336 ( // @[RegFile.scala 66:20:@129694.4]
    .clock(regs_336_clock),
    .reset(regs_336_reset),
    .io_in(regs_336_io_in),
    .io_reset(regs_336_io_reset),
    .io_out(regs_336_io_out),
    .io_enable(regs_336_io_enable)
  );
  FringeFF regs_337 ( // @[RegFile.scala 66:20:@129708.4]
    .clock(regs_337_clock),
    .reset(regs_337_reset),
    .io_in(regs_337_io_in),
    .io_reset(regs_337_io_reset),
    .io_out(regs_337_io_out),
    .io_enable(regs_337_io_enable)
  );
  FringeFF regs_338 ( // @[RegFile.scala 66:20:@129722.4]
    .clock(regs_338_clock),
    .reset(regs_338_reset),
    .io_in(regs_338_io_in),
    .io_reset(regs_338_io_reset),
    .io_out(regs_338_io_out),
    .io_enable(regs_338_io_enable)
  );
  FringeFF regs_339 ( // @[RegFile.scala 66:20:@129736.4]
    .clock(regs_339_clock),
    .reset(regs_339_reset),
    .io_in(regs_339_io_in),
    .io_reset(regs_339_io_reset),
    .io_out(regs_339_io_out),
    .io_enable(regs_339_io_enable)
  );
  FringeFF regs_340 ( // @[RegFile.scala 66:20:@129750.4]
    .clock(regs_340_clock),
    .reset(regs_340_reset),
    .io_in(regs_340_io_in),
    .io_reset(regs_340_io_reset),
    .io_out(regs_340_io_out),
    .io_enable(regs_340_io_enable)
  );
  FringeFF regs_341 ( // @[RegFile.scala 66:20:@129764.4]
    .clock(regs_341_clock),
    .reset(regs_341_reset),
    .io_in(regs_341_io_in),
    .io_reset(regs_341_io_reset),
    .io_out(regs_341_io_out),
    .io_enable(regs_341_io_enable)
  );
  FringeFF regs_342 ( // @[RegFile.scala 66:20:@129778.4]
    .clock(regs_342_clock),
    .reset(regs_342_reset),
    .io_in(regs_342_io_in),
    .io_reset(regs_342_io_reset),
    .io_out(regs_342_io_out),
    .io_enable(regs_342_io_enable)
  );
  FringeFF regs_343 ( // @[RegFile.scala 66:20:@129792.4]
    .clock(regs_343_clock),
    .reset(regs_343_reset),
    .io_in(regs_343_io_in),
    .io_reset(regs_343_io_reset),
    .io_out(regs_343_io_out),
    .io_enable(regs_343_io_enable)
  );
  FringeFF regs_344 ( // @[RegFile.scala 66:20:@129806.4]
    .clock(regs_344_clock),
    .reset(regs_344_reset),
    .io_in(regs_344_io_in),
    .io_reset(regs_344_io_reset),
    .io_out(regs_344_io_out),
    .io_enable(regs_344_io_enable)
  );
  FringeFF regs_345 ( // @[RegFile.scala 66:20:@129820.4]
    .clock(regs_345_clock),
    .reset(regs_345_reset),
    .io_in(regs_345_io_in),
    .io_reset(regs_345_io_reset),
    .io_out(regs_345_io_out),
    .io_enable(regs_345_io_enable)
  );
  FringeFF regs_346 ( // @[RegFile.scala 66:20:@129834.4]
    .clock(regs_346_clock),
    .reset(regs_346_reset),
    .io_in(regs_346_io_in),
    .io_reset(regs_346_io_reset),
    .io_out(regs_346_io_out),
    .io_enable(regs_346_io_enable)
  );
  FringeFF regs_347 ( // @[RegFile.scala 66:20:@129848.4]
    .clock(regs_347_clock),
    .reset(regs_347_reset),
    .io_in(regs_347_io_in),
    .io_reset(regs_347_io_reset),
    .io_out(regs_347_io_out),
    .io_enable(regs_347_io_enable)
  );
  FringeFF regs_348 ( // @[RegFile.scala 66:20:@129862.4]
    .clock(regs_348_clock),
    .reset(regs_348_reset),
    .io_in(regs_348_io_in),
    .io_reset(regs_348_io_reset),
    .io_out(regs_348_io_out),
    .io_enable(regs_348_io_enable)
  );
  FringeFF regs_349 ( // @[RegFile.scala 66:20:@129876.4]
    .clock(regs_349_clock),
    .reset(regs_349_reset),
    .io_in(regs_349_io_in),
    .io_reset(regs_349_io_reset),
    .io_out(regs_349_io_out),
    .io_enable(regs_349_io_enable)
  );
  FringeFF regs_350 ( // @[RegFile.scala 66:20:@129890.4]
    .clock(regs_350_clock),
    .reset(regs_350_reset),
    .io_in(regs_350_io_in),
    .io_reset(regs_350_io_reset),
    .io_out(regs_350_io_out),
    .io_enable(regs_350_io_enable)
  );
  FringeFF regs_351 ( // @[RegFile.scala 66:20:@129904.4]
    .clock(regs_351_clock),
    .reset(regs_351_reset),
    .io_in(regs_351_io_in),
    .io_reset(regs_351_io_reset),
    .io_out(regs_351_io_out),
    .io_enable(regs_351_io_enable)
  );
  FringeFF regs_352 ( // @[RegFile.scala 66:20:@129918.4]
    .clock(regs_352_clock),
    .reset(regs_352_reset),
    .io_in(regs_352_io_in),
    .io_reset(regs_352_io_reset),
    .io_out(regs_352_io_out),
    .io_enable(regs_352_io_enable)
  );
  FringeFF regs_353 ( // @[RegFile.scala 66:20:@129932.4]
    .clock(regs_353_clock),
    .reset(regs_353_reset),
    .io_in(regs_353_io_in),
    .io_reset(regs_353_io_reset),
    .io_out(regs_353_io_out),
    .io_enable(regs_353_io_enable)
  );
  FringeFF regs_354 ( // @[RegFile.scala 66:20:@129946.4]
    .clock(regs_354_clock),
    .reset(regs_354_reset),
    .io_in(regs_354_io_in),
    .io_reset(regs_354_io_reset),
    .io_out(regs_354_io_out),
    .io_enable(regs_354_io_enable)
  );
  FringeFF regs_355 ( // @[RegFile.scala 66:20:@129960.4]
    .clock(regs_355_clock),
    .reset(regs_355_reset),
    .io_in(regs_355_io_in),
    .io_reset(regs_355_io_reset),
    .io_out(regs_355_io_out),
    .io_enable(regs_355_io_enable)
  );
  FringeFF regs_356 ( // @[RegFile.scala 66:20:@129974.4]
    .clock(regs_356_clock),
    .reset(regs_356_reset),
    .io_in(regs_356_io_in),
    .io_reset(regs_356_io_reset),
    .io_out(regs_356_io_out),
    .io_enable(regs_356_io_enable)
  );
  FringeFF regs_357 ( // @[RegFile.scala 66:20:@129988.4]
    .clock(regs_357_clock),
    .reset(regs_357_reset),
    .io_in(regs_357_io_in),
    .io_reset(regs_357_io_reset),
    .io_out(regs_357_io_out),
    .io_enable(regs_357_io_enable)
  );
  FringeFF regs_358 ( // @[RegFile.scala 66:20:@130002.4]
    .clock(regs_358_clock),
    .reset(regs_358_reset),
    .io_in(regs_358_io_in),
    .io_reset(regs_358_io_reset),
    .io_out(regs_358_io_out),
    .io_enable(regs_358_io_enable)
  );
  FringeFF regs_359 ( // @[RegFile.scala 66:20:@130016.4]
    .clock(regs_359_clock),
    .reset(regs_359_reset),
    .io_in(regs_359_io_in),
    .io_reset(regs_359_io_reset),
    .io_out(regs_359_io_out),
    .io_enable(regs_359_io_enable)
  );
  FringeFF regs_360 ( // @[RegFile.scala 66:20:@130030.4]
    .clock(regs_360_clock),
    .reset(regs_360_reset),
    .io_in(regs_360_io_in),
    .io_reset(regs_360_io_reset),
    .io_out(regs_360_io_out),
    .io_enable(regs_360_io_enable)
  );
  FringeFF regs_361 ( // @[RegFile.scala 66:20:@130044.4]
    .clock(regs_361_clock),
    .reset(regs_361_reset),
    .io_in(regs_361_io_in),
    .io_reset(regs_361_io_reset),
    .io_out(regs_361_io_out),
    .io_enable(regs_361_io_enable)
  );
  FringeFF regs_362 ( // @[RegFile.scala 66:20:@130058.4]
    .clock(regs_362_clock),
    .reset(regs_362_reset),
    .io_in(regs_362_io_in),
    .io_reset(regs_362_io_reset),
    .io_out(regs_362_io_out),
    .io_enable(regs_362_io_enable)
  );
  FringeFF regs_363 ( // @[RegFile.scala 66:20:@130072.4]
    .clock(regs_363_clock),
    .reset(regs_363_reset),
    .io_in(regs_363_io_in),
    .io_reset(regs_363_io_reset),
    .io_out(regs_363_io_out),
    .io_enable(regs_363_io_enable)
  );
  FringeFF regs_364 ( // @[RegFile.scala 66:20:@130086.4]
    .clock(regs_364_clock),
    .reset(regs_364_reset),
    .io_in(regs_364_io_in),
    .io_reset(regs_364_io_reset),
    .io_out(regs_364_io_out),
    .io_enable(regs_364_io_enable)
  );
  FringeFF regs_365 ( // @[RegFile.scala 66:20:@130100.4]
    .clock(regs_365_clock),
    .reset(regs_365_reset),
    .io_in(regs_365_io_in),
    .io_reset(regs_365_io_reset),
    .io_out(regs_365_io_out),
    .io_enable(regs_365_io_enable)
  );
  FringeFF regs_366 ( // @[RegFile.scala 66:20:@130114.4]
    .clock(regs_366_clock),
    .reset(regs_366_reset),
    .io_in(regs_366_io_in),
    .io_reset(regs_366_io_reset),
    .io_out(regs_366_io_out),
    .io_enable(regs_366_io_enable)
  );
  FringeFF regs_367 ( // @[RegFile.scala 66:20:@130128.4]
    .clock(regs_367_clock),
    .reset(regs_367_reset),
    .io_in(regs_367_io_in),
    .io_reset(regs_367_io_reset),
    .io_out(regs_367_io_out),
    .io_enable(regs_367_io_enable)
  );
  FringeFF regs_368 ( // @[RegFile.scala 66:20:@130142.4]
    .clock(regs_368_clock),
    .reset(regs_368_reset),
    .io_in(regs_368_io_in),
    .io_reset(regs_368_io_reset),
    .io_out(regs_368_io_out),
    .io_enable(regs_368_io_enable)
  );
  FringeFF regs_369 ( // @[RegFile.scala 66:20:@130156.4]
    .clock(regs_369_clock),
    .reset(regs_369_reset),
    .io_in(regs_369_io_in),
    .io_reset(regs_369_io_reset),
    .io_out(regs_369_io_out),
    .io_enable(regs_369_io_enable)
  );
  FringeFF regs_370 ( // @[RegFile.scala 66:20:@130170.4]
    .clock(regs_370_clock),
    .reset(regs_370_reset),
    .io_in(regs_370_io_in),
    .io_reset(regs_370_io_reset),
    .io_out(regs_370_io_out),
    .io_enable(regs_370_io_enable)
  );
  FringeFF regs_371 ( // @[RegFile.scala 66:20:@130184.4]
    .clock(regs_371_clock),
    .reset(regs_371_reset),
    .io_in(regs_371_io_in),
    .io_reset(regs_371_io_reset),
    .io_out(regs_371_io_out),
    .io_enable(regs_371_io_enable)
  );
  FringeFF regs_372 ( // @[RegFile.scala 66:20:@130198.4]
    .clock(regs_372_clock),
    .reset(regs_372_reset),
    .io_in(regs_372_io_in),
    .io_reset(regs_372_io_reset),
    .io_out(regs_372_io_out),
    .io_enable(regs_372_io_enable)
  );
  FringeFF regs_373 ( // @[RegFile.scala 66:20:@130212.4]
    .clock(regs_373_clock),
    .reset(regs_373_reset),
    .io_in(regs_373_io_in),
    .io_reset(regs_373_io_reset),
    .io_out(regs_373_io_out),
    .io_enable(regs_373_io_enable)
  );
  FringeFF regs_374 ( // @[RegFile.scala 66:20:@130226.4]
    .clock(regs_374_clock),
    .reset(regs_374_reset),
    .io_in(regs_374_io_in),
    .io_reset(regs_374_io_reset),
    .io_out(regs_374_io_out),
    .io_enable(regs_374_io_enable)
  );
  FringeFF regs_375 ( // @[RegFile.scala 66:20:@130240.4]
    .clock(regs_375_clock),
    .reset(regs_375_reset),
    .io_in(regs_375_io_in),
    .io_reset(regs_375_io_reset),
    .io_out(regs_375_io_out),
    .io_enable(regs_375_io_enable)
  );
  FringeFF regs_376 ( // @[RegFile.scala 66:20:@130254.4]
    .clock(regs_376_clock),
    .reset(regs_376_reset),
    .io_in(regs_376_io_in),
    .io_reset(regs_376_io_reset),
    .io_out(regs_376_io_out),
    .io_enable(regs_376_io_enable)
  );
  FringeFF regs_377 ( // @[RegFile.scala 66:20:@130268.4]
    .clock(regs_377_clock),
    .reset(regs_377_reset),
    .io_in(regs_377_io_in),
    .io_reset(regs_377_io_reset),
    .io_out(regs_377_io_out),
    .io_enable(regs_377_io_enable)
  );
  FringeFF regs_378 ( // @[RegFile.scala 66:20:@130282.4]
    .clock(regs_378_clock),
    .reset(regs_378_reset),
    .io_in(regs_378_io_in),
    .io_reset(regs_378_io_reset),
    .io_out(regs_378_io_out),
    .io_enable(regs_378_io_enable)
  );
  FringeFF regs_379 ( // @[RegFile.scala 66:20:@130296.4]
    .clock(regs_379_clock),
    .reset(regs_379_reset),
    .io_in(regs_379_io_in),
    .io_reset(regs_379_io_reset),
    .io_out(regs_379_io_out),
    .io_enable(regs_379_io_enable)
  );
  FringeFF regs_380 ( // @[RegFile.scala 66:20:@130310.4]
    .clock(regs_380_clock),
    .reset(regs_380_reset),
    .io_in(regs_380_io_in),
    .io_reset(regs_380_io_reset),
    .io_out(regs_380_io_out),
    .io_enable(regs_380_io_enable)
  );
  FringeFF regs_381 ( // @[RegFile.scala 66:20:@130324.4]
    .clock(regs_381_clock),
    .reset(regs_381_reset),
    .io_in(regs_381_io_in),
    .io_reset(regs_381_io_reset),
    .io_out(regs_381_io_out),
    .io_enable(regs_381_io_enable)
  );
  FringeFF regs_382 ( // @[RegFile.scala 66:20:@130338.4]
    .clock(regs_382_clock),
    .reset(regs_382_reset),
    .io_in(regs_382_io_in),
    .io_reset(regs_382_io_reset),
    .io_out(regs_382_io_out),
    .io_enable(regs_382_io_enable)
  );
  FringeFF regs_383 ( // @[RegFile.scala 66:20:@130352.4]
    .clock(regs_383_clock),
    .reset(regs_383_reset),
    .io_in(regs_383_io_in),
    .io_reset(regs_383_io_reset),
    .io_out(regs_383_io_out),
    .io_enable(regs_383_io_enable)
  );
  FringeFF regs_384 ( // @[RegFile.scala 66:20:@130366.4]
    .clock(regs_384_clock),
    .reset(regs_384_reset),
    .io_in(regs_384_io_in),
    .io_reset(regs_384_io_reset),
    .io_out(regs_384_io_out),
    .io_enable(regs_384_io_enable)
  );
  FringeFF regs_385 ( // @[RegFile.scala 66:20:@130380.4]
    .clock(regs_385_clock),
    .reset(regs_385_reset),
    .io_in(regs_385_io_in),
    .io_reset(regs_385_io_reset),
    .io_out(regs_385_io_out),
    .io_enable(regs_385_io_enable)
  );
  FringeFF regs_386 ( // @[RegFile.scala 66:20:@130394.4]
    .clock(regs_386_clock),
    .reset(regs_386_reset),
    .io_in(regs_386_io_in),
    .io_reset(regs_386_io_reset),
    .io_out(regs_386_io_out),
    .io_enable(regs_386_io_enable)
  );
  FringeFF regs_387 ( // @[RegFile.scala 66:20:@130408.4]
    .clock(regs_387_clock),
    .reset(regs_387_reset),
    .io_in(regs_387_io_in),
    .io_reset(regs_387_io_reset),
    .io_out(regs_387_io_out),
    .io_enable(regs_387_io_enable)
  );
  FringeFF regs_388 ( // @[RegFile.scala 66:20:@130422.4]
    .clock(regs_388_clock),
    .reset(regs_388_reset),
    .io_in(regs_388_io_in),
    .io_reset(regs_388_io_reset),
    .io_out(regs_388_io_out),
    .io_enable(regs_388_io_enable)
  );
  FringeFF regs_389 ( // @[RegFile.scala 66:20:@130436.4]
    .clock(regs_389_clock),
    .reset(regs_389_reset),
    .io_in(regs_389_io_in),
    .io_reset(regs_389_io_reset),
    .io_out(regs_389_io_out),
    .io_enable(regs_389_io_enable)
  );
  FringeFF regs_390 ( // @[RegFile.scala 66:20:@130450.4]
    .clock(regs_390_clock),
    .reset(regs_390_reset),
    .io_in(regs_390_io_in),
    .io_reset(regs_390_io_reset),
    .io_out(regs_390_io_out),
    .io_enable(regs_390_io_enable)
  );
  FringeFF regs_391 ( // @[RegFile.scala 66:20:@130464.4]
    .clock(regs_391_clock),
    .reset(regs_391_reset),
    .io_in(regs_391_io_in),
    .io_reset(regs_391_io_reset),
    .io_out(regs_391_io_out),
    .io_enable(regs_391_io_enable)
  );
  FringeFF regs_392 ( // @[RegFile.scala 66:20:@130478.4]
    .clock(regs_392_clock),
    .reset(regs_392_reset),
    .io_in(regs_392_io_in),
    .io_reset(regs_392_io_reset),
    .io_out(regs_392_io_out),
    .io_enable(regs_392_io_enable)
  );
  FringeFF regs_393 ( // @[RegFile.scala 66:20:@130492.4]
    .clock(regs_393_clock),
    .reset(regs_393_reset),
    .io_in(regs_393_io_in),
    .io_reset(regs_393_io_reset),
    .io_out(regs_393_io_out),
    .io_enable(regs_393_io_enable)
  );
  FringeFF regs_394 ( // @[RegFile.scala 66:20:@130506.4]
    .clock(regs_394_clock),
    .reset(regs_394_reset),
    .io_in(regs_394_io_in),
    .io_reset(regs_394_io_reset),
    .io_out(regs_394_io_out),
    .io_enable(regs_394_io_enable)
  );
  FringeFF regs_395 ( // @[RegFile.scala 66:20:@130520.4]
    .clock(regs_395_clock),
    .reset(regs_395_reset),
    .io_in(regs_395_io_in),
    .io_reset(regs_395_io_reset),
    .io_out(regs_395_io_out),
    .io_enable(regs_395_io_enable)
  );
  FringeFF regs_396 ( // @[RegFile.scala 66:20:@130534.4]
    .clock(regs_396_clock),
    .reset(regs_396_reset),
    .io_in(regs_396_io_in),
    .io_reset(regs_396_io_reset),
    .io_out(regs_396_io_out),
    .io_enable(regs_396_io_enable)
  );
  FringeFF regs_397 ( // @[RegFile.scala 66:20:@130548.4]
    .clock(regs_397_clock),
    .reset(regs_397_reset),
    .io_in(regs_397_io_in),
    .io_reset(regs_397_io_reset),
    .io_out(regs_397_io_out),
    .io_enable(regs_397_io_enable)
  );
  FringeFF regs_398 ( // @[RegFile.scala 66:20:@130562.4]
    .clock(regs_398_clock),
    .reset(regs_398_reset),
    .io_in(regs_398_io_in),
    .io_reset(regs_398_io_reset),
    .io_out(regs_398_io_out),
    .io_enable(regs_398_io_enable)
  );
  FringeFF regs_399 ( // @[RegFile.scala 66:20:@130576.4]
    .clock(regs_399_clock),
    .reset(regs_399_reset),
    .io_in(regs_399_io_in),
    .io_reset(regs_399_io_reset),
    .io_out(regs_399_io_out),
    .io_enable(regs_399_io_enable)
  );
  FringeFF regs_400 ( // @[RegFile.scala 66:20:@130590.4]
    .clock(regs_400_clock),
    .reset(regs_400_reset),
    .io_in(regs_400_io_in),
    .io_reset(regs_400_io_reset),
    .io_out(regs_400_io_out),
    .io_enable(regs_400_io_enable)
  );
  FringeFF regs_401 ( // @[RegFile.scala 66:20:@130604.4]
    .clock(regs_401_clock),
    .reset(regs_401_reset),
    .io_in(regs_401_io_in),
    .io_reset(regs_401_io_reset),
    .io_out(regs_401_io_out),
    .io_enable(regs_401_io_enable)
  );
  FringeFF regs_402 ( // @[RegFile.scala 66:20:@130618.4]
    .clock(regs_402_clock),
    .reset(regs_402_reset),
    .io_in(regs_402_io_in),
    .io_reset(regs_402_io_reset),
    .io_out(regs_402_io_out),
    .io_enable(regs_402_io_enable)
  );
  FringeFF regs_403 ( // @[RegFile.scala 66:20:@130632.4]
    .clock(regs_403_clock),
    .reset(regs_403_reset),
    .io_in(regs_403_io_in),
    .io_reset(regs_403_io_reset),
    .io_out(regs_403_io_out),
    .io_enable(regs_403_io_enable)
  );
  FringeFF regs_404 ( // @[RegFile.scala 66:20:@130646.4]
    .clock(regs_404_clock),
    .reset(regs_404_reset),
    .io_in(regs_404_io_in),
    .io_reset(regs_404_io_reset),
    .io_out(regs_404_io_out),
    .io_enable(regs_404_io_enable)
  );
  FringeFF regs_405 ( // @[RegFile.scala 66:20:@130660.4]
    .clock(regs_405_clock),
    .reset(regs_405_reset),
    .io_in(regs_405_io_in),
    .io_reset(regs_405_io_reset),
    .io_out(regs_405_io_out),
    .io_enable(regs_405_io_enable)
  );
  FringeFF regs_406 ( // @[RegFile.scala 66:20:@130674.4]
    .clock(regs_406_clock),
    .reset(regs_406_reset),
    .io_in(regs_406_io_in),
    .io_reset(regs_406_io_reset),
    .io_out(regs_406_io_out),
    .io_enable(regs_406_io_enable)
  );
  FringeFF regs_407 ( // @[RegFile.scala 66:20:@130688.4]
    .clock(regs_407_clock),
    .reset(regs_407_reset),
    .io_in(regs_407_io_in),
    .io_reset(regs_407_io_reset),
    .io_out(regs_407_io_out),
    .io_enable(regs_407_io_enable)
  );
  FringeFF regs_408 ( // @[RegFile.scala 66:20:@130702.4]
    .clock(regs_408_clock),
    .reset(regs_408_reset),
    .io_in(regs_408_io_in),
    .io_reset(regs_408_io_reset),
    .io_out(regs_408_io_out),
    .io_enable(regs_408_io_enable)
  );
  FringeFF regs_409 ( // @[RegFile.scala 66:20:@130716.4]
    .clock(regs_409_clock),
    .reset(regs_409_reset),
    .io_in(regs_409_io_in),
    .io_reset(regs_409_io_reset),
    .io_out(regs_409_io_out),
    .io_enable(regs_409_io_enable)
  );
  FringeFF regs_410 ( // @[RegFile.scala 66:20:@130730.4]
    .clock(regs_410_clock),
    .reset(regs_410_reset),
    .io_in(regs_410_io_in),
    .io_reset(regs_410_io_reset),
    .io_out(regs_410_io_out),
    .io_enable(regs_410_io_enable)
  );
  FringeFF regs_411 ( // @[RegFile.scala 66:20:@130744.4]
    .clock(regs_411_clock),
    .reset(regs_411_reset),
    .io_in(regs_411_io_in),
    .io_reset(regs_411_io_reset),
    .io_out(regs_411_io_out),
    .io_enable(regs_411_io_enable)
  );
  FringeFF regs_412 ( // @[RegFile.scala 66:20:@130758.4]
    .clock(regs_412_clock),
    .reset(regs_412_reset),
    .io_in(regs_412_io_in),
    .io_reset(regs_412_io_reset),
    .io_out(regs_412_io_out),
    .io_enable(regs_412_io_enable)
  );
  FringeFF regs_413 ( // @[RegFile.scala 66:20:@130772.4]
    .clock(regs_413_clock),
    .reset(regs_413_reset),
    .io_in(regs_413_io_in),
    .io_reset(regs_413_io_reset),
    .io_out(regs_413_io_out),
    .io_enable(regs_413_io_enable)
  );
  FringeFF regs_414 ( // @[RegFile.scala 66:20:@130786.4]
    .clock(regs_414_clock),
    .reset(regs_414_reset),
    .io_in(regs_414_io_in),
    .io_reset(regs_414_io_reset),
    .io_out(regs_414_io_out),
    .io_enable(regs_414_io_enable)
  );
  FringeFF regs_415 ( // @[RegFile.scala 66:20:@130800.4]
    .clock(regs_415_clock),
    .reset(regs_415_reset),
    .io_in(regs_415_io_in),
    .io_reset(regs_415_io_reset),
    .io_out(regs_415_io_out),
    .io_enable(regs_415_io_enable)
  );
  FringeFF regs_416 ( // @[RegFile.scala 66:20:@130814.4]
    .clock(regs_416_clock),
    .reset(regs_416_reset),
    .io_in(regs_416_io_in),
    .io_reset(regs_416_io_reset),
    .io_out(regs_416_io_out),
    .io_enable(regs_416_io_enable)
  );
  FringeFF regs_417 ( // @[RegFile.scala 66:20:@130828.4]
    .clock(regs_417_clock),
    .reset(regs_417_reset),
    .io_in(regs_417_io_in),
    .io_reset(regs_417_io_reset),
    .io_out(regs_417_io_out),
    .io_enable(regs_417_io_enable)
  );
  FringeFF regs_418 ( // @[RegFile.scala 66:20:@130842.4]
    .clock(regs_418_clock),
    .reset(regs_418_reset),
    .io_in(regs_418_io_in),
    .io_reset(regs_418_io_reset),
    .io_out(regs_418_io_out),
    .io_enable(regs_418_io_enable)
  );
  FringeFF regs_419 ( // @[RegFile.scala 66:20:@130856.4]
    .clock(regs_419_clock),
    .reset(regs_419_reset),
    .io_in(regs_419_io_in),
    .io_reset(regs_419_io_reset),
    .io_out(regs_419_io_out),
    .io_enable(regs_419_io_enable)
  );
  FringeFF regs_420 ( // @[RegFile.scala 66:20:@130870.4]
    .clock(regs_420_clock),
    .reset(regs_420_reset),
    .io_in(regs_420_io_in),
    .io_reset(regs_420_io_reset),
    .io_out(regs_420_io_out),
    .io_enable(regs_420_io_enable)
  );
  FringeFF regs_421 ( // @[RegFile.scala 66:20:@130884.4]
    .clock(regs_421_clock),
    .reset(regs_421_reset),
    .io_in(regs_421_io_in),
    .io_reset(regs_421_io_reset),
    .io_out(regs_421_io_out),
    .io_enable(regs_421_io_enable)
  );
  FringeFF regs_422 ( // @[RegFile.scala 66:20:@130898.4]
    .clock(regs_422_clock),
    .reset(regs_422_reset),
    .io_in(regs_422_io_in),
    .io_reset(regs_422_io_reset),
    .io_out(regs_422_io_out),
    .io_enable(regs_422_io_enable)
  );
  FringeFF regs_423 ( // @[RegFile.scala 66:20:@130912.4]
    .clock(regs_423_clock),
    .reset(regs_423_reset),
    .io_in(regs_423_io_in),
    .io_reset(regs_423_io_reset),
    .io_out(regs_423_io_out),
    .io_enable(regs_423_io_enable)
  );
  FringeFF regs_424 ( // @[RegFile.scala 66:20:@130926.4]
    .clock(regs_424_clock),
    .reset(regs_424_reset),
    .io_in(regs_424_io_in),
    .io_reset(regs_424_io_reset),
    .io_out(regs_424_io_out),
    .io_enable(regs_424_io_enable)
  );
  FringeFF regs_425 ( // @[RegFile.scala 66:20:@130940.4]
    .clock(regs_425_clock),
    .reset(regs_425_reset),
    .io_in(regs_425_io_in),
    .io_reset(regs_425_io_reset),
    .io_out(regs_425_io_out),
    .io_enable(regs_425_io_enable)
  );
  FringeFF regs_426 ( // @[RegFile.scala 66:20:@130954.4]
    .clock(regs_426_clock),
    .reset(regs_426_reset),
    .io_in(regs_426_io_in),
    .io_reset(regs_426_io_reset),
    .io_out(regs_426_io_out),
    .io_enable(regs_426_io_enable)
  );
  FringeFF regs_427 ( // @[RegFile.scala 66:20:@130968.4]
    .clock(regs_427_clock),
    .reset(regs_427_reset),
    .io_in(regs_427_io_in),
    .io_reset(regs_427_io_reset),
    .io_out(regs_427_io_out),
    .io_enable(regs_427_io_enable)
  );
  FringeFF regs_428 ( // @[RegFile.scala 66:20:@130982.4]
    .clock(regs_428_clock),
    .reset(regs_428_reset),
    .io_in(regs_428_io_in),
    .io_reset(regs_428_io_reset),
    .io_out(regs_428_io_out),
    .io_enable(regs_428_io_enable)
  );
  FringeFF regs_429 ( // @[RegFile.scala 66:20:@130996.4]
    .clock(regs_429_clock),
    .reset(regs_429_reset),
    .io_in(regs_429_io_in),
    .io_reset(regs_429_io_reset),
    .io_out(regs_429_io_out),
    .io_enable(regs_429_io_enable)
  );
  FringeFF regs_430 ( // @[RegFile.scala 66:20:@131010.4]
    .clock(regs_430_clock),
    .reset(regs_430_reset),
    .io_in(regs_430_io_in),
    .io_reset(regs_430_io_reset),
    .io_out(regs_430_io_out),
    .io_enable(regs_430_io_enable)
  );
  FringeFF regs_431 ( // @[RegFile.scala 66:20:@131024.4]
    .clock(regs_431_clock),
    .reset(regs_431_reset),
    .io_in(regs_431_io_in),
    .io_reset(regs_431_io_reset),
    .io_out(regs_431_io_out),
    .io_enable(regs_431_io_enable)
  );
  FringeFF regs_432 ( // @[RegFile.scala 66:20:@131038.4]
    .clock(regs_432_clock),
    .reset(regs_432_reset),
    .io_in(regs_432_io_in),
    .io_reset(regs_432_io_reset),
    .io_out(regs_432_io_out),
    .io_enable(regs_432_io_enable)
  );
  FringeFF regs_433 ( // @[RegFile.scala 66:20:@131052.4]
    .clock(regs_433_clock),
    .reset(regs_433_reset),
    .io_in(regs_433_io_in),
    .io_reset(regs_433_io_reset),
    .io_out(regs_433_io_out),
    .io_enable(regs_433_io_enable)
  );
  FringeFF regs_434 ( // @[RegFile.scala 66:20:@131066.4]
    .clock(regs_434_clock),
    .reset(regs_434_reset),
    .io_in(regs_434_io_in),
    .io_reset(regs_434_io_reset),
    .io_out(regs_434_io_out),
    .io_enable(regs_434_io_enable)
  );
  FringeFF regs_435 ( // @[RegFile.scala 66:20:@131080.4]
    .clock(regs_435_clock),
    .reset(regs_435_reset),
    .io_in(regs_435_io_in),
    .io_reset(regs_435_io_reset),
    .io_out(regs_435_io_out),
    .io_enable(regs_435_io_enable)
  );
  FringeFF regs_436 ( // @[RegFile.scala 66:20:@131094.4]
    .clock(regs_436_clock),
    .reset(regs_436_reset),
    .io_in(regs_436_io_in),
    .io_reset(regs_436_io_reset),
    .io_out(regs_436_io_out),
    .io_enable(regs_436_io_enable)
  );
  FringeFF regs_437 ( // @[RegFile.scala 66:20:@131108.4]
    .clock(regs_437_clock),
    .reset(regs_437_reset),
    .io_in(regs_437_io_in),
    .io_reset(regs_437_io_reset),
    .io_out(regs_437_io_out),
    .io_enable(regs_437_io_enable)
  );
  FringeFF regs_438 ( // @[RegFile.scala 66:20:@131122.4]
    .clock(regs_438_clock),
    .reset(regs_438_reset),
    .io_in(regs_438_io_in),
    .io_reset(regs_438_io_reset),
    .io_out(regs_438_io_out),
    .io_enable(regs_438_io_enable)
  );
  FringeFF regs_439 ( // @[RegFile.scala 66:20:@131136.4]
    .clock(regs_439_clock),
    .reset(regs_439_reset),
    .io_in(regs_439_io_in),
    .io_reset(regs_439_io_reset),
    .io_out(regs_439_io_out),
    .io_enable(regs_439_io_enable)
  );
  FringeFF regs_440 ( // @[RegFile.scala 66:20:@131150.4]
    .clock(regs_440_clock),
    .reset(regs_440_reset),
    .io_in(regs_440_io_in),
    .io_reset(regs_440_io_reset),
    .io_out(regs_440_io_out),
    .io_enable(regs_440_io_enable)
  );
  FringeFF regs_441 ( // @[RegFile.scala 66:20:@131164.4]
    .clock(regs_441_clock),
    .reset(regs_441_reset),
    .io_in(regs_441_io_in),
    .io_reset(regs_441_io_reset),
    .io_out(regs_441_io_out),
    .io_enable(regs_441_io_enable)
  );
  FringeFF regs_442 ( // @[RegFile.scala 66:20:@131178.4]
    .clock(regs_442_clock),
    .reset(regs_442_reset),
    .io_in(regs_442_io_in),
    .io_reset(regs_442_io_reset),
    .io_out(regs_442_io_out),
    .io_enable(regs_442_io_enable)
  );
  FringeFF regs_443 ( // @[RegFile.scala 66:20:@131192.4]
    .clock(regs_443_clock),
    .reset(regs_443_reset),
    .io_in(regs_443_io_in),
    .io_reset(regs_443_io_reset),
    .io_out(regs_443_io_out),
    .io_enable(regs_443_io_enable)
  );
  FringeFF regs_444 ( // @[RegFile.scala 66:20:@131206.4]
    .clock(regs_444_clock),
    .reset(regs_444_reset),
    .io_in(regs_444_io_in),
    .io_reset(regs_444_io_reset),
    .io_out(regs_444_io_out),
    .io_enable(regs_444_io_enable)
  );
  FringeFF regs_445 ( // @[RegFile.scala 66:20:@131220.4]
    .clock(regs_445_clock),
    .reset(regs_445_reset),
    .io_in(regs_445_io_in),
    .io_reset(regs_445_io_reset),
    .io_out(regs_445_io_out),
    .io_enable(regs_445_io_enable)
  );
  FringeFF regs_446 ( // @[RegFile.scala 66:20:@131234.4]
    .clock(regs_446_clock),
    .reset(regs_446_reset),
    .io_in(regs_446_io_in),
    .io_reset(regs_446_io_reset),
    .io_out(regs_446_io_out),
    .io_enable(regs_446_io_enable)
  );
  FringeFF regs_447 ( // @[RegFile.scala 66:20:@131248.4]
    .clock(regs_447_clock),
    .reset(regs_447_reset),
    .io_in(regs_447_io_in),
    .io_reset(regs_447_io_reset),
    .io_out(regs_447_io_out),
    .io_enable(regs_447_io_enable)
  );
  FringeFF regs_448 ( // @[RegFile.scala 66:20:@131262.4]
    .clock(regs_448_clock),
    .reset(regs_448_reset),
    .io_in(regs_448_io_in),
    .io_reset(regs_448_io_reset),
    .io_out(regs_448_io_out),
    .io_enable(regs_448_io_enable)
  );
  FringeFF regs_449 ( // @[RegFile.scala 66:20:@131276.4]
    .clock(regs_449_clock),
    .reset(regs_449_reset),
    .io_in(regs_449_io_in),
    .io_reset(regs_449_io_reset),
    .io_out(regs_449_io_out),
    .io_enable(regs_449_io_enable)
  );
  FringeFF regs_450 ( // @[RegFile.scala 66:20:@131290.4]
    .clock(regs_450_clock),
    .reset(regs_450_reset),
    .io_in(regs_450_io_in),
    .io_reset(regs_450_io_reset),
    .io_out(regs_450_io_out),
    .io_enable(regs_450_io_enable)
  );
  FringeFF regs_451 ( // @[RegFile.scala 66:20:@131304.4]
    .clock(regs_451_clock),
    .reset(regs_451_reset),
    .io_in(regs_451_io_in),
    .io_reset(regs_451_io_reset),
    .io_out(regs_451_io_out),
    .io_enable(regs_451_io_enable)
  );
  FringeFF regs_452 ( // @[RegFile.scala 66:20:@131318.4]
    .clock(regs_452_clock),
    .reset(regs_452_reset),
    .io_in(regs_452_io_in),
    .io_reset(regs_452_io_reset),
    .io_out(regs_452_io_out),
    .io_enable(regs_452_io_enable)
  );
  FringeFF regs_453 ( // @[RegFile.scala 66:20:@131332.4]
    .clock(regs_453_clock),
    .reset(regs_453_reset),
    .io_in(regs_453_io_in),
    .io_reset(regs_453_io_reset),
    .io_out(regs_453_io_out),
    .io_enable(regs_453_io_enable)
  );
  FringeFF regs_454 ( // @[RegFile.scala 66:20:@131346.4]
    .clock(regs_454_clock),
    .reset(regs_454_reset),
    .io_in(regs_454_io_in),
    .io_reset(regs_454_io_reset),
    .io_out(regs_454_io_out),
    .io_enable(regs_454_io_enable)
  );
  FringeFF regs_455 ( // @[RegFile.scala 66:20:@131360.4]
    .clock(regs_455_clock),
    .reset(regs_455_reset),
    .io_in(regs_455_io_in),
    .io_reset(regs_455_io_reset),
    .io_out(regs_455_io_out),
    .io_enable(regs_455_io_enable)
  );
  FringeFF regs_456 ( // @[RegFile.scala 66:20:@131374.4]
    .clock(regs_456_clock),
    .reset(regs_456_reset),
    .io_in(regs_456_io_in),
    .io_reset(regs_456_io_reset),
    .io_out(regs_456_io_out),
    .io_enable(regs_456_io_enable)
  );
  FringeFF regs_457 ( // @[RegFile.scala 66:20:@131388.4]
    .clock(regs_457_clock),
    .reset(regs_457_reset),
    .io_in(regs_457_io_in),
    .io_reset(regs_457_io_reset),
    .io_out(regs_457_io_out),
    .io_enable(regs_457_io_enable)
  );
  FringeFF regs_458 ( // @[RegFile.scala 66:20:@131402.4]
    .clock(regs_458_clock),
    .reset(regs_458_reset),
    .io_in(regs_458_io_in),
    .io_reset(regs_458_io_reset),
    .io_out(regs_458_io_out),
    .io_enable(regs_458_io_enable)
  );
  FringeFF regs_459 ( // @[RegFile.scala 66:20:@131416.4]
    .clock(regs_459_clock),
    .reset(regs_459_reset),
    .io_in(regs_459_io_in),
    .io_reset(regs_459_io_reset),
    .io_out(regs_459_io_out),
    .io_enable(regs_459_io_enable)
  );
  FringeFF regs_460 ( // @[RegFile.scala 66:20:@131430.4]
    .clock(regs_460_clock),
    .reset(regs_460_reset),
    .io_in(regs_460_io_in),
    .io_reset(regs_460_io_reset),
    .io_out(regs_460_io_out),
    .io_enable(regs_460_io_enable)
  );
  FringeFF regs_461 ( // @[RegFile.scala 66:20:@131444.4]
    .clock(regs_461_clock),
    .reset(regs_461_reset),
    .io_in(regs_461_io_in),
    .io_reset(regs_461_io_reset),
    .io_out(regs_461_io_out),
    .io_enable(regs_461_io_enable)
  );
  FringeFF regs_462 ( // @[RegFile.scala 66:20:@131458.4]
    .clock(regs_462_clock),
    .reset(regs_462_reset),
    .io_in(regs_462_io_in),
    .io_reset(regs_462_io_reset),
    .io_out(regs_462_io_out),
    .io_enable(regs_462_io_enable)
  );
  FringeFF regs_463 ( // @[RegFile.scala 66:20:@131472.4]
    .clock(regs_463_clock),
    .reset(regs_463_reset),
    .io_in(regs_463_io_in),
    .io_reset(regs_463_io_reset),
    .io_out(regs_463_io_out),
    .io_enable(regs_463_io_enable)
  );
  FringeFF regs_464 ( // @[RegFile.scala 66:20:@131486.4]
    .clock(regs_464_clock),
    .reset(regs_464_reset),
    .io_in(regs_464_io_in),
    .io_reset(regs_464_io_reset),
    .io_out(regs_464_io_out),
    .io_enable(regs_464_io_enable)
  );
  FringeFF regs_465 ( // @[RegFile.scala 66:20:@131500.4]
    .clock(regs_465_clock),
    .reset(regs_465_reset),
    .io_in(regs_465_io_in),
    .io_reset(regs_465_io_reset),
    .io_out(regs_465_io_out),
    .io_enable(regs_465_io_enable)
  );
  FringeFF regs_466 ( // @[RegFile.scala 66:20:@131514.4]
    .clock(regs_466_clock),
    .reset(regs_466_reset),
    .io_in(regs_466_io_in),
    .io_reset(regs_466_io_reset),
    .io_out(regs_466_io_out),
    .io_enable(regs_466_io_enable)
  );
  FringeFF regs_467 ( // @[RegFile.scala 66:20:@131528.4]
    .clock(regs_467_clock),
    .reset(regs_467_reset),
    .io_in(regs_467_io_in),
    .io_reset(regs_467_io_reset),
    .io_out(regs_467_io_out),
    .io_enable(regs_467_io_enable)
  );
  FringeFF regs_468 ( // @[RegFile.scala 66:20:@131542.4]
    .clock(regs_468_clock),
    .reset(regs_468_reset),
    .io_in(regs_468_io_in),
    .io_reset(regs_468_io_reset),
    .io_out(regs_468_io_out),
    .io_enable(regs_468_io_enable)
  );
  FringeFF regs_469 ( // @[RegFile.scala 66:20:@131556.4]
    .clock(regs_469_clock),
    .reset(regs_469_reset),
    .io_in(regs_469_io_in),
    .io_reset(regs_469_io_reset),
    .io_out(regs_469_io_out),
    .io_enable(regs_469_io_enable)
  );
  FringeFF regs_470 ( // @[RegFile.scala 66:20:@131570.4]
    .clock(regs_470_clock),
    .reset(regs_470_reset),
    .io_in(regs_470_io_in),
    .io_reset(regs_470_io_reset),
    .io_out(regs_470_io_out),
    .io_enable(regs_470_io_enable)
  );
  FringeFF regs_471 ( // @[RegFile.scala 66:20:@131584.4]
    .clock(regs_471_clock),
    .reset(regs_471_reset),
    .io_in(regs_471_io_in),
    .io_reset(regs_471_io_reset),
    .io_out(regs_471_io_out),
    .io_enable(regs_471_io_enable)
  );
  FringeFF regs_472 ( // @[RegFile.scala 66:20:@131598.4]
    .clock(regs_472_clock),
    .reset(regs_472_reset),
    .io_in(regs_472_io_in),
    .io_reset(regs_472_io_reset),
    .io_out(regs_472_io_out),
    .io_enable(regs_472_io_enable)
  );
  FringeFF regs_473 ( // @[RegFile.scala 66:20:@131612.4]
    .clock(regs_473_clock),
    .reset(regs_473_reset),
    .io_in(regs_473_io_in),
    .io_reset(regs_473_io_reset),
    .io_out(regs_473_io_out),
    .io_enable(regs_473_io_enable)
  );
  FringeFF regs_474 ( // @[RegFile.scala 66:20:@131626.4]
    .clock(regs_474_clock),
    .reset(regs_474_reset),
    .io_in(regs_474_io_in),
    .io_reset(regs_474_io_reset),
    .io_out(regs_474_io_out),
    .io_enable(regs_474_io_enable)
  );
  FringeFF regs_475 ( // @[RegFile.scala 66:20:@131640.4]
    .clock(regs_475_clock),
    .reset(regs_475_reset),
    .io_in(regs_475_io_in),
    .io_reset(regs_475_io_reset),
    .io_out(regs_475_io_out),
    .io_enable(regs_475_io_enable)
  );
  FringeFF regs_476 ( // @[RegFile.scala 66:20:@131654.4]
    .clock(regs_476_clock),
    .reset(regs_476_reset),
    .io_in(regs_476_io_in),
    .io_reset(regs_476_io_reset),
    .io_out(regs_476_io_out),
    .io_enable(regs_476_io_enable)
  );
  FringeFF regs_477 ( // @[RegFile.scala 66:20:@131668.4]
    .clock(regs_477_clock),
    .reset(regs_477_reset),
    .io_in(regs_477_io_in),
    .io_reset(regs_477_io_reset),
    .io_out(regs_477_io_out),
    .io_enable(regs_477_io_enable)
  );
  FringeFF regs_478 ( // @[RegFile.scala 66:20:@131682.4]
    .clock(regs_478_clock),
    .reset(regs_478_reset),
    .io_in(regs_478_io_in),
    .io_reset(regs_478_io_reset),
    .io_out(regs_478_io_out),
    .io_enable(regs_478_io_enable)
  );
  FringeFF regs_479 ( // @[RegFile.scala 66:20:@131696.4]
    .clock(regs_479_clock),
    .reset(regs_479_reset),
    .io_in(regs_479_io_in),
    .io_reset(regs_479_io_reset),
    .io_out(regs_479_io_out),
    .io_enable(regs_479_io_enable)
  );
  FringeFF regs_480 ( // @[RegFile.scala 66:20:@131710.4]
    .clock(regs_480_clock),
    .reset(regs_480_reset),
    .io_in(regs_480_io_in),
    .io_reset(regs_480_io_reset),
    .io_out(regs_480_io_out),
    .io_enable(regs_480_io_enable)
  );
  FringeFF regs_481 ( // @[RegFile.scala 66:20:@131724.4]
    .clock(regs_481_clock),
    .reset(regs_481_reset),
    .io_in(regs_481_io_in),
    .io_reset(regs_481_io_reset),
    .io_out(regs_481_io_out),
    .io_enable(regs_481_io_enable)
  );
  FringeFF regs_482 ( // @[RegFile.scala 66:20:@131738.4]
    .clock(regs_482_clock),
    .reset(regs_482_reset),
    .io_in(regs_482_io_in),
    .io_reset(regs_482_io_reset),
    .io_out(regs_482_io_out),
    .io_enable(regs_482_io_enable)
  );
  FringeFF regs_483 ( // @[RegFile.scala 66:20:@131752.4]
    .clock(regs_483_clock),
    .reset(regs_483_reset),
    .io_in(regs_483_io_in),
    .io_reset(regs_483_io_reset),
    .io_out(regs_483_io_out),
    .io_enable(regs_483_io_enable)
  );
  FringeFF regs_484 ( // @[RegFile.scala 66:20:@131766.4]
    .clock(regs_484_clock),
    .reset(regs_484_reset),
    .io_in(regs_484_io_in),
    .io_reset(regs_484_io_reset),
    .io_out(regs_484_io_out),
    .io_enable(regs_484_io_enable)
  );
  FringeFF regs_485 ( // @[RegFile.scala 66:20:@131780.4]
    .clock(regs_485_clock),
    .reset(regs_485_reset),
    .io_in(regs_485_io_in),
    .io_reset(regs_485_io_reset),
    .io_out(regs_485_io_out),
    .io_enable(regs_485_io_enable)
  );
  FringeFF regs_486 ( // @[RegFile.scala 66:20:@131794.4]
    .clock(regs_486_clock),
    .reset(regs_486_reset),
    .io_in(regs_486_io_in),
    .io_reset(regs_486_io_reset),
    .io_out(regs_486_io_out),
    .io_enable(regs_486_io_enable)
  );
  FringeFF regs_487 ( // @[RegFile.scala 66:20:@131808.4]
    .clock(regs_487_clock),
    .reset(regs_487_reset),
    .io_in(regs_487_io_in),
    .io_reset(regs_487_io_reset),
    .io_out(regs_487_io_out),
    .io_enable(regs_487_io_enable)
  );
  FringeFF regs_488 ( // @[RegFile.scala 66:20:@131822.4]
    .clock(regs_488_clock),
    .reset(regs_488_reset),
    .io_in(regs_488_io_in),
    .io_reset(regs_488_io_reset),
    .io_out(regs_488_io_out),
    .io_enable(regs_488_io_enable)
  );
  FringeFF regs_489 ( // @[RegFile.scala 66:20:@131836.4]
    .clock(regs_489_clock),
    .reset(regs_489_reset),
    .io_in(regs_489_io_in),
    .io_reset(regs_489_io_reset),
    .io_out(regs_489_io_out),
    .io_enable(regs_489_io_enable)
  );
  FringeFF regs_490 ( // @[RegFile.scala 66:20:@131850.4]
    .clock(regs_490_clock),
    .reset(regs_490_reset),
    .io_in(regs_490_io_in),
    .io_reset(regs_490_io_reset),
    .io_out(regs_490_io_out),
    .io_enable(regs_490_io_enable)
  );
  FringeFF regs_491 ( // @[RegFile.scala 66:20:@131864.4]
    .clock(regs_491_clock),
    .reset(regs_491_reset),
    .io_in(regs_491_io_in),
    .io_reset(regs_491_io_reset),
    .io_out(regs_491_io_out),
    .io_enable(regs_491_io_enable)
  );
  FringeFF regs_492 ( // @[RegFile.scala 66:20:@131878.4]
    .clock(regs_492_clock),
    .reset(regs_492_reset),
    .io_in(regs_492_io_in),
    .io_reset(regs_492_io_reset),
    .io_out(regs_492_io_out),
    .io_enable(regs_492_io_enable)
  );
  FringeFF regs_493 ( // @[RegFile.scala 66:20:@131892.4]
    .clock(regs_493_clock),
    .reset(regs_493_reset),
    .io_in(regs_493_io_in),
    .io_reset(regs_493_io_reset),
    .io_out(regs_493_io_out),
    .io_enable(regs_493_io_enable)
  );
  FringeFF regs_494 ( // @[RegFile.scala 66:20:@131906.4]
    .clock(regs_494_clock),
    .reset(regs_494_reset),
    .io_in(regs_494_io_in),
    .io_reset(regs_494_io_reset),
    .io_out(regs_494_io_out),
    .io_enable(regs_494_io_enable)
  );
  FringeFF regs_495 ( // @[RegFile.scala 66:20:@131920.4]
    .clock(regs_495_clock),
    .reset(regs_495_reset),
    .io_in(regs_495_io_in),
    .io_reset(regs_495_io_reset),
    .io_out(regs_495_io_out),
    .io_enable(regs_495_io_enable)
  );
  FringeFF regs_496 ( // @[RegFile.scala 66:20:@131934.4]
    .clock(regs_496_clock),
    .reset(regs_496_reset),
    .io_in(regs_496_io_in),
    .io_reset(regs_496_io_reset),
    .io_out(regs_496_io_out),
    .io_enable(regs_496_io_enable)
  );
  FringeFF regs_497 ( // @[RegFile.scala 66:20:@131948.4]
    .clock(regs_497_clock),
    .reset(regs_497_reset),
    .io_in(regs_497_io_in),
    .io_reset(regs_497_io_reset),
    .io_out(regs_497_io_out),
    .io_enable(regs_497_io_enable)
  );
  FringeFF regs_498 ( // @[RegFile.scala 66:20:@131962.4]
    .clock(regs_498_clock),
    .reset(regs_498_reset),
    .io_in(regs_498_io_in),
    .io_reset(regs_498_io_reset),
    .io_out(regs_498_io_out),
    .io_enable(regs_498_io_enable)
  );
  FringeFF regs_499 ( // @[RegFile.scala 66:20:@131976.4]
    .clock(regs_499_clock),
    .reset(regs_499_reset),
    .io_in(regs_499_io_in),
    .io_reset(regs_499_io_reset),
    .io_out(regs_499_io_out),
    .io_enable(regs_499_io_enable)
  );
  FringeFF regs_500 ( // @[RegFile.scala 66:20:@131990.4]
    .clock(regs_500_clock),
    .reset(regs_500_reset),
    .io_in(regs_500_io_in),
    .io_reset(regs_500_io_reset),
    .io_out(regs_500_io_out),
    .io_enable(regs_500_io_enable)
  );
  FringeFF regs_501 ( // @[RegFile.scala 66:20:@132004.4]
    .clock(regs_501_clock),
    .reset(regs_501_reset),
    .io_in(regs_501_io_in),
    .io_reset(regs_501_io_reset),
    .io_out(regs_501_io_out),
    .io_enable(regs_501_io_enable)
  );
  FringeFF regs_502 ( // @[RegFile.scala 66:20:@132018.4]
    .clock(regs_502_clock),
    .reset(regs_502_reset),
    .io_in(regs_502_io_in),
    .io_reset(regs_502_io_reset),
    .io_out(regs_502_io_out),
    .io_enable(regs_502_io_enable)
  );
  MuxN rport ( // @[RegFile.scala 95:21:@132032.4]
    .io_ins_0(rport_io_ins_0),
    .io_ins_1(rport_io_ins_1),
    .io_ins_2(rport_io_ins_2),
    .io_ins_3(rport_io_ins_3),
    .io_ins_4(rport_io_ins_4),
    .io_ins_5(rport_io_ins_5),
    .io_ins_6(rport_io_ins_6),
    .io_ins_7(rport_io_ins_7),
    .io_ins_8(rport_io_ins_8),
    .io_ins_9(rport_io_ins_9),
    .io_ins_10(rport_io_ins_10),
    .io_ins_11(rport_io_ins_11),
    .io_ins_12(rport_io_ins_12),
    .io_ins_13(rport_io_ins_13),
    .io_ins_14(rport_io_ins_14),
    .io_ins_15(rport_io_ins_15),
    .io_ins_16(rport_io_ins_16),
    .io_ins_17(rport_io_ins_17),
    .io_ins_18(rport_io_ins_18),
    .io_ins_19(rport_io_ins_19),
    .io_ins_20(rport_io_ins_20),
    .io_ins_21(rport_io_ins_21),
    .io_ins_22(rport_io_ins_22),
    .io_ins_23(rport_io_ins_23),
    .io_ins_24(rport_io_ins_24),
    .io_ins_25(rport_io_ins_25),
    .io_ins_26(rport_io_ins_26),
    .io_ins_27(rport_io_ins_27),
    .io_ins_28(rport_io_ins_28),
    .io_ins_29(rport_io_ins_29),
    .io_ins_30(rport_io_ins_30),
    .io_ins_31(rport_io_ins_31),
    .io_ins_32(rport_io_ins_32),
    .io_ins_33(rport_io_ins_33),
    .io_ins_34(rport_io_ins_34),
    .io_ins_35(rport_io_ins_35),
    .io_ins_36(rport_io_ins_36),
    .io_ins_37(rport_io_ins_37),
    .io_ins_38(rport_io_ins_38),
    .io_ins_39(rport_io_ins_39),
    .io_ins_40(rport_io_ins_40),
    .io_ins_41(rport_io_ins_41),
    .io_ins_42(rport_io_ins_42),
    .io_ins_43(rport_io_ins_43),
    .io_ins_44(rport_io_ins_44),
    .io_ins_45(rport_io_ins_45),
    .io_ins_46(rport_io_ins_46),
    .io_ins_47(rport_io_ins_47),
    .io_ins_48(rport_io_ins_48),
    .io_ins_49(rport_io_ins_49),
    .io_ins_50(rport_io_ins_50),
    .io_ins_51(rport_io_ins_51),
    .io_ins_52(rport_io_ins_52),
    .io_ins_53(rport_io_ins_53),
    .io_ins_54(rport_io_ins_54),
    .io_ins_55(rport_io_ins_55),
    .io_ins_56(rport_io_ins_56),
    .io_ins_57(rport_io_ins_57),
    .io_ins_58(rport_io_ins_58),
    .io_ins_59(rport_io_ins_59),
    .io_ins_60(rport_io_ins_60),
    .io_ins_61(rport_io_ins_61),
    .io_ins_62(rport_io_ins_62),
    .io_ins_63(rport_io_ins_63),
    .io_ins_64(rport_io_ins_64),
    .io_ins_65(rport_io_ins_65),
    .io_ins_66(rport_io_ins_66),
    .io_ins_67(rport_io_ins_67),
    .io_ins_68(rport_io_ins_68),
    .io_ins_69(rport_io_ins_69),
    .io_ins_70(rport_io_ins_70),
    .io_ins_71(rport_io_ins_71),
    .io_ins_72(rport_io_ins_72),
    .io_ins_73(rport_io_ins_73),
    .io_ins_74(rport_io_ins_74),
    .io_ins_75(rport_io_ins_75),
    .io_ins_76(rport_io_ins_76),
    .io_ins_77(rport_io_ins_77),
    .io_ins_78(rport_io_ins_78),
    .io_ins_79(rport_io_ins_79),
    .io_ins_80(rport_io_ins_80),
    .io_ins_81(rport_io_ins_81),
    .io_ins_82(rport_io_ins_82),
    .io_ins_83(rport_io_ins_83),
    .io_ins_84(rport_io_ins_84),
    .io_ins_85(rport_io_ins_85),
    .io_ins_86(rport_io_ins_86),
    .io_ins_87(rport_io_ins_87),
    .io_ins_88(rport_io_ins_88),
    .io_ins_89(rport_io_ins_89),
    .io_ins_90(rport_io_ins_90),
    .io_ins_91(rport_io_ins_91),
    .io_ins_92(rport_io_ins_92),
    .io_ins_93(rport_io_ins_93),
    .io_ins_94(rport_io_ins_94),
    .io_ins_95(rport_io_ins_95),
    .io_ins_96(rport_io_ins_96),
    .io_ins_97(rport_io_ins_97),
    .io_ins_98(rport_io_ins_98),
    .io_ins_99(rport_io_ins_99),
    .io_ins_100(rport_io_ins_100),
    .io_ins_101(rport_io_ins_101),
    .io_ins_102(rport_io_ins_102),
    .io_ins_103(rport_io_ins_103),
    .io_ins_104(rport_io_ins_104),
    .io_ins_105(rport_io_ins_105),
    .io_ins_106(rport_io_ins_106),
    .io_ins_107(rport_io_ins_107),
    .io_ins_108(rport_io_ins_108),
    .io_ins_109(rport_io_ins_109),
    .io_ins_110(rport_io_ins_110),
    .io_ins_111(rport_io_ins_111),
    .io_ins_112(rport_io_ins_112),
    .io_ins_113(rport_io_ins_113),
    .io_ins_114(rport_io_ins_114),
    .io_ins_115(rport_io_ins_115),
    .io_ins_116(rport_io_ins_116),
    .io_ins_117(rport_io_ins_117),
    .io_ins_118(rport_io_ins_118),
    .io_ins_119(rport_io_ins_119),
    .io_ins_120(rport_io_ins_120),
    .io_ins_121(rport_io_ins_121),
    .io_ins_122(rport_io_ins_122),
    .io_ins_123(rport_io_ins_123),
    .io_ins_124(rport_io_ins_124),
    .io_ins_125(rport_io_ins_125),
    .io_ins_126(rport_io_ins_126),
    .io_ins_127(rport_io_ins_127),
    .io_ins_128(rport_io_ins_128),
    .io_ins_129(rport_io_ins_129),
    .io_ins_130(rport_io_ins_130),
    .io_ins_131(rport_io_ins_131),
    .io_ins_132(rport_io_ins_132),
    .io_ins_133(rport_io_ins_133),
    .io_ins_134(rport_io_ins_134),
    .io_ins_135(rport_io_ins_135),
    .io_ins_136(rport_io_ins_136),
    .io_ins_137(rport_io_ins_137),
    .io_ins_138(rport_io_ins_138),
    .io_ins_139(rport_io_ins_139),
    .io_ins_140(rport_io_ins_140),
    .io_ins_141(rport_io_ins_141),
    .io_ins_142(rport_io_ins_142),
    .io_ins_143(rport_io_ins_143),
    .io_ins_144(rport_io_ins_144),
    .io_ins_145(rport_io_ins_145),
    .io_ins_146(rport_io_ins_146),
    .io_ins_147(rport_io_ins_147),
    .io_ins_148(rport_io_ins_148),
    .io_ins_149(rport_io_ins_149),
    .io_ins_150(rport_io_ins_150),
    .io_ins_151(rport_io_ins_151),
    .io_ins_152(rport_io_ins_152),
    .io_ins_153(rport_io_ins_153),
    .io_ins_154(rport_io_ins_154),
    .io_ins_155(rport_io_ins_155),
    .io_ins_156(rport_io_ins_156),
    .io_ins_157(rport_io_ins_157),
    .io_ins_158(rport_io_ins_158),
    .io_ins_159(rport_io_ins_159),
    .io_ins_160(rport_io_ins_160),
    .io_ins_161(rport_io_ins_161),
    .io_ins_162(rport_io_ins_162),
    .io_ins_163(rport_io_ins_163),
    .io_ins_164(rport_io_ins_164),
    .io_ins_165(rport_io_ins_165),
    .io_ins_166(rport_io_ins_166),
    .io_ins_167(rport_io_ins_167),
    .io_ins_168(rport_io_ins_168),
    .io_ins_169(rport_io_ins_169),
    .io_ins_170(rport_io_ins_170),
    .io_ins_171(rport_io_ins_171),
    .io_ins_172(rport_io_ins_172),
    .io_ins_173(rport_io_ins_173),
    .io_ins_174(rport_io_ins_174),
    .io_ins_175(rport_io_ins_175),
    .io_ins_176(rport_io_ins_176),
    .io_ins_177(rport_io_ins_177),
    .io_ins_178(rport_io_ins_178),
    .io_ins_179(rport_io_ins_179),
    .io_ins_180(rport_io_ins_180),
    .io_ins_181(rport_io_ins_181),
    .io_ins_182(rport_io_ins_182),
    .io_ins_183(rport_io_ins_183),
    .io_ins_184(rport_io_ins_184),
    .io_ins_185(rport_io_ins_185),
    .io_ins_186(rport_io_ins_186),
    .io_ins_187(rport_io_ins_187),
    .io_ins_188(rport_io_ins_188),
    .io_ins_189(rport_io_ins_189),
    .io_ins_190(rport_io_ins_190),
    .io_ins_191(rport_io_ins_191),
    .io_ins_192(rport_io_ins_192),
    .io_ins_193(rport_io_ins_193),
    .io_ins_194(rport_io_ins_194),
    .io_ins_195(rport_io_ins_195),
    .io_ins_196(rport_io_ins_196),
    .io_ins_197(rport_io_ins_197),
    .io_ins_198(rport_io_ins_198),
    .io_ins_199(rport_io_ins_199),
    .io_ins_200(rport_io_ins_200),
    .io_ins_201(rport_io_ins_201),
    .io_ins_202(rport_io_ins_202),
    .io_ins_203(rport_io_ins_203),
    .io_ins_204(rport_io_ins_204),
    .io_ins_205(rport_io_ins_205),
    .io_ins_206(rport_io_ins_206),
    .io_ins_207(rport_io_ins_207),
    .io_ins_208(rport_io_ins_208),
    .io_ins_209(rport_io_ins_209),
    .io_ins_210(rport_io_ins_210),
    .io_ins_211(rport_io_ins_211),
    .io_ins_212(rport_io_ins_212),
    .io_ins_213(rport_io_ins_213),
    .io_ins_214(rport_io_ins_214),
    .io_ins_215(rport_io_ins_215),
    .io_ins_216(rport_io_ins_216),
    .io_ins_217(rport_io_ins_217),
    .io_ins_218(rport_io_ins_218),
    .io_ins_219(rport_io_ins_219),
    .io_ins_220(rport_io_ins_220),
    .io_ins_221(rport_io_ins_221),
    .io_ins_222(rport_io_ins_222),
    .io_ins_223(rport_io_ins_223),
    .io_ins_224(rport_io_ins_224),
    .io_ins_225(rport_io_ins_225),
    .io_ins_226(rport_io_ins_226),
    .io_ins_227(rport_io_ins_227),
    .io_ins_228(rport_io_ins_228),
    .io_ins_229(rport_io_ins_229),
    .io_ins_230(rport_io_ins_230),
    .io_ins_231(rport_io_ins_231),
    .io_ins_232(rport_io_ins_232),
    .io_ins_233(rport_io_ins_233),
    .io_ins_234(rport_io_ins_234),
    .io_ins_235(rport_io_ins_235),
    .io_ins_236(rport_io_ins_236),
    .io_ins_237(rport_io_ins_237),
    .io_ins_238(rport_io_ins_238),
    .io_ins_239(rport_io_ins_239),
    .io_ins_240(rport_io_ins_240),
    .io_ins_241(rport_io_ins_241),
    .io_ins_242(rport_io_ins_242),
    .io_ins_243(rport_io_ins_243),
    .io_ins_244(rport_io_ins_244),
    .io_ins_245(rport_io_ins_245),
    .io_ins_246(rport_io_ins_246),
    .io_ins_247(rport_io_ins_247),
    .io_ins_248(rport_io_ins_248),
    .io_ins_249(rport_io_ins_249),
    .io_ins_250(rport_io_ins_250),
    .io_ins_251(rport_io_ins_251),
    .io_ins_252(rport_io_ins_252),
    .io_ins_253(rport_io_ins_253),
    .io_ins_254(rport_io_ins_254),
    .io_ins_255(rport_io_ins_255),
    .io_ins_256(rport_io_ins_256),
    .io_ins_257(rport_io_ins_257),
    .io_ins_258(rport_io_ins_258),
    .io_ins_259(rport_io_ins_259),
    .io_ins_260(rport_io_ins_260),
    .io_ins_261(rport_io_ins_261),
    .io_ins_262(rport_io_ins_262),
    .io_ins_263(rport_io_ins_263),
    .io_ins_264(rport_io_ins_264),
    .io_ins_265(rport_io_ins_265),
    .io_ins_266(rport_io_ins_266),
    .io_ins_267(rport_io_ins_267),
    .io_ins_268(rport_io_ins_268),
    .io_ins_269(rport_io_ins_269),
    .io_ins_270(rport_io_ins_270),
    .io_ins_271(rport_io_ins_271),
    .io_ins_272(rport_io_ins_272),
    .io_ins_273(rport_io_ins_273),
    .io_ins_274(rport_io_ins_274),
    .io_ins_275(rport_io_ins_275),
    .io_ins_276(rport_io_ins_276),
    .io_ins_277(rport_io_ins_277),
    .io_ins_278(rport_io_ins_278),
    .io_ins_279(rport_io_ins_279),
    .io_ins_280(rport_io_ins_280),
    .io_ins_281(rport_io_ins_281),
    .io_ins_282(rport_io_ins_282),
    .io_ins_283(rport_io_ins_283),
    .io_ins_284(rport_io_ins_284),
    .io_ins_285(rport_io_ins_285),
    .io_ins_286(rport_io_ins_286),
    .io_ins_287(rport_io_ins_287),
    .io_ins_288(rport_io_ins_288),
    .io_ins_289(rport_io_ins_289),
    .io_ins_290(rport_io_ins_290),
    .io_ins_291(rport_io_ins_291),
    .io_ins_292(rport_io_ins_292),
    .io_ins_293(rport_io_ins_293),
    .io_ins_294(rport_io_ins_294),
    .io_ins_295(rport_io_ins_295),
    .io_ins_296(rport_io_ins_296),
    .io_ins_297(rport_io_ins_297),
    .io_ins_298(rport_io_ins_298),
    .io_ins_299(rport_io_ins_299),
    .io_ins_300(rport_io_ins_300),
    .io_ins_301(rport_io_ins_301),
    .io_ins_302(rport_io_ins_302),
    .io_ins_303(rport_io_ins_303),
    .io_ins_304(rport_io_ins_304),
    .io_ins_305(rport_io_ins_305),
    .io_ins_306(rport_io_ins_306),
    .io_ins_307(rport_io_ins_307),
    .io_ins_308(rport_io_ins_308),
    .io_ins_309(rport_io_ins_309),
    .io_ins_310(rport_io_ins_310),
    .io_ins_311(rport_io_ins_311),
    .io_ins_312(rport_io_ins_312),
    .io_ins_313(rport_io_ins_313),
    .io_ins_314(rport_io_ins_314),
    .io_ins_315(rport_io_ins_315),
    .io_ins_316(rport_io_ins_316),
    .io_ins_317(rport_io_ins_317),
    .io_ins_318(rport_io_ins_318),
    .io_ins_319(rport_io_ins_319),
    .io_ins_320(rport_io_ins_320),
    .io_ins_321(rport_io_ins_321),
    .io_ins_322(rport_io_ins_322),
    .io_ins_323(rport_io_ins_323),
    .io_ins_324(rport_io_ins_324),
    .io_ins_325(rport_io_ins_325),
    .io_ins_326(rport_io_ins_326),
    .io_ins_327(rport_io_ins_327),
    .io_ins_328(rport_io_ins_328),
    .io_ins_329(rport_io_ins_329),
    .io_ins_330(rport_io_ins_330),
    .io_ins_331(rport_io_ins_331),
    .io_ins_332(rport_io_ins_332),
    .io_ins_333(rport_io_ins_333),
    .io_ins_334(rport_io_ins_334),
    .io_ins_335(rport_io_ins_335),
    .io_ins_336(rport_io_ins_336),
    .io_ins_337(rport_io_ins_337),
    .io_ins_338(rport_io_ins_338),
    .io_ins_339(rport_io_ins_339),
    .io_ins_340(rport_io_ins_340),
    .io_ins_341(rport_io_ins_341),
    .io_ins_342(rport_io_ins_342),
    .io_ins_343(rport_io_ins_343),
    .io_ins_344(rport_io_ins_344),
    .io_ins_345(rport_io_ins_345),
    .io_ins_346(rport_io_ins_346),
    .io_ins_347(rport_io_ins_347),
    .io_ins_348(rport_io_ins_348),
    .io_ins_349(rport_io_ins_349),
    .io_ins_350(rport_io_ins_350),
    .io_ins_351(rport_io_ins_351),
    .io_ins_352(rport_io_ins_352),
    .io_ins_353(rport_io_ins_353),
    .io_ins_354(rport_io_ins_354),
    .io_ins_355(rport_io_ins_355),
    .io_ins_356(rport_io_ins_356),
    .io_ins_357(rport_io_ins_357),
    .io_ins_358(rport_io_ins_358),
    .io_ins_359(rport_io_ins_359),
    .io_ins_360(rport_io_ins_360),
    .io_ins_361(rport_io_ins_361),
    .io_ins_362(rport_io_ins_362),
    .io_ins_363(rport_io_ins_363),
    .io_ins_364(rport_io_ins_364),
    .io_ins_365(rport_io_ins_365),
    .io_ins_366(rport_io_ins_366),
    .io_ins_367(rport_io_ins_367),
    .io_ins_368(rport_io_ins_368),
    .io_ins_369(rport_io_ins_369),
    .io_ins_370(rport_io_ins_370),
    .io_ins_371(rport_io_ins_371),
    .io_ins_372(rport_io_ins_372),
    .io_ins_373(rport_io_ins_373),
    .io_ins_374(rport_io_ins_374),
    .io_ins_375(rport_io_ins_375),
    .io_ins_376(rport_io_ins_376),
    .io_ins_377(rport_io_ins_377),
    .io_ins_378(rport_io_ins_378),
    .io_ins_379(rport_io_ins_379),
    .io_ins_380(rport_io_ins_380),
    .io_ins_381(rport_io_ins_381),
    .io_ins_382(rport_io_ins_382),
    .io_ins_383(rport_io_ins_383),
    .io_ins_384(rport_io_ins_384),
    .io_ins_385(rport_io_ins_385),
    .io_ins_386(rport_io_ins_386),
    .io_ins_387(rport_io_ins_387),
    .io_ins_388(rport_io_ins_388),
    .io_ins_389(rport_io_ins_389),
    .io_ins_390(rport_io_ins_390),
    .io_ins_391(rport_io_ins_391),
    .io_ins_392(rport_io_ins_392),
    .io_ins_393(rport_io_ins_393),
    .io_ins_394(rport_io_ins_394),
    .io_ins_395(rport_io_ins_395),
    .io_ins_396(rport_io_ins_396),
    .io_ins_397(rport_io_ins_397),
    .io_ins_398(rport_io_ins_398),
    .io_ins_399(rport_io_ins_399),
    .io_ins_400(rport_io_ins_400),
    .io_ins_401(rport_io_ins_401),
    .io_ins_402(rport_io_ins_402),
    .io_ins_403(rport_io_ins_403),
    .io_ins_404(rport_io_ins_404),
    .io_ins_405(rport_io_ins_405),
    .io_ins_406(rport_io_ins_406),
    .io_ins_407(rport_io_ins_407),
    .io_ins_408(rport_io_ins_408),
    .io_ins_409(rport_io_ins_409),
    .io_ins_410(rport_io_ins_410),
    .io_ins_411(rport_io_ins_411),
    .io_ins_412(rport_io_ins_412),
    .io_ins_413(rport_io_ins_413),
    .io_ins_414(rport_io_ins_414),
    .io_ins_415(rport_io_ins_415),
    .io_ins_416(rport_io_ins_416),
    .io_ins_417(rport_io_ins_417),
    .io_ins_418(rport_io_ins_418),
    .io_ins_419(rport_io_ins_419),
    .io_ins_420(rport_io_ins_420),
    .io_ins_421(rport_io_ins_421),
    .io_ins_422(rport_io_ins_422),
    .io_ins_423(rport_io_ins_423),
    .io_ins_424(rport_io_ins_424),
    .io_ins_425(rport_io_ins_425),
    .io_ins_426(rport_io_ins_426),
    .io_ins_427(rport_io_ins_427),
    .io_ins_428(rport_io_ins_428),
    .io_ins_429(rport_io_ins_429),
    .io_ins_430(rport_io_ins_430),
    .io_ins_431(rport_io_ins_431),
    .io_ins_432(rport_io_ins_432),
    .io_ins_433(rport_io_ins_433),
    .io_ins_434(rport_io_ins_434),
    .io_ins_435(rport_io_ins_435),
    .io_ins_436(rport_io_ins_436),
    .io_ins_437(rport_io_ins_437),
    .io_ins_438(rport_io_ins_438),
    .io_ins_439(rport_io_ins_439),
    .io_ins_440(rport_io_ins_440),
    .io_ins_441(rport_io_ins_441),
    .io_ins_442(rport_io_ins_442),
    .io_ins_443(rport_io_ins_443),
    .io_ins_444(rport_io_ins_444),
    .io_ins_445(rport_io_ins_445),
    .io_ins_446(rport_io_ins_446),
    .io_ins_447(rport_io_ins_447),
    .io_ins_448(rport_io_ins_448),
    .io_ins_449(rport_io_ins_449),
    .io_ins_450(rport_io_ins_450),
    .io_ins_451(rport_io_ins_451),
    .io_ins_452(rport_io_ins_452),
    .io_ins_453(rport_io_ins_453),
    .io_ins_454(rport_io_ins_454),
    .io_ins_455(rport_io_ins_455),
    .io_ins_456(rport_io_ins_456),
    .io_ins_457(rport_io_ins_457),
    .io_ins_458(rport_io_ins_458),
    .io_ins_459(rport_io_ins_459),
    .io_ins_460(rport_io_ins_460),
    .io_ins_461(rport_io_ins_461),
    .io_ins_462(rport_io_ins_462),
    .io_ins_463(rport_io_ins_463),
    .io_ins_464(rport_io_ins_464),
    .io_ins_465(rport_io_ins_465),
    .io_ins_466(rport_io_ins_466),
    .io_ins_467(rport_io_ins_467),
    .io_ins_468(rport_io_ins_468),
    .io_ins_469(rport_io_ins_469),
    .io_ins_470(rport_io_ins_470),
    .io_ins_471(rport_io_ins_471),
    .io_ins_472(rport_io_ins_472),
    .io_ins_473(rport_io_ins_473),
    .io_ins_474(rport_io_ins_474),
    .io_ins_475(rport_io_ins_475),
    .io_ins_476(rport_io_ins_476),
    .io_ins_477(rport_io_ins_477),
    .io_ins_478(rport_io_ins_478),
    .io_ins_479(rport_io_ins_479),
    .io_ins_480(rport_io_ins_480),
    .io_ins_481(rport_io_ins_481),
    .io_ins_482(rport_io_ins_482),
    .io_ins_483(rport_io_ins_483),
    .io_ins_484(rport_io_ins_484),
    .io_ins_485(rport_io_ins_485),
    .io_ins_486(rport_io_ins_486),
    .io_ins_487(rport_io_ins_487),
    .io_ins_488(rport_io_ins_488),
    .io_ins_489(rport_io_ins_489),
    .io_ins_490(rport_io_ins_490),
    .io_ins_491(rport_io_ins_491),
    .io_ins_492(rport_io_ins_492),
    .io_ins_493(rport_io_ins_493),
    .io_ins_494(rport_io_ins_494),
    .io_ins_495(rport_io_ins_495),
    .io_ins_496(rport_io_ins_496),
    .io_ins_497(rport_io_ins_497),
    .io_ins_498(rport_io_ins_498),
    .io_ins_499(rport_io_ins_499),
    .io_ins_500(rport_io_ins_500),
    .io_ins_501(rport_io_ins_501),
    .io_ins_502(rport_io_ins_502),
    .io_sel(rport_io_sel),
    .io_out(rport_io_out)
  );
  assign _T_3078 = io_waddr == 32'h0; // @[RegFile.scala 80:42:@124994.4]
  assign _T_3084 = io_waddr == 32'h1; // @[RegFile.scala 68:46:@125006.4]
  assign _T_3085 = io_wen & _T_3084; // @[RegFile.scala 68:34:@125007.4]
  assign _T_3098 = io_waddr == 32'h2; // @[RegFile.scala 80:42:@125025.4]
  assign _T_3104 = io_waddr == 32'h3; // @[RegFile.scala 80:42:@125037.4]
  assign _T_3110 = io_waddr == 32'h4; // @[RegFile.scala 74:80:@125049.4]
  assign _T_3111 = io_wen & _T_3110; // @[RegFile.scala 74:68:@125050.4]
  assign io_rdata = rport_io_out; // @[RegFile.scala 107:14:@133043.4]
  assign io_argIns_0 = regs_0_io_out; // @[RegFile.scala 111:13:@133049.4]
  assign io_argIns_1 = regs_1_io_out; // @[RegFile.scala 111:13:@133050.4]
  assign io_argIns_2 = regs_2_io_out; // @[RegFile.scala 111:13:@133051.4]
  assign io_argIns_3 = regs_3_io_out; // @[RegFile.scala 111:13:@133052.4]
  assign regs_0_clock = clock; // @[:@124992.4]
  assign regs_0_reset = reset; // @[:@124993.4 RegFile.scala 82:16:@124999.4]
  assign regs_0_io_in = io_wdata; // @[RegFile.scala 81:16:@124997.4]
  assign regs_0_io_reset = reset; // @[RegFile.scala 83:19:@125001.4]
  assign regs_0_io_enable = io_wen & _T_3078; // @[RegFile.scala 80:20:@124996.4]
  assign regs_1_clock = clock; // @[:@125004.4]
  assign regs_1_reset = reset; // @[:@125005.4 RegFile.scala 70:16:@125017.4]
  assign regs_1_io_in = _T_3085 ? io_wdata : io_argOuts_0_bits; // @[RegFile.scala 69:16:@125015.4]
  assign regs_1_io_reset = reset; // @[RegFile.scala 72:19:@125020.4]
  assign regs_1_io_enable = _T_3085 ? _T_3085 : io_argOuts_0_valid; // @[RegFile.scala 68:20:@125011.4]
  assign regs_2_clock = clock; // @[:@125023.4]
  assign regs_2_reset = reset; // @[:@125024.4 RegFile.scala 82:16:@125030.4]
  assign regs_2_io_in = io_wdata; // @[RegFile.scala 81:16:@125028.4]
  assign regs_2_io_reset = reset; // @[RegFile.scala 83:19:@125032.4]
  assign regs_2_io_enable = io_wen & _T_3098; // @[RegFile.scala 80:20:@125027.4]
  assign regs_3_clock = clock; // @[:@125035.4]
  assign regs_3_reset = reset; // @[:@125036.4 RegFile.scala 82:16:@125042.4]
  assign regs_3_io_in = io_wdata; // @[RegFile.scala 81:16:@125040.4]
  assign regs_3_io_reset = reset; // @[RegFile.scala 83:19:@125044.4]
  assign regs_3_io_enable = io_wen & _T_3104; // @[RegFile.scala 80:20:@125039.4]
  assign regs_4_clock = clock; // @[:@125047.4]
  assign regs_4_reset = io_reset; // @[:@125048.4 RegFile.scala 76:16:@125055.4]
  assign regs_4_io_in = io_argOuts_1_valid ? io_argOuts_1_bits : io_wdata; // @[RegFile.scala 75:16:@125054.4]
  assign regs_4_io_reset = reset; // @[RegFile.scala 78:19:@125058.4]
  assign regs_4_io_enable = io_argOuts_1_valid | _T_3111; // @[RegFile.scala 74:20:@125052.4]
  assign regs_5_clock = clock; // @[:@125061.4]
  assign regs_5_reset = io_reset; // @[:@125062.4 RegFile.scala 76:16:@125069.4]
  assign regs_5_io_in = 64'h0; // @[RegFile.scala 75:16:@125068.4]
  assign regs_5_io_reset = reset; // @[RegFile.scala 78:19:@125072.4]
  assign regs_5_io_enable = 1'h1; // @[RegFile.scala 74:20:@125066.4]
  assign regs_6_clock = clock; // @[:@125075.4]
  assign regs_6_reset = io_reset; // @[:@125076.4 RegFile.scala 76:16:@125083.4]
  assign regs_6_io_in = 64'h0; // @[RegFile.scala 75:16:@125082.4]
  assign regs_6_io_reset = reset; // @[RegFile.scala 78:19:@125086.4]
  assign regs_6_io_enable = 1'h1; // @[RegFile.scala 74:20:@125080.4]
  assign regs_7_clock = clock; // @[:@125089.4]
  assign regs_7_reset = io_reset; // @[:@125090.4 RegFile.scala 76:16:@125097.4]
  assign regs_7_io_in = 64'h0; // @[RegFile.scala 75:16:@125096.4]
  assign regs_7_io_reset = reset; // @[RegFile.scala 78:19:@125100.4]
  assign regs_7_io_enable = 1'h1; // @[RegFile.scala 74:20:@125094.4]
  assign regs_8_clock = clock; // @[:@125103.4]
  assign regs_8_reset = io_reset; // @[:@125104.4 RegFile.scala 76:16:@125111.4]
  assign regs_8_io_in = 64'h0; // @[RegFile.scala 75:16:@125110.4]
  assign regs_8_io_reset = reset; // @[RegFile.scala 78:19:@125114.4]
  assign regs_8_io_enable = 1'h1; // @[RegFile.scala 74:20:@125108.4]
  assign regs_9_clock = clock; // @[:@125117.4]
  assign regs_9_reset = io_reset; // @[:@125118.4 RegFile.scala 76:16:@125125.4]
  assign regs_9_io_in = 64'h0; // @[RegFile.scala 75:16:@125124.4]
  assign regs_9_io_reset = reset; // @[RegFile.scala 78:19:@125128.4]
  assign regs_9_io_enable = 1'h1; // @[RegFile.scala 74:20:@125122.4]
  assign regs_10_clock = clock; // @[:@125131.4]
  assign regs_10_reset = io_reset; // @[:@125132.4 RegFile.scala 76:16:@125139.4]
  assign regs_10_io_in = 64'h0; // @[RegFile.scala 75:16:@125138.4]
  assign regs_10_io_reset = reset; // @[RegFile.scala 78:19:@125142.4]
  assign regs_10_io_enable = 1'h1; // @[RegFile.scala 74:20:@125136.4]
  assign regs_11_clock = clock; // @[:@125145.4]
  assign regs_11_reset = io_reset; // @[:@125146.4 RegFile.scala 76:16:@125153.4]
  assign regs_11_io_in = 64'h0; // @[RegFile.scala 75:16:@125152.4]
  assign regs_11_io_reset = reset; // @[RegFile.scala 78:19:@125156.4]
  assign regs_11_io_enable = 1'h1; // @[RegFile.scala 74:20:@125150.4]
  assign regs_12_clock = clock; // @[:@125159.4]
  assign regs_12_reset = io_reset; // @[:@125160.4 RegFile.scala 76:16:@125167.4]
  assign regs_12_io_in = 64'h0; // @[RegFile.scala 75:16:@125166.4]
  assign regs_12_io_reset = reset; // @[RegFile.scala 78:19:@125170.4]
  assign regs_12_io_enable = 1'h1; // @[RegFile.scala 74:20:@125164.4]
  assign regs_13_clock = clock; // @[:@125173.4]
  assign regs_13_reset = io_reset; // @[:@125174.4 RegFile.scala 76:16:@125181.4]
  assign regs_13_io_in = 64'h0; // @[RegFile.scala 75:16:@125180.4]
  assign regs_13_io_reset = reset; // @[RegFile.scala 78:19:@125184.4]
  assign regs_13_io_enable = 1'h1; // @[RegFile.scala 74:20:@125178.4]
  assign regs_14_clock = clock; // @[:@125187.4]
  assign regs_14_reset = io_reset; // @[:@125188.4 RegFile.scala 76:16:@125195.4]
  assign regs_14_io_in = 64'h0; // @[RegFile.scala 75:16:@125194.4]
  assign regs_14_io_reset = reset; // @[RegFile.scala 78:19:@125198.4]
  assign regs_14_io_enable = 1'h1; // @[RegFile.scala 74:20:@125192.4]
  assign regs_15_clock = clock; // @[:@125201.4]
  assign regs_15_reset = io_reset; // @[:@125202.4 RegFile.scala 76:16:@125209.4]
  assign regs_15_io_in = 64'h0; // @[RegFile.scala 75:16:@125208.4]
  assign regs_15_io_reset = reset; // @[RegFile.scala 78:19:@125212.4]
  assign regs_15_io_enable = 1'h1; // @[RegFile.scala 74:20:@125206.4]
  assign regs_16_clock = clock; // @[:@125215.4]
  assign regs_16_reset = io_reset; // @[:@125216.4 RegFile.scala 76:16:@125223.4]
  assign regs_16_io_in = 64'h0; // @[RegFile.scala 75:16:@125222.4]
  assign regs_16_io_reset = reset; // @[RegFile.scala 78:19:@125226.4]
  assign regs_16_io_enable = 1'h1; // @[RegFile.scala 74:20:@125220.4]
  assign regs_17_clock = clock; // @[:@125229.4]
  assign regs_17_reset = io_reset; // @[:@125230.4 RegFile.scala 76:16:@125237.4]
  assign regs_17_io_in = 64'h0; // @[RegFile.scala 75:16:@125236.4]
  assign regs_17_io_reset = reset; // @[RegFile.scala 78:19:@125240.4]
  assign regs_17_io_enable = 1'h1; // @[RegFile.scala 74:20:@125234.4]
  assign regs_18_clock = clock; // @[:@125243.4]
  assign regs_18_reset = io_reset; // @[:@125244.4 RegFile.scala 76:16:@125251.4]
  assign regs_18_io_in = 64'h0; // @[RegFile.scala 75:16:@125250.4]
  assign regs_18_io_reset = reset; // @[RegFile.scala 78:19:@125254.4]
  assign regs_18_io_enable = 1'h1; // @[RegFile.scala 74:20:@125248.4]
  assign regs_19_clock = clock; // @[:@125257.4]
  assign regs_19_reset = io_reset; // @[:@125258.4 RegFile.scala 76:16:@125265.4]
  assign regs_19_io_in = 64'h0; // @[RegFile.scala 75:16:@125264.4]
  assign regs_19_io_reset = reset; // @[RegFile.scala 78:19:@125268.4]
  assign regs_19_io_enable = 1'h1; // @[RegFile.scala 74:20:@125262.4]
  assign regs_20_clock = clock; // @[:@125271.4]
  assign regs_20_reset = io_reset; // @[:@125272.4 RegFile.scala 76:16:@125279.4]
  assign regs_20_io_in = 64'h0; // @[RegFile.scala 75:16:@125278.4]
  assign regs_20_io_reset = reset; // @[RegFile.scala 78:19:@125282.4]
  assign regs_20_io_enable = 1'h1; // @[RegFile.scala 74:20:@125276.4]
  assign regs_21_clock = clock; // @[:@125285.4]
  assign regs_21_reset = io_reset; // @[:@125286.4 RegFile.scala 76:16:@125293.4]
  assign regs_21_io_in = 64'h0; // @[RegFile.scala 75:16:@125292.4]
  assign regs_21_io_reset = reset; // @[RegFile.scala 78:19:@125296.4]
  assign regs_21_io_enable = 1'h1; // @[RegFile.scala 74:20:@125290.4]
  assign regs_22_clock = clock; // @[:@125299.4]
  assign regs_22_reset = io_reset; // @[:@125300.4 RegFile.scala 76:16:@125307.4]
  assign regs_22_io_in = 64'h0; // @[RegFile.scala 75:16:@125306.4]
  assign regs_22_io_reset = reset; // @[RegFile.scala 78:19:@125310.4]
  assign regs_22_io_enable = 1'h1; // @[RegFile.scala 74:20:@125304.4]
  assign regs_23_clock = clock; // @[:@125313.4]
  assign regs_23_reset = io_reset; // @[:@125314.4 RegFile.scala 76:16:@125321.4]
  assign regs_23_io_in = 64'h0; // @[RegFile.scala 75:16:@125320.4]
  assign regs_23_io_reset = reset; // @[RegFile.scala 78:19:@125324.4]
  assign regs_23_io_enable = 1'h1; // @[RegFile.scala 74:20:@125318.4]
  assign regs_24_clock = clock; // @[:@125327.4]
  assign regs_24_reset = io_reset; // @[:@125328.4 RegFile.scala 76:16:@125335.4]
  assign regs_24_io_in = 64'h0; // @[RegFile.scala 75:16:@125334.4]
  assign regs_24_io_reset = reset; // @[RegFile.scala 78:19:@125338.4]
  assign regs_24_io_enable = 1'h1; // @[RegFile.scala 74:20:@125332.4]
  assign regs_25_clock = clock; // @[:@125341.4]
  assign regs_25_reset = io_reset; // @[:@125342.4 RegFile.scala 76:16:@125349.4]
  assign regs_25_io_in = 64'h0; // @[RegFile.scala 75:16:@125348.4]
  assign regs_25_io_reset = reset; // @[RegFile.scala 78:19:@125352.4]
  assign regs_25_io_enable = 1'h1; // @[RegFile.scala 74:20:@125346.4]
  assign regs_26_clock = clock; // @[:@125355.4]
  assign regs_26_reset = io_reset; // @[:@125356.4 RegFile.scala 76:16:@125363.4]
  assign regs_26_io_in = 64'h0; // @[RegFile.scala 75:16:@125362.4]
  assign regs_26_io_reset = reset; // @[RegFile.scala 78:19:@125366.4]
  assign regs_26_io_enable = 1'h1; // @[RegFile.scala 74:20:@125360.4]
  assign regs_27_clock = clock; // @[:@125369.4]
  assign regs_27_reset = io_reset; // @[:@125370.4 RegFile.scala 76:16:@125377.4]
  assign regs_27_io_in = 64'h0; // @[RegFile.scala 75:16:@125376.4]
  assign regs_27_io_reset = reset; // @[RegFile.scala 78:19:@125380.4]
  assign regs_27_io_enable = 1'h1; // @[RegFile.scala 74:20:@125374.4]
  assign regs_28_clock = clock; // @[:@125383.4]
  assign regs_28_reset = io_reset; // @[:@125384.4 RegFile.scala 76:16:@125391.4]
  assign regs_28_io_in = 64'h0; // @[RegFile.scala 75:16:@125390.4]
  assign regs_28_io_reset = reset; // @[RegFile.scala 78:19:@125394.4]
  assign regs_28_io_enable = 1'h1; // @[RegFile.scala 74:20:@125388.4]
  assign regs_29_clock = clock; // @[:@125397.4]
  assign regs_29_reset = io_reset; // @[:@125398.4 RegFile.scala 76:16:@125405.4]
  assign regs_29_io_in = 64'h0; // @[RegFile.scala 75:16:@125404.4]
  assign regs_29_io_reset = reset; // @[RegFile.scala 78:19:@125408.4]
  assign regs_29_io_enable = 1'h1; // @[RegFile.scala 74:20:@125402.4]
  assign regs_30_clock = clock; // @[:@125411.4]
  assign regs_30_reset = io_reset; // @[:@125412.4 RegFile.scala 76:16:@125419.4]
  assign regs_30_io_in = 64'h0; // @[RegFile.scala 75:16:@125418.4]
  assign regs_30_io_reset = reset; // @[RegFile.scala 78:19:@125422.4]
  assign regs_30_io_enable = 1'h1; // @[RegFile.scala 74:20:@125416.4]
  assign regs_31_clock = clock; // @[:@125425.4]
  assign regs_31_reset = io_reset; // @[:@125426.4 RegFile.scala 76:16:@125433.4]
  assign regs_31_io_in = 64'h0; // @[RegFile.scala 75:16:@125432.4]
  assign regs_31_io_reset = reset; // @[RegFile.scala 78:19:@125436.4]
  assign regs_31_io_enable = 1'h1; // @[RegFile.scala 74:20:@125430.4]
  assign regs_32_clock = clock; // @[:@125439.4]
  assign regs_32_reset = io_reset; // @[:@125440.4 RegFile.scala 76:16:@125447.4]
  assign regs_32_io_in = 64'h0; // @[RegFile.scala 75:16:@125446.4]
  assign regs_32_io_reset = reset; // @[RegFile.scala 78:19:@125450.4]
  assign regs_32_io_enable = 1'h1; // @[RegFile.scala 74:20:@125444.4]
  assign regs_33_clock = clock; // @[:@125453.4]
  assign regs_33_reset = io_reset; // @[:@125454.4 RegFile.scala 76:16:@125461.4]
  assign regs_33_io_in = 64'h0; // @[RegFile.scala 75:16:@125460.4]
  assign regs_33_io_reset = reset; // @[RegFile.scala 78:19:@125464.4]
  assign regs_33_io_enable = 1'h1; // @[RegFile.scala 74:20:@125458.4]
  assign regs_34_clock = clock; // @[:@125467.4]
  assign regs_34_reset = io_reset; // @[:@125468.4 RegFile.scala 76:16:@125475.4]
  assign regs_34_io_in = 64'h0; // @[RegFile.scala 75:16:@125474.4]
  assign regs_34_io_reset = reset; // @[RegFile.scala 78:19:@125478.4]
  assign regs_34_io_enable = 1'h1; // @[RegFile.scala 74:20:@125472.4]
  assign regs_35_clock = clock; // @[:@125481.4]
  assign regs_35_reset = io_reset; // @[:@125482.4 RegFile.scala 76:16:@125489.4]
  assign regs_35_io_in = 64'h0; // @[RegFile.scala 75:16:@125488.4]
  assign regs_35_io_reset = reset; // @[RegFile.scala 78:19:@125492.4]
  assign regs_35_io_enable = 1'h1; // @[RegFile.scala 74:20:@125486.4]
  assign regs_36_clock = clock; // @[:@125495.4]
  assign regs_36_reset = io_reset; // @[:@125496.4 RegFile.scala 76:16:@125503.4]
  assign regs_36_io_in = 64'h0; // @[RegFile.scala 75:16:@125502.4]
  assign regs_36_io_reset = reset; // @[RegFile.scala 78:19:@125506.4]
  assign regs_36_io_enable = 1'h1; // @[RegFile.scala 74:20:@125500.4]
  assign regs_37_clock = clock; // @[:@125509.4]
  assign regs_37_reset = io_reset; // @[:@125510.4 RegFile.scala 76:16:@125517.4]
  assign regs_37_io_in = 64'h0; // @[RegFile.scala 75:16:@125516.4]
  assign regs_37_io_reset = reset; // @[RegFile.scala 78:19:@125520.4]
  assign regs_37_io_enable = 1'h1; // @[RegFile.scala 74:20:@125514.4]
  assign regs_38_clock = clock; // @[:@125523.4]
  assign regs_38_reset = io_reset; // @[:@125524.4 RegFile.scala 76:16:@125531.4]
  assign regs_38_io_in = 64'h0; // @[RegFile.scala 75:16:@125530.4]
  assign regs_38_io_reset = reset; // @[RegFile.scala 78:19:@125534.4]
  assign regs_38_io_enable = 1'h1; // @[RegFile.scala 74:20:@125528.4]
  assign regs_39_clock = clock; // @[:@125537.4]
  assign regs_39_reset = io_reset; // @[:@125538.4 RegFile.scala 76:16:@125545.4]
  assign regs_39_io_in = 64'h0; // @[RegFile.scala 75:16:@125544.4]
  assign regs_39_io_reset = reset; // @[RegFile.scala 78:19:@125548.4]
  assign regs_39_io_enable = 1'h1; // @[RegFile.scala 74:20:@125542.4]
  assign regs_40_clock = clock; // @[:@125551.4]
  assign regs_40_reset = io_reset; // @[:@125552.4 RegFile.scala 76:16:@125559.4]
  assign regs_40_io_in = 64'h0; // @[RegFile.scala 75:16:@125558.4]
  assign regs_40_io_reset = reset; // @[RegFile.scala 78:19:@125562.4]
  assign regs_40_io_enable = 1'h1; // @[RegFile.scala 74:20:@125556.4]
  assign regs_41_clock = clock; // @[:@125565.4]
  assign regs_41_reset = io_reset; // @[:@125566.4 RegFile.scala 76:16:@125573.4]
  assign regs_41_io_in = 64'h0; // @[RegFile.scala 75:16:@125572.4]
  assign regs_41_io_reset = reset; // @[RegFile.scala 78:19:@125576.4]
  assign regs_41_io_enable = 1'h1; // @[RegFile.scala 74:20:@125570.4]
  assign regs_42_clock = clock; // @[:@125579.4]
  assign regs_42_reset = io_reset; // @[:@125580.4 RegFile.scala 76:16:@125587.4]
  assign regs_42_io_in = 64'h0; // @[RegFile.scala 75:16:@125586.4]
  assign regs_42_io_reset = reset; // @[RegFile.scala 78:19:@125590.4]
  assign regs_42_io_enable = 1'h1; // @[RegFile.scala 74:20:@125584.4]
  assign regs_43_clock = clock; // @[:@125593.4]
  assign regs_43_reset = io_reset; // @[:@125594.4 RegFile.scala 76:16:@125601.4]
  assign regs_43_io_in = 64'h0; // @[RegFile.scala 75:16:@125600.4]
  assign regs_43_io_reset = reset; // @[RegFile.scala 78:19:@125604.4]
  assign regs_43_io_enable = 1'h1; // @[RegFile.scala 74:20:@125598.4]
  assign regs_44_clock = clock; // @[:@125607.4]
  assign regs_44_reset = io_reset; // @[:@125608.4 RegFile.scala 76:16:@125615.4]
  assign regs_44_io_in = 64'h0; // @[RegFile.scala 75:16:@125614.4]
  assign regs_44_io_reset = reset; // @[RegFile.scala 78:19:@125618.4]
  assign regs_44_io_enable = 1'h1; // @[RegFile.scala 74:20:@125612.4]
  assign regs_45_clock = clock; // @[:@125621.4]
  assign regs_45_reset = io_reset; // @[:@125622.4 RegFile.scala 76:16:@125629.4]
  assign regs_45_io_in = 64'h0; // @[RegFile.scala 75:16:@125628.4]
  assign regs_45_io_reset = reset; // @[RegFile.scala 78:19:@125632.4]
  assign regs_45_io_enable = 1'h1; // @[RegFile.scala 74:20:@125626.4]
  assign regs_46_clock = clock; // @[:@125635.4]
  assign regs_46_reset = io_reset; // @[:@125636.4 RegFile.scala 76:16:@125643.4]
  assign regs_46_io_in = 64'h0; // @[RegFile.scala 75:16:@125642.4]
  assign regs_46_io_reset = reset; // @[RegFile.scala 78:19:@125646.4]
  assign regs_46_io_enable = 1'h1; // @[RegFile.scala 74:20:@125640.4]
  assign regs_47_clock = clock; // @[:@125649.4]
  assign regs_47_reset = io_reset; // @[:@125650.4 RegFile.scala 76:16:@125657.4]
  assign regs_47_io_in = 64'h0; // @[RegFile.scala 75:16:@125656.4]
  assign regs_47_io_reset = reset; // @[RegFile.scala 78:19:@125660.4]
  assign regs_47_io_enable = 1'h1; // @[RegFile.scala 74:20:@125654.4]
  assign regs_48_clock = clock; // @[:@125663.4]
  assign regs_48_reset = io_reset; // @[:@125664.4 RegFile.scala 76:16:@125671.4]
  assign regs_48_io_in = 64'h0; // @[RegFile.scala 75:16:@125670.4]
  assign regs_48_io_reset = reset; // @[RegFile.scala 78:19:@125674.4]
  assign regs_48_io_enable = 1'h1; // @[RegFile.scala 74:20:@125668.4]
  assign regs_49_clock = clock; // @[:@125677.4]
  assign regs_49_reset = io_reset; // @[:@125678.4 RegFile.scala 76:16:@125685.4]
  assign regs_49_io_in = 64'h0; // @[RegFile.scala 75:16:@125684.4]
  assign regs_49_io_reset = reset; // @[RegFile.scala 78:19:@125688.4]
  assign regs_49_io_enable = 1'h1; // @[RegFile.scala 74:20:@125682.4]
  assign regs_50_clock = clock; // @[:@125691.4]
  assign regs_50_reset = io_reset; // @[:@125692.4 RegFile.scala 76:16:@125699.4]
  assign regs_50_io_in = 64'h0; // @[RegFile.scala 75:16:@125698.4]
  assign regs_50_io_reset = reset; // @[RegFile.scala 78:19:@125702.4]
  assign regs_50_io_enable = 1'h1; // @[RegFile.scala 74:20:@125696.4]
  assign regs_51_clock = clock; // @[:@125705.4]
  assign regs_51_reset = io_reset; // @[:@125706.4 RegFile.scala 76:16:@125713.4]
  assign regs_51_io_in = 64'h0; // @[RegFile.scala 75:16:@125712.4]
  assign regs_51_io_reset = reset; // @[RegFile.scala 78:19:@125716.4]
  assign regs_51_io_enable = 1'h1; // @[RegFile.scala 74:20:@125710.4]
  assign regs_52_clock = clock; // @[:@125719.4]
  assign regs_52_reset = io_reset; // @[:@125720.4 RegFile.scala 76:16:@125727.4]
  assign regs_52_io_in = 64'h0; // @[RegFile.scala 75:16:@125726.4]
  assign regs_52_io_reset = reset; // @[RegFile.scala 78:19:@125730.4]
  assign regs_52_io_enable = 1'h1; // @[RegFile.scala 74:20:@125724.4]
  assign regs_53_clock = clock; // @[:@125733.4]
  assign regs_53_reset = io_reset; // @[:@125734.4 RegFile.scala 76:16:@125741.4]
  assign regs_53_io_in = 64'h0; // @[RegFile.scala 75:16:@125740.4]
  assign regs_53_io_reset = reset; // @[RegFile.scala 78:19:@125744.4]
  assign regs_53_io_enable = 1'h1; // @[RegFile.scala 74:20:@125738.4]
  assign regs_54_clock = clock; // @[:@125747.4]
  assign regs_54_reset = io_reset; // @[:@125748.4 RegFile.scala 76:16:@125755.4]
  assign regs_54_io_in = 64'h0; // @[RegFile.scala 75:16:@125754.4]
  assign regs_54_io_reset = reset; // @[RegFile.scala 78:19:@125758.4]
  assign regs_54_io_enable = 1'h1; // @[RegFile.scala 74:20:@125752.4]
  assign regs_55_clock = clock; // @[:@125761.4]
  assign regs_55_reset = io_reset; // @[:@125762.4 RegFile.scala 76:16:@125769.4]
  assign regs_55_io_in = 64'h0; // @[RegFile.scala 75:16:@125768.4]
  assign regs_55_io_reset = reset; // @[RegFile.scala 78:19:@125772.4]
  assign regs_55_io_enable = 1'h1; // @[RegFile.scala 74:20:@125766.4]
  assign regs_56_clock = clock; // @[:@125775.4]
  assign regs_56_reset = io_reset; // @[:@125776.4 RegFile.scala 76:16:@125783.4]
  assign regs_56_io_in = 64'h0; // @[RegFile.scala 75:16:@125782.4]
  assign regs_56_io_reset = reset; // @[RegFile.scala 78:19:@125786.4]
  assign regs_56_io_enable = 1'h1; // @[RegFile.scala 74:20:@125780.4]
  assign regs_57_clock = clock; // @[:@125789.4]
  assign regs_57_reset = io_reset; // @[:@125790.4 RegFile.scala 76:16:@125797.4]
  assign regs_57_io_in = 64'h0; // @[RegFile.scala 75:16:@125796.4]
  assign regs_57_io_reset = reset; // @[RegFile.scala 78:19:@125800.4]
  assign regs_57_io_enable = 1'h1; // @[RegFile.scala 74:20:@125794.4]
  assign regs_58_clock = clock; // @[:@125803.4]
  assign regs_58_reset = io_reset; // @[:@125804.4 RegFile.scala 76:16:@125811.4]
  assign regs_58_io_in = 64'h0; // @[RegFile.scala 75:16:@125810.4]
  assign regs_58_io_reset = reset; // @[RegFile.scala 78:19:@125814.4]
  assign regs_58_io_enable = 1'h1; // @[RegFile.scala 74:20:@125808.4]
  assign regs_59_clock = clock; // @[:@125817.4]
  assign regs_59_reset = io_reset; // @[:@125818.4 RegFile.scala 76:16:@125825.4]
  assign regs_59_io_in = 64'h0; // @[RegFile.scala 75:16:@125824.4]
  assign regs_59_io_reset = reset; // @[RegFile.scala 78:19:@125828.4]
  assign regs_59_io_enable = 1'h1; // @[RegFile.scala 74:20:@125822.4]
  assign regs_60_clock = clock; // @[:@125831.4]
  assign regs_60_reset = io_reset; // @[:@125832.4 RegFile.scala 76:16:@125839.4]
  assign regs_60_io_in = 64'h0; // @[RegFile.scala 75:16:@125838.4]
  assign regs_60_io_reset = reset; // @[RegFile.scala 78:19:@125842.4]
  assign regs_60_io_enable = 1'h1; // @[RegFile.scala 74:20:@125836.4]
  assign regs_61_clock = clock; // @[:@125845.4]
  assign regs_61_reset = io_reset; // @[:@125846.4 RegFile.scala 76:16:@125853.4]
  assign regs_61_io_in = 64'h0; // @[RegFile.scala 75:16:@125852.4]
  assign regs_61_io_reset = reset; // @[RegFile.scala 78:19:@125856.4]
  assign regs_61_io_enable = 1'h1; // @[RegFile.scala 74:20:@125850.4]
  assign regs_62_clock = clock; // @[:@125859.4]
  assign regs_62_reset = io_reset; // @[:@125860.4 RegFile.scala 76:16:@125867.4]
  assign regs_62_io_in = 64'h0; // @[RegFile.scala 75:16:@125866.4]
  assign regs_62_io_reset = reset; // @[RegFile.scala 78:19:@125870.4]
  assign regs_62_io_enable = 1'h1; // @[RegFile.scala 74:20:@125864.4]
  assign regs_63_clock = clock; // @[:@125873.4]
  assign regs_63_reset = io_reset; // @[:@125874.4 RegFile.scala 76:16:@125881.4]
  assign regs_63_io_in = 64'h0; // @[RegFile.scala 75:16:@125880.4]
  assign regs_63_io_reset = reset; // @[RegFile.scala 78:19:@125884.4]
  assign regs_63_io_enable = 1'h1; // @[RegFile.scala 74:20:@125878.4]
  assign regs_64_clock = clock; // @[:@125887.4]
  assign regs_64_reset = io_reset; // @[:@125888.4 RegFile.scala 76:16:@125895.4]
  assign regs_64_io_in = 64'h0; // @[RegFile.scala 75:16:@125894.4]
  assign regs_64_io_reset = reset; // @[RegFile.scala 78:19:@125898.4]
  assign regs_64_io_enable = 1'h1; // @[RegFile.scala 74:20:@125892.4]
  assign regs_65_clock = clock; // @[:@125901.4]
  assign regs_65_reset = io_reset; // @[:@125902.4 RegFile.scala 76:16:@125909.4]
  assign regs_65_io_in = 64'h0; // @[RegFile.scala 75:16:@125908.4]
  assign regs_65_io_reset = reset; // @[RegFile.scala 78:19:@125912.4]
  assign regs_65_io_enable = 1'h1; // @[RegFile.scala 74:20:@125906.4]
  assign regs_66_clock = clock; // @[:@125915.4]
  assign regs_66_reset = io_reset; // @[:@125916.4 RegFile.scala 76:16:@125923.4]
  assign regs_66_io_in = 64'h0; // @[RegFile.scala 75:16:@125922.4]
  assign regs_66_io_reset = reset; // @[RegFile.scala 78:19:@125926.4]
  assign regs_66_io_enable = 1'h1; // @[RegFile.scala 74:20:@125920.4]
  assign regs_67_clock = clock; // @[:@125929.4]
  assign regs_67_reset = io_reset; // @[:@125930.4 RegFile.scala 76:16:@125937.4]
  assign regs_67_io_in = 64'h0; // @[RegFile.scala 75:16:@125936.4]
  assign regs_67_io_reset = reset; // @[RegFile.scala 78:19:@125940.4]
  assign regs_67_io_enable = 1'h1; // @[RegFile.scala 74:20:@125934.4]
  assign regs_68_clock = clock; // @[:@125943.4]
  assign regs_68_reset = io_reset; // @[:@125944.4 RegFile.scala 76:16:@125951.4]
  assign regs_68_io_in = 64'h0; // @[RegFile.scala 75:16:@125950.4]
  assign regs_68_io_reset = reset; // @[RegFile.scala 78:19:@125954.4]
  assign regs_68_io_enable = 1'h1; // @[RegFile.scala 74:20:@125948.4]
  assign regs_69_clock = clock; // @[:@125957.4]
  assign regs_69_reset = io_reset; // @[:@125958.4 RegFile.scala 76:16:@125965.4]
  assign regs_69_io_in = 64'h0; // @[RegFile.scala 75:16:@125964.4]
  assign regs_69_io_reset = reset; // @[RegFile.scala 78:19:@125968.4]
  assign regs_69_io_enable = 1'h1; // @[RegFile.scala 74:20:@125962.4]
  assign regs_70_clock = clock; // @[:@125971.4]
  assign regs_70_reset = io_reset; // @[:@125972.4 RegFile.scala 76:16:@125979.4]
  assign regs_70_io_in = 64'h0; // @[RegFile.scala 75:16:@125978.4]
  assign regs_70_io_reset = reset; // @[RegFile.scala 78:19:@125982.4]
  assign regs_70_io_enable = 1'h1; // @[RegFile.scala 74:20:@125976.4]
  assign regs_71_clock = clock; // @[:@125985.4]
  assign regs_71_reset = io_reset; // @[:@125986.4 RegFile.scala 76:16:@125993.4]
  assign regs_71_io_in = 64'h0; // @[RegFile.scala 75:16:@125992.4]
  assign regs_71_io_reset = reset; // @[RegFile.scala 78:19:@125996.4]
  assign regs_71_io_enable = 1'h1; // @[RegFile.scala 74:20:@125990.4]
  assign regs_72_clock = clock; // @[:@125999.4]
  assign regs_72_reset = io_reset; // @[:@126000.4 RegFile.scala 76:16:@126007.4]
  assign regs_72_io_in = 64'h0; // @[RegFile.scala 75:16:@126006.4]
  assign regs_72_io_reset = reset; // @[RegFile.scala 78:19:@126010.4]
  assign regs_72_io_enable = 1'h1; // @[RegFile.scala 74:20:@126004.4]
  assign regs_73_clock = clock; // @[:@126013.4]
  assign regs_73_reset = io_reset; // @[:@126014.4 RegFile.scala 76:16:@126021.4]
  assign regs_73_io_in = 64'h0; // @[RegFile.scala 75:16:@126020.4]
  assign regs_73_io_reset = reset; // @[RegFile.scala 78:19:@126024.4]
  assign regs_73_io_enable = 1'h1; // @[RegFile.scala 74:20:@126018.4]
  assign regs_74_clock = clock; // @[:@126027.4]
  assign regs_74_reset = io_reset; // @[:@126028.4 RegFile.scala 76:16:@126035.4]
  assign regs_74_io_in = 64'h0; // @[RegFile.scala 75:16:@126034.4]
  assign regs_74_io_reset = reset; // @[RegFile.scala 78:19:@126038.4]
  assign regs_74_io_enable = 1'h1; // @[RegFile.scala 74:20:@126032.4]
  assign regs_75_clock = clock; // @[:@126041.4]
  assign regs_75_reset = io_reset; // @[:@126042.4 RegFile.scala 76:16:@126049.4]
  assign regs_75_io_in = 64'h0; // @[RegFile.scala 75:16:@126048.4]
  assign regs_75_io_reset = reset; // @[RegFile.scala 78:19:@126052.4]
  assign regs_75_io_enable = 1'h1; // @[RegFile.scala 74:20:@126046.4]
  assign regs_76_clock = clock; // @[:@126055.4]
  assign regs_76_reset = io_reset; // @[:@126056.4 RegFile.scala 76:16:@126063.4]
  assign regs_76_io_in = 64'h0; // @[RegFile.scala 75:16:@126062.4]
  assign regs_76_io_reset = reset; // @[RegFile.scala 78:19:@126066.4]
  assign regs_76_io_enable = 1'h1; // @[RegFile.scala 74:20:@126060.4]
  assign regs_77_clock = clock; // @[:@126069.4]
  assign regs_77_reset = io_reset; // @[:@126070.4 RegFile.scala 76:16:@126077.4]
  assign regs_77_io_in = 64'h0; // @[RegFile.scala 75:16:@126076.4]
  assign regs_77_io_reset = reset; // @[RegFile.scala 78:19:@126080.4]
  assign regs_77_io_enable = 1'h1; // @[RegFile.scala 74:20:@126074.4]
  assign regs_78_clock = clock; // @[:@126083.4]
  assign regs_78_reset = io_reset; // @[:@126084.4 RegFile.scala 76:16:@126091.4]
  assign regs_78_io_in = 64'h0; // @[RegFile.scala 75:16:@126090.4]
  assign regs_78_io_reset = reset; // @[RegFile.scala 78:19:@126094.4]
  assign regs_78_io_enable = 1'h1; // @[RegFile.scala 74:20:@126088.4]
  assign regs_79_clock = clock; // @[:@126097.4]
  assign regs_79_reset = io_reset; // @[:@126098.4 RegFile.scala 76:16:@126105.4]
  assign regs_79_io_in = 64'h0; // @[RegFile.scala 75:16:@126104.4]
  assign regs_79_io_reset = reset; // @[RegFile.scala 78:19:@126108.4]
  assign regs_79_io_enable = 1'h1; // @[RegFile.scala 74:20:@126102.4]
  assign regs_80_clock = clock; // @[:@126111.4]
  assign regs_80_reset = io_reset; // @[:@126112.4 RegFile.scala 76:16:@126119.4]
  assign regs_80_io_in = 64'h0; // @[RegFile.scala 75:16:@126118.4]
  assign regs_80_io_reset = reset; // @[RegFile.scala 78:19:@126122.4]
  assign regs_80_io_enable = 1'h1; // @[RegFile.scala 74:20:@126116.4]
  assign regs_81_clock = clock; // @[:@126125.4]
  assign regs_81_reset = io_reset; // @[:@126126.4 RegFile.scala 76:16:@126133.4]
  assign regs_81_io_in = 64'h0; // @[RegFile.scala 75:16:@126132.4]
  assign regs_81_io_reset = reset; // @[RegFile.scala 78:19:@126136.4]
  assign regs_81_io_enable = 1'h1; // @[RegFile.scala 74:20:@126130.4]
  assign regs_82_clock = clock; // @[:@126139.4]
  assign regs_82_reset = io_reset; // @[:@126140.4 RegFile.scala 76:16:@126147.4]
  assign regs_82_io_in = 64'h0; // @[RegFile.scala 75:16:@126146.4]
  assign regs_82_io_reset = reset; // @[RegFile.scala 78:19:@126150.4]
  assign regs_82_io_enable = 1'h1; // @[RegFile.scala 74:20:@126144.4]
  assign regs_83_clock = clock; // @[:@126153.4]
  assign regs_83_reset = io_reset; // @[:@126154.4 RegFile.scala 76:16:@126161.4]
  assign regs_83_io_in = 64'h0; // @[RegFile.scala 75:16:@126160.4]
  assign regs_83_io_reset = reset; // @[RegFile.scala 78:19:@126164.4]
  assign regs_83_io_enable = 1'h1; // @[RegFile.scala 74:20:@126158.4]
  assign regs_84_clock = clock; // @[:@126167.4]
  assign regs_84_reset = io_reset; // @[:@126168.4 RegFile.scala 76:16:@126175.4]
  assign regs_84_io_in = 64'h0; // @[RegFile.scala 75:16:@126174.4]
  assign regs_84_io_reset = reset; // @[RegFile.scala 78:19:@126178.4]
  assign regs_84_io_enable = 1'h1; // @[RegFile.scala 74:20:@126172.4]
  assign regs_85_clock = clock; // @[:@126181.4]
  assign regs_85_reset = io_reset; // @[:@126182.4 RegFile.scala 76:16:@126189.4]
  assign regs_85_io_in = 64'h0; // @[RegFile.scala 75:16:@126188.4]
  assign regs_85_io_reset = reset; // @[RegFile.scala 78:19:@126192.4]
  assign regs_85_io_enable = 1'h1; // @[RegFile.scala 74:20:@126186.4]
  assign regs_86_clock = clock; // @[:@126195.4]
  assign regs_86_reset = io_reset; // @[:@126196.4 RegFile.scala 76:16:@126203.4]
  assign regs_86_io_in = 64'h0; // @[RegFile.scala 75:16:@126202.4]
  assign regs_86_io_reset = reset; // @[RegFile.scala 78:19:@126206.4]
  assign regs_86_io_enable = 1'h1; // @[RegFile.scala 74:20:@126200.4]
  assign regs_87_clock = clock; // @[:@126209.4]
  assign regs_87_reset = io_reset; // @[:@126210.4 RegFile.scala 76:16:@126217.4]
  assign regs_87_io_in = 64'h0; // @[RegFile.scala 75:16:@126216.4]
  assign regs_87_io_reset = reset; // @[RegFile.scala 78:19:@126220.4]
  assign regs_87_io_enable = 1'h1; // @[RegFile.scala 74:20:@126214.4]
  assign regs_88_clock = clock; // @[:@126223.4]
  assign regs_88_reset = io_reset; // @[:@126224.4 RegFile.scala 76:16:@126231.4]
  assign regs_88_io_in = 64'h0; // @[RegFile.scala 75:16:@126230.4]
  assign regs_88_io_reset = reset; // @[RegFile.scala 78:19:@126234.4]
  assign regs_88_io_enable = 1'h1; // @[RegFile.scala 74:20:@126228.4]
  assign regs_89_clock = clock; // @[:@126237.4]
  assign regs_89_reset = io_reset; // @[:@126238.4 RegFile.scala 76:16:@126245.4]
  assign regs_89_io_in = 64'h0; // @[RegFile.scala 75:16:@126244.4]
  assign regs_89_io_reset = reset; // @[RegFile.scala 78:19:@126248.4]
  assign regs_89_io_enable = 1'h1; // @[RegFile.scala 74:20:@126242.4]
  assign regs_90_clock = clock; // @[:@126251.4]
  assign regs_90_reset = io_reset; // @[:@126252.4 RegFile.scala 76:16:@126259.4]
  assign regs_90_io_in = 64'h0; // @[RegFile.scala 75:16:@126258.4]
  assign regs_90_io_reset = reset; // @[RegFile.scala 78:19:@126262.4]
  assign regs_90_io_enable = 1'h1; // @[RegFile.scala 74:20:@126256.4]
  assign regs_91_clock = clock; // @[:@126265.4]
  assign regs_91_reset = io_reset; // @[:@126266.4 RegFile.scala 76:16:@126273.4]
  assign regs_91_io_in = 64'h0; // @[RegFile.scala 75:16:@126272.4]
  assign regs_91_io_reset = reset; // @[RegFile.scala 78:19:@126276.4]
  assign regs_91_io_enable = 1'h1; // @[RegFile.scala 74:20:@126270.4]
  assign regs_92_clock = clock; // @[:@126279.4]
  assign regs_92_reset = io_reset; // @[:@126280.4 RegFile.scala 76:16:@126287.4]
  assign regs_92_io_in = 64'h0; // @[RegFile.scala 75:16:@126286.4]
  assign regs_92_io_reset = reset; // @[RegFile.scala 78:19:@126290.4]
  assign regs_92_io_enable = 1'h1; // @[RegFile.scala 74:20:@126284.4]
  assign regs_93_clock = clock; // @[:@126293.4]
  assign regs_93_reset = io_reset; // @[:@126294.4 RegFile.scala 76:16:@126301.4]
  assign regs_93_io_in = 64'h0; // @[RegFile.scala 75:16:@126300.4]
  assign regs_93_io_reset = reset; // @[RegFile.scala 78:19:@126304.4]
  assign regs_93_io_enable = 1'h1; // @[RegFile.scala 74:20:@126298.4]
  assign regs_94_clock = clock; // @[:@126307.4]
  assign regs_94_reset = io_reset; // @[:@126308.4 RegFile.scala 76:16:@126315.4]
  assign regs_94_io_in = 64'h0; // @[RegFile.scala 75:16:@126314.4]
  assign regs_94_io_reset = reset; // @[RegFile.scala 78:19:@126318.4]
  assign regs_94_io_enable = 1'h1; // @[RegFile.scala 74:20:@126312.4]
  assign regs_95_clock = clock; // @[:@126321.4]
  assign regs_95_reset = io_reset; // @[:@126322.4 RegFile.scala 76:16:@126329.4]
  assign regs_95_io_in = 64'h0; // @[RegFile.scala 75:16:@126328.4]
  assign regs_95_io_reset = reset; // @[RegFile.scala 78:19:@126332.4]
  assign regs_95_io_enable = 1'h1; // @[RegFile.scala 74:20:@126326.4]
  assign regs_96_clock = clock; // @[:@126335.4]
  assign regs_96_reset = io_reset; // @[:@126336.4 RegFile.scala 76:16:@126343.4]
  assign regs_96_io_in = 64'h0; // @[RegFile.scala 75:16:@126342.4]
  assign regs_96_io_reset = reset; // @[RegFile.scala 78:19:@126346.4]
  assign regs_96_io_enable = 1'h1; // @[RegFile.scala 74:20:@126340.4]
  assign regs_97_clock = clock; // @[:@126349.4]
  assign regs_97_reset = io_reset; // @[:@126350.4 RegFile.scala 76:16:@126357.4]
  assign regs_97_io_in = 64'h0; // @[RegFile.scala 75:16:@126356.4]
  assign regs_97_io_reset = reset; // @[RegFile.scala 78:19:@126360.4]
  assign regs_97_io_enable = 1'h1; // @[RegFile.scala 74:20:@126354.4]
  assign regs_98_clock = clock; // @[:@126363.4]
  assign regs_98_reset = io_reset; // @[:@126364.4 RegFile.scala 76:16:@126371.4]
  assign regs_98_io_in = 64'h0; // @[RegFile.scala 75:16:@126370.4]
  assign regs_98_io_reset = reset; // @[RegFile.scala 78:19:@126374.4]
  assign regs_98_io_enable = 1'h1; // @[RegFile.scala 74:20:@126368.4]
  assign regs_99_clock = clock; // @[:@126377.4]
  assign regs_99_reset = io_reset; // @[:@126378.4 RegFile.scala 76:16:@126385.4]
  assign regs_99_io_in = 64'h0; // @[RegFile.scala 75:16:@126384.4]
  assign regs_99_io_reset = reset; // @[RegFile.scala 78:19:@126388.4]
  assign regs_99_io_enable = 1'h1; // @[RegFile.scala 74:20:@126382.4]
  assign regs_100_clock = clock; // @[:@126391.4]
  assign regs_100_reset = io_reset; // @[:@126392.4 RegFile.scala 76:16:@126399.4]
  assign regs_100_io_in = 64'h0; // @[RegFile.scala 75:16:@126398.4]
  assign regs_100_io_reset = reset; // @[RegFile.scala 78:19:@126402.4]
  assign regs_100_io_enable = 1'h1; // @[RegFile.scala 74:20:@126396.4]
  assign regs_101_clock = clock; // @[:@126405.4]
  assign regs_101_reset = io_reset; // @[:@126406.4 RegFile.scala 76:16:@126413.4]
  assign regs_101_io_in = 64'h0; // @[RegFile.scala 75:16:@126412.4]
  assign regs_101_io_reset = reset; // @[RegFile.scala 78:19:@126416.4]
  assign regs_101_io_enable = 1'h1; // @[RegFile.scala 74:20:@126410.4]
  assign regs_102_clock = clock; // @[:@126419.4]
  assign regs_102_reset = io_reset; // @[:@126420.4 RegFile.scala 76:16:@126427.4]
  assign regs_102_io_in = 64'h0; // @[RegFile.scala 75:16:@126426.4]
  assign regs_102_io_reset = reset; // @[RegFile.scala 78:19:@126430.4]
  assign regs_102_io_enable = 1'h1; // @[RegFile.scala 74:20:@126424.4]
  assign regs_103_clock = clock; // @[:@126433.4]
  assign regs_103_reset = io_reset; // @[:@126434.4 RegFile.scala 76:16:@126441.4]
  assign regs_103_io_in = 64'h0; // @[RegFile.scala 75:16:@126440.4]
  assign regs_103_io_reset = reset; // @[RegFile.scala 78:19:@126444.4]
  assign regs_103_io_enable = 1'h1; // @[RegFile.scala 74:20:@126438.4]
  assign regs_104_clock = clock; // @[:@126447.4]
  assign regs_104_reset = io_reset; // @[:@126448.4 RegFile.scala 76:16:@126455.4]
  assign regs_104_io_in = 64'h0; // @[RegFile.scala 75:16:@126454.4]
  assign regs_104_io_reset = reset; // @[RegFile.scala 78:19:@126458.4]
  assign regs_104_io_enable = 1'h1; // @[RegFile.scala 74:20:@126452.4]
  assign regs_105_clock = clock; // @[:@126461.4]
  assign regs_105_reset = io_reset; // @[:@126462.4 RegFile.scala 76:16:@126469.4]
  assign regs_105_io_in = 64'h0; // @[RegFile.scala 75:16:@126468.4]
  assign regs_105_io_reset = reset; // @[RegFile.scala 78:19:@126472.4]
  assign regs_105_io_enable = 1'h1; // @[RegFile.scala 74:20:@126466.4]
  assign regs_106_clock = clock; // @[:@126475.4]
  assign regs_106_reset = io_reset; // @[:@126476.4 RegFile.scala 76:16:@126483.4]
  assign regs_106_io_in = 64'h0; // @[RegFile.scala 75:16:@126482.4]
  assign regs_106_io_reset = reset; // @[RegFile.scala 78:19:@126486.4]
  assign regs_106_io_enable = 1'h1; // @[RegFile.scala 74:20:@126480.4]
  assign regs_107_clock = clock; // @[:@126489.4]
  assign regs_107_reset = io_reset; // @[:@126490.4 RegFile.scala 76:16:@126497.4]
  assign regs_107_io_in = 64'h0; // @[RegFile.scala 75:16:@126496.4]
  assign regs_107_io_reset = reset; // @[RegFile.scala 78:19:@126500.4]
  assign regs_107_io_enable = 1'h1; // @[RegFile.scala 74:20:@126494.4]
  assign regs_108_clock = clock; // @[:@126503.4]
  assign regs_108_reset = io_reset; // @[:@126504.4 RegFile.scala 76:16:@126511.4]
  assign regs_108_io_in = 64'h0; // @[RegFile.scala 75:16:@126510.4]
  assign regs_108_io_reset = reset; // @[RegFile.scala 78:19:@126514.4]
  assign regs_108_io_enable = 1'h1; // @[RegFile.scala 74:20:@126508.4]
  assign regs_109_clock = clock; // @[:@126517.4]
  assign regs_109_reset = io_reset; // @[:@126518.4 RegFile.scala 76:16:@126525.4]
  assign regs_109_io_in = 64'h0; // @[RegFile.scala 75:16:@126524.4]
  assign regs_109_io_reset = reset; // @[RegFile.scala 78:19:@126528.4]
  assign regs_109_io_enable = 1'h1; // @[RegFile.scala 74:20:@126522.4]
  assign regs_110_clock = clock; // @[:@126531.4]
  assign regs_110_reset = io_reset; // @[:@126532.4 RegFile.scala 76:16:@126539.4]
  assign regs_110_io_in = 64'h0; // @[RegFile.scala 75:16:@126538.4]
  assign regs_110_io_reset = reset; // @[RegFile.scala 78:19:@126542.4]
  assign regs_110_io_enable = 1'h1; // @[RegFile.scala 74:20:@126536.4]
  assign regs_111_clock = clock; // @[:@126545.4]
  assign regs_111_reset = io_reset; // @[:@126546.4 RegFile.scala 76:16:@126553.4]
  assign regs_111_io_in = 64'h0; // @[RegFile.scala 75:16:@126552.4]
  assign regs_111_io_reset = reset; // @[RegFile.scala 78:19:@126556.4]
  assign regs_111_io_enable = 1'h1; // @[RegFile.scala 74:20:@126550.4]
  assign regs_112_clock = clock; // @[:@126559.4]
  assign regs_112_reset = io_reset; // @[:@126560.4 RegFile.scala 76:16:@126567.4]
  assign regs_112_io_in = 64'h0; // @[RegFile.scala 75:16:@126566.4]
  assign regs_112_io_reset = reset; // @[RegFile.scala 78:19:@126570.4]
  assign regs_112_io_enable = 1'h1; // @[RegFile.scala 74:20:@126564.4]
  assign regs_113_clock = clock; // @[:@126573.4]
  assign regs_113_reset = io_reset; // @[:@126574.4 RegFile.scala 76:16:@126581.4]
  assign regs_113_io_in = 64'h0; // @[RegFile.scala 75:16:@126580.4]
  assign regs_113_io_reset = reset; // @[RegFile.scala 78:19:@126584.4]
  assign regs_113_io_enable = 1'h1; // @[RegFile.scala 74:20:@126578.4]
  assign regs_114_clock = clock; // @[:@126587.4]
  assign regs_114_reset = io_reset; // @[:@126588.4 RegFile.scala 76:16:@126595.4]
  assign regs_114_io_in = 64'h0; // @[RegFile.scala 75:16:@126594.4]
  assign regs_114_io_reset = reset; // @[RegFile.scala 78:19:@126598.4]
  assign regs_114_io_enable = 1'h1; // @[RegFile.scala 74:20:@126592.4]
  assign regs_115_clock = clock; // @[:@126601.4]
  assign regs_115_reset = io_reset; // @[:@126602.4 RegFile.scala 76:16:@126609.4]
  assign regs_115_io_in = 64'h0; // @[RegFile.scala 75:16:@126608.4]
  assign regs_115_io_reset = reset; // @[RegFile.scala 78:19:@126612.4]
  assign regs_115_io_enable = 1'h1; // @[RegFile.scala 74:20:@126606.4]
  assign regs_116_clock = clock; // @[:@126615.4]
  assign regs_116_reset = io_reset; // @[:@126616.4 RegFile.scala 76:16:@126623.4]
  assign regs_116_io_in = 64'h0; // @[RegFile.scala 75:16:@126622.4]
  assign regs_116_io_reset = reset; // @[RegFile.scala 78:19:@126626.4]
  assign regs_116_io_enable = 1'h1; // @[RegFile.scala 74:20:@126620.4]
  assign regs_117_clock = clock; // @[:@126629.4]
  assign regs_117_reset = io_reset; // @[:@126630.4 RegFile.scala 76:16:@126637.4]
  assign regs_117_io_in = 64'h0; // @[RegFile.scala 75:16:@126636.4]
  assign regs_117_io_reset = reset; // @[RegFile.scala 78:19:@126640.4]
  assign regs_117_io_enable = 1'h1; // @[RegFile.scala 74:20:@126634.4]
  assign regs_118_clock = clock; // @[:@126643.4]
  assign regs_118_reset = io_reset; // @[:@126644.4 RegFile.scala 76:16:@126651.4]
  assign regs_118_io_in = 64'h0; // @[RegFile.scala 75:16:@126650.4]
  assign regs_118_io_reset = reset; // @[RegFile.scala 78:19:@126654.4]
  assign regs_118_io_enable = 1'h1; // @[RegFile.scala 74:20:@126648.4]
  assign regs_119_clock = clock; // @[:@126657.4]
  assign regs_119_reset = io_reset; // @[:@126658.4 RegFile.scala 76:16:@126665.4]
  assign regs_119_io_in = 64'h0; // @[RegFile.scala 75:16:@126664.4]
  assign regs_119_io_reset = reset; // @[RegFile.scala 78:19:@126668.4]
  assign regs_119_io_enable = 1'h1; // @[RegFile.scala 74:20:@126662.4]
  assign regs_120_clock = clock; // @[:@126671.4]
  assign regs_120_reset = io_reset; // @[:@126672.4 RegFile.scala 76:16:@126679.4]
  assign regs_120_io_in = 64'h0; // @[RegFile.scala 75:16:@126678.4]
  assign regs_120_io_reset = reset; // @[RegFile.scala 78:19:@126682.4]
  assign regs_120_io_enable = 1'h1; // @[RegFile.scala 74:20:@126676.4]
  assign regs_121_clock = clock; // @[:@126685.4]
  assign regs_121_reset = io_reset; // @[:@126686.4 RegFile.scala 76:16:@126693.4]
  assign regs_121_io_in = 64'h0; // @[RegFile.scala 75:16:@126692.4]
  assign regs_121_io_reset = reset; // @[RegFile.scala 78:19:@126696.4]
  assign regs_121_io_enable = 1'h1; // @[RegFile.scala 74:20:@126690.4]
  assign regs_122_clock = clock; // @[:@126699.4]
  assign regs_122_reset = io_reset; // @[:@126700.4 RegFile.scala 76:16:@126707.4]
  assign regs_122_io_in = 64'h0; // @[RegFile.scala 75:16:@126706.4]
  assign regs_122_io_reset = reset; // @[RegFile.scala 78:19:@126710.4]
  assign regs_122_io_enable = 1'h1; // @[RegFile.scala 74:20:@126704.4]
  assign regs_123_clock = clock; // @[:@126713.4]
  assign regs_123_reset = io_reset; // @[:@126714.4 RegFile.scala 76:16:@126721.4]
  assign regs_123_io_in = 64'h0; // @[RegFile.scala 75:16:@126720.4]
  assign regs_123_io_reset = reset; // @[RegFile.scala 78:19:@126724.4]
  assign regs_123_io_enable = 1'h1; // @[RegFile.scala 74:20:@126718.4]
  assign regs_124_clock = clock; // @[:@126727.4]
  assign regs_124_reset = io_reset; // @[:@126728.4 RegFile.scala 76:16:@126735.4]
  assign regs_124_io_in = 64'h0; // @[RegFile.scala 75:16:@126734.4]
  assign regs_124_io_reset = reset; // @[RegFile.scala 78:19:@126738.4]
  assign regs_124_io_enable = 1'h1; // @[RegFile.scala 74:20:@126732.4]
  assign regs_125_clock = clock; // @[:@126741.4]
  assign regs_125_reset = io_reset; // @[:@126742.4 RegFile.scala 76:16:@126749.4]
  assign regs_125_io_in = 64'h0; // @[RegFile.scala 75:16:@126748.4]
  assign regs_125_io_reset = reset; // @[RegFile.scala 78:19:@126752.4]
  assign regs_125_io_enable = 1'h1; // @[RegFile.scala 74:20:@126746.4]
  assign regs_126_clock = clock; // @[:@126755.4]
  assign regs_126_reset = io_reset; // @[:@126756.4 RegFile.scala 76:16:@126763.4]
  assign regs_126_io_in = 64'h0; // @[RegFile.scala 75:16:@126762.4]
  assign regs_126_io_reset = reset; // @[RegFile.scala 78:19:@126766.4]
  assign regs_126_io_enable = 1'h1; // @[RegFile.scala 74:20:@126760.4]
  assign regs_127_clock = clock; // @[:@126769.4]
  assign regs_127_reset = io_reset; // @[:@126770.4 RegFile.scala 76:16:@126777.4]
  assign regs_127_io_in = 64'h0; // @[RegFile.scala 75:16:@126776.4]
  assign regs_127_io_reset = reset; // @[RegFile.scala 78:19:@126780.4]
  assign regs_127_io_enable = 1'h1; // @[RegFile.scala 74:20:@126774.4]
  assign regs_128_clock = clock; // @[:@126783.4]
  assign regs_128_reset = io_reset; // @[:@126784.4 RegFile.scala 76:16:@126791.4]
  assign regs_128_io_in = 64'h0; // @[RegFile.scala 75:16:@126790.4]
  assign regs_128_io_reset = reset; // @[RegFile.scala 78:19:@126794.4]
  assign regs_128_io_enable = 1'h1; // @[RegFile.scala 74:20:@126788.4]
  assign regs_129_clock = clock; // @[:@126797.4]
  assign regs_129_reset = io_reset; // @[:@126798.4 RegFile.scala 76:16:@126805.4]
  assign regs_129_io_in = 64'h0; // @[RegFile.scala 75:16:@126804.4]
  assign regs_129_io_reset = reset; // @[RegFile.scala 78:19:@126808.4]
  assign regs_129_io_enable = 1'h1; // @[RegFile.scala 74:20:@126802.4]
  assign regs_130_clock = clock; // @[:@126811.4]
  assign regs_130_reset = io_reset; // @[:@126812.4 RegFile.scala 76:16:@126819.4]
  assign regs_130_io_in = 64'h0; // @[RegFile.scala 75:16:@126818.4]
  assign regs_130_io_reset = reset; // @[RegFile.scala 78:19:@126822.4]
  assign regs_130_io_enable = 1'h1; // @[RegFile.scala 74:20:@126816.4]
  assign regs_131_clock = clock; // @[:@126825.4]
  assign regs_131_reset = io_reset; // @[:@126826.4 RegFile.scala 76:16:@126833.4]
  assign regs_131_io_in = 64'h0; // @[RegFile.scala 75:16:@126832.4]
  assign regs_131_io_reset = reset; // @[RegFile.scala 78:19:@126836.4]
  assign regs_131_io_enable = 1'h1; // @[RegFile.scala 74:20:@126830.4]
  assign regs_132_clock = clock; // @[:@126839.4]
  assign regs_132_reset = io_reset; // @[:@126840.4 RegFile.scala 76:16:@126847.4]
  assign regs_132_io_in = 64'h0; // @[RegFile.scala 75:16:@126846.4]
  assign regs_132_io_reset = reset; // @[RegFile.scala 78:19:@126850.4]
  assign regs_132_io_enable = 1'h1; // @[RegFile.scala 74:20:@126844.4]
  assign regs_133_clock = clock; // @[:@126853.4]
  assign regs_133_reset = io_reset; // @[:@126854.4 RegFile.scala 76:16:@126861.4]
  assign regs_133_io_in = 64'h0; // @[RegFile.scala 75:16:@126860.4]
  assign regs_133_io_reset = reset; // @[RegFile.scala 78:19:@126864.4]
  assign regs_133_io_enable = 1'h1; // @[RegFile.scala 74:20:@126858.4]
  assign regs_134_clock = clock; // @[:@126867.4]
  assign regs_134_reset = io_reset; // @[:@126868.4 RegFile.scala 76:16:@126875.4]
  assign regs_134_io_in = 64'h0; // @[RegFile.scala 75:16:@126874.4]
  assign regs_134_io_reset = reset; // @[RegFile.scala 78:19:@126878.4]
  assign regs_134_io_enable = 1'h1; // @[RegFile.scala 74:20:@126872.4]
  assign regs_135_clock = clock; // @[:@126881.4]
  assign regs_135_reset = io_reset; // @[:@126882.4 RegFile.scala 76:16:@126889.4]
  assign regs_135_io_in = 64'h0; // @[RegFile.scala 75:16:@126888.4]
  assign regs_135_io_reset = reset; // @[RegFile.scala 78:19:@126892.4]
  assign regs_135_io_enable = 1'h1; // @[RegFile.scala 74:20:@126886.4]
  assign regs_136_clock = clock; // @[:@126895.4]
  assign regs_136_reset = io_reset; // @[:@126896.4 RegFile.scala 76:16:@126903.4]
  assign regs_136_io_in = 64'h0; // @[RegFile.scala 75:16:@126902.4]
  assign regs_136_io_reset = reset; // @[RegFile.scala 78:19:@126906.4]
  assign regs_136_io_enable = 1'h1; // @[RegFile.scala 74:20:@126900.4]
  assign regs_137_clock = clock; // @[:@126909.4]
  assign regs_137_reset = io_reset; // @[:@126910.4 RegFile.scala 76:16:@126917.4]
  assign regs_137_io_in = 64'h0; // @[RegFile.scala 75:16:@126916.4]
  assign regs_137_io_reset = reset; // @[RegFile.scala 78:19:@126920.4]
  assign regs_137_io_enable = 1'h1; // @[RegFile.scala 74:20:@126914.4]
  assign regs_138_clock = clock; // @[:@126923.4]
  assign regs_138_reset = io_reset; // @[:@126924.4 RegFile.scala 76:16:@126931.4]
  assign regs_138_io_in = 64'h0; // @[RegFile.scala 75:16:@126930.4]
  assign regs_138_io_reset = reset; // @[RegFile.scala 78:19:@126934.4]
  assign regs_138_io_enable = 1'h1; // @[RegFile.scala 74:20:@126928.4]
  assign regs_139_clock = clock; // @[:@126937.4]
  assign regs_139_reset = io_reset; // @[:@126938.4 RegFile.scala 76:16:@126945.4]
  assign regs_139_io_in = 64'h0; // @[RegFile.scala 75:16:@126944.4]
  assign regs_139_io_reset = reset; // @[RegFile.scala 78:19:@126948.4]
  assign regs_139_io_enable = 1'h1; // @[RegFile.scala 74:20:@126942.4]
  assign regs_140_clock = clock; // @[:@126951.4]
  assign regs_140_reset = io_reset; // @[:@126952.4 RegFile.scala 76:16:@126959.4]
  assign regs_140_io_in = 64'h0; // @[RegFile.scala 75:16:@126958.4]
  assign regs_140_io_reset = reset; // @[RegFile.scala 78:19:@126962.4]
  assign regs_140_io_enable = 1'h1; // @[RegFile.scala 74:20:@126956.4]
  assign regs_141_clock = clock; // @[:@126965.4]
  assign regs_141_reset = io_reset; // @[:@126966.4 RegFile.scala 76:16:@126973.4]
  assign regs_141_io_in = 64'h0; // @[RegFile.scala 75:16:@126972.4]
  assign regs_141_io_reset = reset; // @[RegFile.scala 78:19:@126976.4]
  assign regs_141_io_enable = 1'h1; // @[RegFile.scala 74:20:@126970.4]
  assign regs_142_clock = clock; // @[:@126979.4]
  assign regs_142_reset = io_reset; // @[:@126980.4 RegFile.scala 76:16:@126987.4]
  assign regs_142_io_in = 64'h0; // @[RegFile.scala 75:16:@126986.4]
  assign regs_142_io_reset = reset; // @[RegFile.scala 78:19:@126990.4]
  assign regs_142_io_enable = 1'h1; // @[RegFile.scala 74:20:@126984.4]
  assign regs_143_clock = clock; // @[:@126993.4]
  assign regs_143_reset = io_reset; // @[:@126994.4 RegFile.scala 76:16:@127001.4]
  assign regs_143_io_in = 64'h0; // @[RegFile.scala 75:16:@127000.4]
  assign regs_143_io_reset = reset; // @[RegFile.scala 78:19:@127004.4]
  assign regs_143_io_enable = 1'h1; // @[RegFile.scala 74:20:@126998.4]
  assign regs_144_clock = clock; // @[:@127007.4]
  assign regs_144_reset = io_reset; // @[:@127008.4 RegFile.scala 76:16:@127015.4]
  assign regs_144_io_in = 64'h0; // @[RegFile.scala 75:16:@127014.4]
  assign regs_144_io_reset = reset; // @[RegFile.scala 78:19:@127018.4]
  assign regs_144_io_enable = 1'h1; // @[RegFile.scala 74:20:@127012.4]
  assign regs_145_clock = clock; // @[:@127021.4]
  assign regs_145_reset = io_reset; // @[:@127022.4 RegFile.scala 76:16:@127029.4]
  assign regs_145_io_in = 64'h0; // @[RegFile.scala 75:16:@127028.4]
  assign regs_145_io_reset = reset; // @[RegFile.scala 78:19:@127032.4]
  assign regs_145_io_enable = 1'h1; // @[RegFile.scala 74:20:@127026.4]
  assign regs_146_clock = clock; // @[:@127035.4]
  assign regs_146_reset = io_reset; // @[:@127036.4 RegFile.scala 76:16:@127043.4]
  assign regs_146_io_in = 64'h0; // @[RegFile.scala 75:16:@127042.4]
  assign regs_146_io_reset = reset; // @[RegFile.scala 78:19:@127046.4]
  assign regs_146_io_enable = 1'h1; // @[RegFile.scala 74:20:@127040.4]
  assign regs_147_clock = clock; // @[:@127049.4]
  assign regs_147_reset = io_reset; // @[:@127050.4 RegFile.scala 76:16:@127057.4]
  assign regs_147_io_in = 64'h0; // @[RegFile.scala 75:16:@127056.4]
  assign regs_147_io_reset = reset; // @[RegFile.scala 78:19:@127060.4]
  assign regs_147_io_enable = 1'h1; // @[RegFile.scala 74:20:@127054.4]
  assign regs_148_clock = clock; // @[:@127063.4]
  assign regs_148_reset = io_reset; // @[:@127064.4 RegFile.scala 76:16:@127071.4]
  assign regs_148_io_in = 64'h0; // @[RegFile.scala 75:16:@127070.4]
  assign regs_148_io_reset = reset; // @[RegFile.scala 78:19:@127074.4]
  assign regs_148_io_enable = 1'h1; // @[RegFile.scala 74:20:@127068.4]
  assign regs_149_clock = clock; // @[:@127077.4]
  assign regs_149_reset = io_reset; // @[:@127078.4 RegFile.scala 76:16:@127085.4]
  assign regs_149_io_in = 64'h0; // @[RegFile.scala 75:16:@127084.4]
  assign regs_149_io_reset = reset; // @[RegFile.scala 78:19:@127088.4]
  assign regs_149_io_enable = 1'h1; // @[RegFile.scala 74:20:@127082.4]
  assign regs_150_clock = clock; // @[:@127091.4]
  assign regs_150_reset = io_reset; // @[:@127092.4 RegFile.scala 76:16:@127099.4]
  assign regs_150_io_in = 64'h0; // @[RegFile.scala 75:16:@127098.4]
  assign regs_150_io_reset = reset; // @[RegFile.scala 78:19:@127102.4]
  assign regs_150_io_enable = 1'h1; // @[RegFile.scala 74:20:@127096.4]
  assign regs_151_clock = clock; // @[:@127105.4]
  assign regs_151_reset = io_reset; // @[:@127106.4 RegFile.scala 76:16:@127113.4]
  assign regs_151_io_in = 64'h0; // @[RegFile.scala 75:16:@127112.4]
  assign regs_151_io_reset = reset; // @[RegFile.scala 78:19:@127116.4]
  assign regs_151_io_enable = 1'h1; // @[RegFile.scala 74:20:@127110.4]
  assign regs_152_clock = clock; // @[:@127119.4]
  assign regs_152_reset = io_reset; // @[:@127120.4 RegFile.scala 76:16:@127127.4]
  assign regs_152_io_in = 64'h0; // @[RegFile.scala 75:16:@127126.4]
  assign regs_152_io_reset = reset; // @[RegFile.scala 78:19:@127130.4]
  assign regs_152_io_enable = 1'h1; // @[RegFile.scala 74:20:@127124.4]
  assign regs_153_clock = clock; // @[:@127133.4]
  assign regs_153_reset = io_reset; // @[:@127134.4 RegFile.scala 76:16:@127141.4]
  assign regs_153_io_in = 64'h0; // @[RegFile.scala 75:16:@127140.4]
  assign regs_153_io_reset = reset; // @[RegFile.scala 78:19:@127144.4]
  assign regs_153_io_enable = 1'h1; // @[RegFile.scala 74:20:@127138.4]
  assign regs_154_clock = clock; // @[:@127147.4]
  assign regs_154_reset = io_reset; // @[:@127148.4 RegFile.scala 76:16:@127155.4]
  assign regs_154_io_in = 64'h0; // @[RegFile.scala 75:16:@127154.4]
  assign regs_154_io_reset = reset; // @[RegFile.scala 78:19:@127158.4]
  assign regs_154_io_enable = 1'h1; // @[RegFile.scala 74:20:@127152.4]
  assign regs_155_clock = clock; // @[:@127161.4]
  assign regs_155_reset = io_reset; // @[:@127162.4 RegFile.scala 76:16:@127169.4]
  assign regs_155_io_in = 64'h0; // @[RegFile.scala 75:16:@127168.4]
  assign regs_155_io_reset = reset; // @[RegFile.scala 78:19:@127172.4]
  assign regs_155_io_enable = 1'h1; // @[RegFile.scala 74:20:@127166.4]
  assign regs_156_clock = clock; // @[:@127175.4]
  assign regs_156_reset = io_reset; // @[:@127176.4 RegFile.scala 76:16:@127183.4]
  assign regs_156_io_in = 64'h0; // @[RegFile.scala 75:16:@127182.4]
  assign regs_156_io_reset = reset; // @[RegFile.scala 78:19:@127186.4]
  assign regs_156_io_enable = 1'h1; // @[RegFile.scala 74:20:@127180.4]
  assign regs_157_clock = clock; // @[:@127189.4]
  assign regs_157_reset = io_reset; // @[:@127190.4 RegFile.scala 76:16:@127197.4]
  assign regs_157_io_in = 64'h0; // @[RegFile.scala 75:16:@127196.4]
  assign regs_157_io_reset = reset; // @[RegFile.scala 78:19:@127200.4]
  assign regs_157_io_enable = 1'h1; // @[RegFile.scala 74:20:@127194.4]
  assign regs_158_clock = clock; // @[:@127203.4]
  assign regs_158_reset = io_reset; // @[:@127204.4 RegFile.scala 76:16:@127211.4]
  assign regs_158_io_in = 64'h0; // @[RegFile.scala 75:16:@127210.4]
  assign regs_158_io_reset = reset; // @[RegFile.scala 78:19:@127214.4]
  assign regs_158_io_enable = 1'h1; // @[RegFile.scala 74:20:@127208.4]
  assign regs_159_clock = clock; // @[:@127217.4]
  assign regs_159_reset = io_reset; // @[:@127218.4 RegFile.scala 76:16:@127225.4]
  assign regs_159_io_in = 64'h0; // @[RegFile.scala 75:16:@127224.4]
  assign regs_159_io_reset = reset; // @[RegFile.scala 78:19:@127228.4]
  assign regs_159_io_enable = 1'h1; // @[RegFile.scala 74:20:@127222.4]
  assign regs_160_clock = clock; // @[:@127231.4]
  assign regs_160_reset = io_reset; // @[:@127232.4 RegFile.scala 76:16:@127239.4]
  assign regs_160_io_in = 64'h0; // @[RegFile.scala 75:16:@127238.4]
  assign regs_160_io_reset = reset; // @[RegFile.scala 78:19:@127242.4]
  assign regs_160_io_enable = 1'h1; // @[RegFile.scala 74:20:@127236.4]
  assign regs_161_clock = clock; // @[:@127245.4]
  assign regs_161_reset = io_reset; // @[:@127246.4 RegFile.scala 76:16:@127253.4]
  assign regs_161_io_in = 64'h0; // @[RegFile.scala 75:16:@127252.4]
  assign regs_161_io_reset = reset; // @[RegFile.scala 78:19:@127256.4]
  assign regs_161_io_enable = 1'h1; // @[RegFile.scala 74:20:@127250.4]
  assign regs_162_clock = clock; // @[:@127259.4]
  assign regs_162_reset = io_reset; // @[:@127260.4 RegFile.scala 76:16:@127267.4]
  assign regs_162_io_in = 64'h0; // @[RegFile.scala 75:16:@127266.4]
  assign regs_162_io_reset = reset; // @[RegFile.scala 78:19:@127270.4]
  assign regs_162_io_enable = 1'h1; // @[RegFile.scala 74:20:@127264.4]
  assign regs_163_clock = clock; // @[:@127273.4]
  assign regs_163_reset = io_reset; // @[:@127274.4 RegFile.scala 76:16:@127281.4]
  assign regs_163_io_in = 64'h0; // @[RegFile.scala 75:16:@127280.4]
  assign regs_163_io_reset = reset; // @[RegFile.scala 78:19:@127284.4]
  assign regs_163_io_enable = 1'h1; // @[RegFile.scala 74:20:@127278.4]
  assign regs_164_clock = clock; // @[:@127287.4]
  assign regs_164_reset = io_reset; // @[:@127288.4 RegFile.scala 76:16:@127295.4]
  assign regs_164_io_in = 64'h0; // @[RegFile.scala 75:16:@127294.4]
  assign regs_164_io_reset = reset; // @[RegFile.scala 78:19:@127298.4]
  assign regs_164_io_enable = 1'h1; // @[RegFile.scala 74:20:@127292.4]
  assign regs_165_clock = clock; // @[:@127301.4]
  assign regs_165_reset = io_reset; // @[:@127302.4 RegFile.scala 76:16:@127309.4]
  assign regs_165_io_in = 64'h0; // @[RegFile.scala 75:16:@127308.4]
  assign regs_165_io_reset = reset; // @[RegFile.scala 78:19:@127312.4]
  assign regs_165_io_enable = 1'h1; // @[RegFile.scala 74:20:@127306.4]
  assign regs_166_clock = clock; // @[:@127315.4]
  assign regs_166_reset = io_reset; // @[:@127316.4 RegFile.scala 76:16:@127323.4]
  assign regs_166_io_in = 64'h0; // @[RegFile.scala 75:16:@127322.4]
  assign regs_166_io_reset = reset; // @[RegFile.scala 78:19:@127326.4]
  assign regs_166_io_enable = 1'h1; // @[RegFile.scala 74:20:@127320.4]
  assign regs_167_clock = clock; // @[:@127329.4]
  assign regs_167_reset = io_reset; // @[:@127330.4 RegFile.scala 76:16:@127337.4]
  assign regs_167_io_in = 64'h0; // @[RegFile.scala 75:16:@127336.4]
  assign regs_167_io_reset = reset; // @[RegFile.scala 78:19:@127340.4]
  assign regs_167_io_enable = 1'h1; // @[RegFile.scala 74:20:@127334.4]
  assign regs_168_clock = clock; // @[:@127343.4]
  assign regs_168_reset = io_reset; // @[:@127344.4 RegFile.scala 76:16:@127351.4]
  assign regs_168_io_in = 64'h0; // @[RegFile.scala 75:16:@127350.4]
  assign regs_168_io_reset = reset; // @[RegFile.scala 78:19:@127354.4]
  assign regs_168_io_enable = 1'h1; // @[RegFile.scala 74:20:@127348.4]
  assign regs_169_clock = clock; // @[:@127357.4]
  assign regs_169_reset = io_reset; // @[:@127358.4 RegFile.scala 76:16:@127365.4]
  assign regs_169_io_in = 64'h0; // @[RegFile.scala 75:16:@127364.4]
  assign regs_169_io_reset = reset; // @[RegFile.scala 78:19:@127368.4]
  assign regs_169_io_enable = 1'h1; // @[RegFile.scala 74:20:@127362.4]
  assign regs_170_clock = clock; // @[:@127371.4]
  assign regs_170_reset = io_reset; // @[:@127372.4 RegFile.scala 76:16:@127379.4]
  assign regs_170_io_in = 64'h0; // @[RegFile.scala 75:16:@127378.4]
  assign regs_170_io_reset = reset; // @[RegFile.scala 78:19:@127382.4]
  assign regs_170_io_enable = 1'h1; // @[RegFile.scala 74:20:@127376.4]
  assign regs_171_clock = clock; // @[:@127385.4]
  assign regs_171_reset = io_reset; // @[:@127386.4 RegFile.scala 76:16:@127393.4]
  assign regs_171_io_in = 64'h0; // @[RegFile.scala 75:16:@127392.4]
  assign regs_171_io_reset = reset; // @[RegFile.scala 78:19:@127396.4]
  assign regs_171_io_enable = 1'h1; // @[RegFile.scala 74:20:@127390.4]
  assign regs_172_clock = clock; // @[:@127399.4]
  assign regs_172_reset = io_reset; // @[:@127400.4 RegFile.scala 76:16:@127407.4]
  assign regs_172_io_in = 64'h0; // @[RegFile.scala 75:16:@127406.4]
  assign regs_172_io_reset = reset; // @[RegFile.scala 78:19:@127410.4]
  assign regs_172_io_enable = 1'h1; // @[RegFile.scala 74:20:@127404.4]
  assign regs_173_clock = clock; // @[:@127413.4]
  assign regs_173_reset = io_reset; // @[:@127414.4 RegFile.scala 76:16:@127421.4]
  assign regs_173_io_in = 64'h0; // @[RegFile.scala 75:16:@127420.4]
  assign regs_173_io_reset = reset; // @[RegFile.scala 78:19:@127424.4]
  assign regs_173_io_enable = 1'h1; // @[RegFile.scala 74:20:@127418.4]
  assign regs_174_clock = clock; // @[:@127427.4]
  assign regs_174_reset = io_reset; // @[:@127428.4 RegFile.scala 76:16:@127435.4]
  assign regs_174_io_in = 64'h0; // @[RegFile.scala 75:16:@127434.4]
  assign regs_174_io_reset = reset; // @[RegFile.scala 78:19:@127438.4]
  assign regs_174_io_enable = 1'h1; // @[RegFile.scala 74:20:@127432.4]
  assign regs_175_clock = clock; // @[:@127441.4]
  assign regs_175_reset = io_reset; // @[:@127442.4 RegFile.scala 76:16:@127449.4]
  assign regs_175_io_in = 64'h0; // @[RegFile.scala 75:16:@127448.4]
  assign regs_175_io_reset = reset; // @[RegFile.scala 78:19:@127452.4]
  assign regs_175_io_enable = 1'h1; // @[RegFile.scala 74:20:@127446.4]
  assign regs_176_clock = clock; // @[:@127455.4]
  assign regs_176_reset = io_reset; // @[:@127456.4 RegFile.scala 76:16:@127463.4]
  assign regs_176_io_in = 64'h0; // @[RegFile.scala 75:16:@127462.4]
  assign regs_176_io_reset = reset; // @[RegFile.scala 78:19:@127466.4]
  assign regs_176_io_enable = 1'h1; // @[RegFile.scala 74:20:@127460.4]
  assign regs_177_clock = clock; // @[:@127469.4]
  assign regs_177_reset = io_reset; // @[:@127470.4 RegFile.scala 76:16:@127477.4]
  assign regs_177_io_in = 64'h0; // @[RegFile.scala 75:16:@127476.4]
  assign regs_177_io_reset = reset; // @[RegFile.scala 78:19:@127480.4]
  assign regs_177_io_enable = 1'h1; // @[RegFile.scala 74:20:@127474.4]
  assign regs_178_clock = clock; // @[:@127483.4]
  assign regs_178_reset = io_reset; // @[:@127484.4 RegFile.scala 76:16:@127491.4]
  assign regs_178_io_in = 64'h0; // @[RegFile.scala 75:16:@127490.4]
  assign regs_178_io_reset = reset; // @[RegFile.scala 78:19:@127494.4]
  assign regs_178_io_enable = 1'h1; // @[RegFile.scala 74:20:@127488.4]
  assign regs_179_clock = clock; // @[:@127497.4]
  assign regs_179_reset = io_reset; // @[:@127498.4 RegFile.scala 76:16:@127505.4]
  assign regs_179_io_in = 64'h0; // @[RegFile.scala 75:16:@127504.4]
  assign regs_179_io_reset = reset; // @[RegFile.scala 78:19:@127508.4]
  assign regs_179_io_enable = 1'h1; // @[RegFile.scala 74:20:@127502.4]
  assign regs_180_clock = clock; // @[:@127511.4]
  assign regs_180_reset = io_reset; // @[:@127512.4 RegFile.scala 76:16:@127519.4]
  assign regs_180_io_in = 64'h0; // @[RegFile.scala 75:16:@127518.4]
  assign regs_180_io_reset = reset; // @[RegFile.scala 78:19:@127522.4]
  assign regs_180_io_enable = 1'h1; // @[RegFile.scala 74:20:@127516.4]
  assign regs_181_clock = clock; // @[:@127525.4]
  assign regs_181_reset = io_reset; // @[:@127526.4 RegFile.scala 76:16:@127533.4]
  assign regs_181_io_in = 64'h0; // @[RegFile.scala 75:16:@127532.4]
  assign regs_181_io_reset = reset; // @[RegFile.scala 78:19:@127536.4]
  assign regs_181_io_enable = 1'h1; // @[RegFile.scala 74:20:@127530.4]
  assign regs_182_clock = clock; // @[:@127539.4]
  assign regs_182_reset = io_reset; // @[:@127540.4 RegFile.scala 76:16:@127547.4]
  assign regs_182_io_in = 64'h0; // @[RegFile.scala 75:16:@127546.4]
  assign regs_182_io_reset = reset; // @[RegFile.scala 78:19:@127550.4]
  assign regs_182_io_enable = 1'h1; // @[RegFile.scala 74:20:@127544.4]
  assign regs_183_clock = clock; // @[:@127553.4]
  assign regs_183_reset = io_reset; // @[:@127554.4 RegFile.scala 76:16:@127561.4]
  assign regs_183_io_in = 64'h0; // @[RegFile.scala 75:16:@127560.4]
  assign regs_183_io_reset = reset; // @[RegFile.scala 78:19:@127564.4]
  assign regs_183_io_enable = 1'h1; // @[RegFile.scala 74:20:@127558.4]
  assign regs_184_clock = clock; // @[:@127567.4]
  assign regs_184_reset = io_reset; // @[:@127568.4 RegFile.scala 76:16:@127575.4]
  assign regs_184_io_in = 64'h0; // @[RegFile.scala 75:16:@127574.4]
  assign regs_184_io_reset = reset; // @[RegFile.scala 78:19:@127578.4]
  assign regs_184_io_enable = 1'h1; // @[RegFile.scala 74:20:@127572.4]
  assign regs_185_clock = clock; // @[:@127581.4]
  assign regs_185_reset = io_reset; // @[:@127582.4 RegFile.scala 76:16:@127589.4]
  assign regs_185_io_in = 64'h0; // @[RegFile.scala 75:16:@127588.4]
  assign regs_185_io_reset = reset; // @[RegFile.scala 78:19:@127592.4]
  assign regs_185_io_enable = 1'h1; // @[RegFile.scala 74:20:@127586.4]
  assign regs_186_clock = clock; // @[:@127595.4]
  assign regs_186_reset = io_reset; // @[:@127596.4 RegFile.scala 76:16:@127603.4]
  assign regs_186_io_in = 64'h0; // @[RegFile.scala 75:16:@127602.4]
  assign regs_186_io_reset = reset; // @[RegFile.scala 78:19:@127606.4]
  assign regs_186_io_enable = 1'h1; // @[RegFile.scala 74:20:@127600.4]
  assign regs_187_clock = clock; // @[:@127609.4]
  assign regs_187_reset = io_reset; // @[:@127610.4 RegFile.scala 76:16:@127617.4]
  assign regs_187_io_in = 64'h0; // @[RegFile.scala 75:16:@127616.4]
  assign regs_187_io_reset = reset; // @[RegFile.scala 78:19:@127620.4]
  assign regs_187_io_enable = 1'h1; // @[RegFile.scala 74:20:@127614.4]
  assign regs_188_clock = clock; // @[:@127623.4]
  assign regs_188_reset = io_reset; // @[:@127624.4 RegFile.scala 76:16:@127631.4]
  assign regs_188_io_in = 64'h0; // @[RegFile.scala 75:16:@127630.4]
  assign regs_188_io_reset = reset; // @[RegFile.scala 78:19:@127634.4]
  assign regs_188_io_enable = 1'h1; // @[RegFile.scala 74:20:@127628.4]
  assign regs_189_clock = clock; // @[:@127637.4]
  assign regs_189_reset = io_reset; // @[:@127638.4 RegFile.scala 76:16:@127645.4]
  assign regs_189_io_in = 64'h0; // @[RegFile.scala 75:16:@127644.4]
  assign regs_189_io_reset = reset; // @[RegFile.scala 78:19:@127648.4]
  assign regs_189_io_enable = 1'h1; // @[RegFile.scala 74:20:@127642.4]
  assign regs_190_clock = clock; // @[:@127651.4]
  assign regs_190_reset = io_reset; // @[:@127652.4 RegFile.scala 76:16:@127659.4]
  assign regs_190_io_in = 64'h0; // @[RegFile.scala 75:16:@127658.4]
  assign regs_190_io_reset = reset; // @[RegFile.scala 78:19:@127662.4]
  assign regs_190_io_enable = 1'h1; // @[RegFile.scala 74:20:@127656.4]
  assign regs_191_clock = clock; // @[:@127665.4]
  assign regs_191_reset = io_reset; // @[:@127666.4 RegFile.scala 76:16:@127673.4]
  assign regs_191_io_in = 64'h0; // @[RegFile.scala 75:16:@127672.4]
  assign regs_191_io_reset = reset; // @[RegFile.scala 78:19:@127676.4]
  assign regs_191_io_enable = 1'h1; // @[RegFile.scala 74:20:@127670.4]
  assign regs_192_clock = clock; // @[:@127679.4]
  assign regs_192_reset = io_reset; // @[:@127680.4 RegFile.scala 76:16:@127687.4]
  assign regs_192_io_in = 64'h0; // @[RegFile.scala 75:16:@127686.4]
  assign regs_192_io_reset = reset; // @[RegFile.scala 78:19:@127690.4]
  assign regs_192_io_enable = 1'h1; // @[RegFile.scala 74:20:@127684.4]
  assign regs_193_clock = clock; // @[:@127693.4]
  assign regs_193_reset = io_reset; // @[:@127694.4 RegFile.scala 76:16:@127701.4]
  assign regs_193_io_in = 64'h0; // @[RegFile.scala 75:16:@127700.4]
  assign regs_193_io_reset = reset; // @[RegFile.scala 78:19:@127704.4]
  assign regs_193_io_enable = 1'h1; // @[RegFile.scala 74:20:@127698.4]
  assign regs_194_clock = clock; // @[:@127707.4]
  assign regs_194_reset = io_reset; // @[:@127708.4 RegFile.scala 76:16:@127715.4]
  assign regs_194_io_in = 64'h0; // @[RegFile.scala 75:16:@127714.4]
  assign regs_194_io_reset = reset; // @[RegFile.scala 78:19:@127718.4]
  assign regs_194_io_enable = 1'h1; // @[RegFile.scala 74:20:@127712.4]
  assign regs_195_clock = clock; // @[:@127721.4]
  assign regs_195_reset = io_reset; // @[:@127722.4 RegFile.scala 76:16:@127729.4]
  assign regs_195_io_in = 64'h0; // @[RegFile.scala 75:16:@127728.4]
  assign regs_195_io_reset = reset; // @[RegFile.scala 78:19:@127732.4]
  assign regs_195_io_enable = 1'h1; // @[RegFile.scala 74:20:@127726.4]
  assign regs_196_clock = clock; // @[:@127735.4]
  assign regs_196_reset = io_reset; // @[:@127736.4 RegFile.scala 76:16:@127743.4]
  assign regs_196_io_in = 64'h0; // @[RegFile.scala 75:16:@127742.4]
  assign regs_196_io_reset = reset; // @[RegFile.scala 78:19:@127746.4]
  assign regs_196_io_enable = 1'h1; // @[RegFile.scala 74:20:@127740.4]
  assign regs_197_clock = clock; // @[:@127749.4]
  assign regs_197_reset = io_reset; // @[:@127750.4 RegFile.scala 76:16:@127757.4]
  assign regs_197_io_in = 64'h0; // @[RegFile.scala 75:16:@127756.4]
  assign regs_197_io_reset = reset; // @[RegFile.scala 78:19:@127760.4]
  assign regs_197_io_enable = 1'h1; // @[RegFile.scala 74:20:@127754.4]
  assign regs_198_clock = clock; // @[:@127763.4]
  assign regs_198_reset = io_reset; // @[:@127764.4 RegFile.scala 76:16:@127771.4]
  assign regs_198_io_in = 64'h0; // @[RegFile.scala 75:16:@127770.4]
  assign regs_198_io_reset = reset; // @[RegFile.scala 78:19:@127774.4]
  assign regs_198_io_enable = 1'h1; // @[RegFile.scala 74:20:@127768.4]
  assign regs_199_clock = clock; // @[:@127777.4]
  assign regs_199_reset = io_reset; // @[:@127778.4 RegFile.scala 76:16:@127785.4]
  assign regs_199_io_in = 64'h0; // @[RegFile.scala 75:16:@127784.4]
  assign regs_199_io_reset = reset; // @[RegFile.scala 78:19:@127788.4]
  assign regs_199_io_enable = 1'h1; // @[RegFile.scala 74:20:@127782.4]
  assign regs_200_clock = clock; // @[:@127791.4]
  assign regs_200_reset = io_reset; // @[:@127792.4 RegFile.scala 76:16:@127799.4]
  assign regs_200_io_in = 64'h0; // @[RegFile.scala 75:16:@127798.4]
  assign regs_200_io_reset = reset; // @[RegFile.scala 78:19:@127802.4]
  assign regs_200_io_enable = 1'h1; // @[RegFile.scala 74:20:@127796.4]
  assign regs_201_clock = clock; // @[:@127805.4]
  assign regs_201_reset = io_reset; // @[:@127806.4 RegFile.scala 76:16:@127813.4]
  assign regs_201_io_in = 64'h0; // @[RegFile.scala 75:16:@127812.4]
  assign regs_201_io_reset = reset; // @[RegFile.scala 78:19:@127816.4]
  assign regs_201_io_enable = 1'h1; // @[RegFile.scala 74:20:@127810.4]
  assign regs_202_clock = clock; // @[:@127819.4]
  assign regs_202_reset = io_reset; // @[:@127820.4 RegFile.scala 76:16:@127827.4]
  assign regs_202_io_in = 64'h0; // @[RegFile.scala 75:16:@127826.4]
  assign regs_202_io_reset = reset; // @[RegFile.scala 78:19:@127830.4]
  assign regs_202_io_enable = 1'h1; // @[RegFile.scala 74:20:@127824.4]
  assign regs_203_clock = clock; // @[:@127833.4]
  assign regs_203_reset = io_reset; // @[:@127834.4 RegFile.scala 76:16:@127841.4]
  assign regs_203_io_in = 64'h0; // @[RegFile.scala 75:16:@127840.4]
  assign regs_203_io_reset = reset; // @[RegFile.scala 78:19:@127844.4]
  assign regs_203_io_enable = 1'h1; // @[RegFile.scala 74:20:@127838.4]
  assign regs_204_clock = clock; // @[:@127847.4]
  assign regs_204_reset = io_reset; // @[:@127848.4 RegFile.scala 76:16:@127855.4]
  assign regs_204_io_in = 64'h0; // @[RegFile.scala 75:16:@127854.4]
  assign regs_204_io_reset = reset; // @[RegFile.scala 78:19:@127858.4]
  assign regs_204_io_enable = 1'h1; // @[RegFile.scala 74:20:@127852.4]
  assign regs_205_clock = clock; // @[:@127861.4]
  assign regs_205_reset = io_reset; // @[:@127862.4 RegFile.scala 76:16:@127869.4]
  assign regs_205_io_in = 64'h0; // @[RegFile.scala 75:16:@127868.4]
  assign regs_205_io_reset = reset; // @[RegFile.scala 78:19:@127872.4]
  assign regs_205_io_enable = 1'h1; // @[RegFile.scala 74:20:@127866.4]
  assign regs_206_clock = clock; // @[:@127875.4]
  assign regs_206_reset = io_reset; // @[:@127876.4 RegFile.scala 76:16:@127883.4]
  assign regs_206_io_in = 64'h0; // @[RegFile.scala 75:16:@127882.4]
  assign regs_206_io_reset = reset; // @[RegFile.scala 78:19:@127886.4]
  assign regs_206_io_enable = 1'h1; // @[RegFile.scala 74:20:@127880.4]
  assign regs_207_clock = clock; // @[:@127889.4]
  assign regs_207_reset = io_reset; // @[:@127890.4 RegFile.scala 76:16:@127897.4]
  assign regs_207_io_in = 64'h0; // @[RegFile.scala 75:16:@127896.4]
  assign regs_207_io_reset = reset; // @[RegFile.scala 78:19:@127900.4]
  assign regs_207_io_enable = 1'h1; // @[RegFile.scala 74:20:@127894.4]
  assign regs_208_clock = clock; // @[:@127903.4]
  assign regs_208_reset = io_reset; // @[:@127904.4 RegFile.scala 76:16:@127911.4]
  assign regs_208_io_in = 64'h0; // @[RegFile.scala 75:16:@127910.4]
  assign regs_208_io_reset = reset; // @[RegFile.scala 78:19:@127914.4]
  assign regs_208_io_enable = 1'h1; // @[RegFile.scala 74:20:@127908.4]
  assign regs_209_clock = clock; // @[:@127917.4]
  assign regs_209_reset = io_reset; // @[:@127918.4 RegFile.scala 76:16:@127925.4]
  assign regs_209_io_in = 64'h0; // @[RegFile.scala 75:16:@127924.4]
  assign regs_209_io_reset = reset; // @[RegFile.scala 78:19:@127928.4]
  assign regs_209_io_enable = 1'h1; // @[RegFile.scala 74:20:@127922.4]
  assign regs_210_clock = clock; // @[:@127931.4]
  assign regs_210_reset = io_reset; // @[:@127932.4 RegFile.scala 76:16:@127939.4]
  assign regs_210_io_in = 64'h0; // @[RegFile.scala 75:16:@127938.4]
  assign regs_210_io_reset = reset; // @[RegFile.scala 78:19:@127942.4]
  assign regs_210_io_enable = 1'h1; // @[RegFile.scala 74:20:@127936.4]
  assign regs_211_clock = clock; // @[:@127945.4]
  assign regs_211_reset = io_reset; // @[:@127946.4 RegFile.scala 76:16:@127953.4]
  assign regs_211_io_in = 64'h0; // @[RegFile.scala 75:16:@127952.4]
  assign regs_211_io_reset = reset; // @[RegFile.scala 78:19:@127956.4]
  assign regs_211_io_enable = 1'h1; // @[RegFile.scala 74:20:@127950.4]
  assign regs_212_clock = clock; // @[:@127959.4]
  assign regs_212_reset = io_reset; // @[:@127960.4 RegFile.scala 76:16:@127967.4]
  assign regs_212_io_in = 64'h0; // @[RegFile.scala 75:16:@127966.4]
  assign regs_212_io_reset = reset; // @[RegFile.scala 78:19:@127970.4]
  assign regs_212_io_enable = 1'h1; // @[RegFile.scala 74:20:@127964.4]
  assign regs_213_clock = clock; // @[:@127973.4]
  assign regs_213_reset = io_reset; // @[:@127974.4 RegFile.scala 76:16:@127981.4]
  assign regs_213_io_in = 64'h0; // @[RegFile.scala 75:16:@127980.4]
  assign regs_213_io_reset = reset; // @[RegFile.scala 78:19:@127984.4]
  assign regs_213_io_enable = 1'h1; // @[RegFile.scala 74:20:@127978.4]
  assign regs_214_clock = clock; // @[:@127987.4]
  assign regs_214_reset = io_reset; // @[:@127988.4 RegFile.scala 76:16:@127995.4]
  assign regs_214_io_in = 64'h0; // @[RegFile.scala 75:16:@127994.4]
  assign regs_214_io_reset = reset; // @[RegFile.scala 78:19:@127998.4]
  assign regs_214_io_enable = 1'h1; // @[RegFile.scala 74:20:@127992.4]
  assign regs_215_clock = clock; // @[:@128001.4]
  assign regs_215_reset = io_reset; // @[:@128002.4 RegFile.scala 76:16:@128009.4]
  assign regs_215_io_in = 64'h0; // @[RegFile.scala 75:16:@128008.4]
  assign regs_215_io_reset = reset; // @[RegFile.scala 78:19:@128012.4]
  assign regs_215_io_enable = 1'h1; // @[RegFile.scala 74:20:@128006.4]
  assign regs_216_clock = clock; // @[:@128015.4]
  assign regs_216_reset = io_reset; // @[:@128016.4 RegFile.scala 76:16:@128023.4]
  assign regs_216_io_in = 64'h0; // @[RegFile.scala 75:16:@128022.4]
  assign regs_216_io_reset = reset; // @[RegFile.scala 78:19:@128026.4]
  assign regs_216_io_enable = 1'h1; // @[RegFile.scala 74:20:@128020.4]
  assign regs_217_clock = clock; // @[:@128029.4]
  assign regs_217_reset = io_reset; // @[:@128030.4 RegFile.scala 76:16:@128037.4]
  assign regs_217_io_in = 64'h0; // @[RegFile.scala 75:16:@128036.4]
  assign regs_217_io_reset = reset; // @[RegFile.scala 78:19:@128040.4]
  assign regs_217_io_enable = 1'h1; // @[RegFile.scala 74:20:@128034.4]
  assign regs_218_clock = clock; // @[:@128043.4]
  assign regs_218_reset = io_reset; // @[:@128044.4 RegFile.scala 76:16:@128051.4]
  assign regs_218_io_in = 64'h0; // @[RegFile.scala 75:16:@128050.4]
  assign regs_218_io_reset = reset; // @[RegFile.scala 78:19:@128054.4]
  assign regs_218_io_enable = 1'h1; // @[RegFile.scala 74:20:@128048.4]
  assign regs_219_clock = clock; // @[:@128057.4]
  assign regs_219_reset = io_reset; // @[:@128058.4 RegFile.scala 76:16:@128065.4]
  assign regs_219_io_in = 64'h0; // @[RegFile.scala 75:16:@128064.4]
  assign regs_219_io_reset = reset; // @[RegFile.scala 78:19:@128068.4]
  assign regs_219_io_enable = 1'h1; // @[RegFile.scala 74:20:@128062.4]
  assign regs_220_clock = clock; // @[:@128071.4]
  assign regs_220_reset = io_reset; // @[:@128072.4 RegFile.scala 76:16:@128079.4]
  assign regs_220_io_in = 64'h0; // @[RegFile.scala 75:16:@128078.4]
  assign regs_220_io_reset = reset; // @[RegFile.scala 78:19:@128082.4]
  assign regs_220_io_enable = 1'h1; // @[RegFile.scala 74:20:@128076.4]
  assign regs_221_clock = clock; // @[:@128085.4]
  assign regs_221_reset = io_reset; // @[:@128086.4 RegFile.scala 76:16:@128093.4]
  assign regs_221_io_in = 64'h0; // @[RegFile.scala 75:16:@128092.4]
  assign regs_221_io_reset = reset; // @[RegFile.scala 78:19:@128096.4]
  assign regs_221_io_enable = 1'h1; // @[RegFile.scala 74:20:@128090.4]
  assign regs_222_clock = clock; // @[:@128099.4]
  assign regs_222_reset = io_reset; // @[:@128100.4 RegFile.scala 76:16:@128107.4]
  assign regs_222_io_in = 64'h0; // @[RegFile.scala 75:16:@128106.4]
  assign regs_222_io_reset = reset; // @[RegFile.scala 78:19:@128110.4]
  assign regs_222_io_enable = 1'h1; // @[RegFile.scala 74:20:@128104.4]
  assign regs_223_clock = clock; // @[:@128113.4]
  assign regs_223_reset = io_reset; // @[:@128114.4 RegFile.scala 76:16:@128121.4]
  assign regs_223_io_in = 64'h0; // @[RegFile.scala 75:16:@128120.4]
  assign regs_223_io_reset = reset; // @[RegFile.scala 78:19:@128124.4]
  assign regs_223_io_enable = 1'h1; // @[RegFile.scala 74:20:@128118.4]
  assign regs_224_clock = clock; // @[:@128127.4]
  assign regs_224_reset = io_reset; // @[:@128128.4 RegFile.scala 76:16:@128135.4]
  assign regs_224_io_in = 64'h0; // @[RegFile.scala 75:16:@128134.4]
  assign regs_224_io_reset = reset; // @[RegFile.scala 78:19:@128138.4]
  assign regs_224_io_enable = 1'h1; // @[RegFile.scala 74:20:@128132.4]
  assign regs_225_clock = clock; // @[:@128141.4]
  assign regs_225_reset = io_reset; // @[:@128142.4 RegFile.scala 76:16:@128149.4]
  assign regs_225_io_in = 64'h0; // @[RegFile.scala 75:16:@128148.4]
  assign regs_225_io_reset = reset; // @[RegFile.scala 78:19:@128152.4]
  assign regs_225_io_enable = 1'h1; // @[RegFile.scala 74:20:@128146.4]
  assign regs_226_clock = clock; // @[:@128155.4]
  assign regs_226_reset = io_reset; // @[:@128156.4 RegFile.scala 76:16:@128163.4]
  assign regs_226_io_in = 64'h0; // @[RegFile.scala 75:16:@128162.4]
  assign regs_226_io_reset = reset; // @[RegFile.scala 78:19:@128166.4]
  assign regs_226_io_enable = 1'h1; // @[RegFile.scala 74:20:@128160.4]
  assign regs_227_clock = clock; // @[:@128169.4]
  assign regs_227_reset = io_reset; // @[:@128170.4 RegFile.scala 76:16:@128177.4]
  assign regs_227_io_in = 64'h0; // @[RegFile.scala 75:16:@128176.4]
  assign regs_227_io_reset = reset; // @[RegFile.scala 78:19:@128180.4]
  assign regs_227_io_enable = 1'h1; // @[RegFile.scala 74:20:@128174.4]
  assign regs_228_clock = clock; // @[:@128183.4]
  assign regs_228_reset = io_reset; // @[:@128184.4 RegFile.scala 76:16:@128191.4]
  assign regs_228_io_in = 64'h0; // @[RegFile.scala 75:16:@128190.4]
  assign regs_228_io_reset = reset; // @[RegFile.scala 78:19:@128194.4]
  assign regs_228_io_enable = 1'h1; // @[RegFile.scala 74:20:@128188.4]
  assign regs_229_clock = clock; // @[:@128197.4]
  assign regs_229_reset = io_reset; // @[:@128198.4 RegFile.scala 76:16:@128205.4]
  assign regs_229_io_in = 64'h0; // @[RegFile.scala 75:16:@128204.4]
  assign regs_229_io_reset = reset; // @[RegFile.scala 78:19:@128208.4]
  assign regs_229_io_enable = 1'h1; // @[RegFile.scala 74:20:@128202.4]
  assign regs_230_clock = clock; // @[:@128211.4]
  assign regs_230_reset = io_reset; // @[:@128212.4 RegFile.scala 76:16:@128219.4]
  assign regs_230_io_in = 64'h0; // @[RegFile.scala 75:16:@128218.4]
  assign regs_230_io_reset = reset; // @[RegFile.scala 78:19:@128222.4]
  assign regs_230_io_enable = 1'h1; // @[RegFile.scala 74:20:@128216.4]
  assign regs_231_clock = clock; // @[:@128225.4]
  assign regs_231_reset = io_reset; // @[:@128226.4 RegFile.scala 76:16:@128233.4]
  assign regs_231_io_in = 64'h0; // @[RegFile.scala 75:16:@128232.4]
  assign regs_231_io_reset = reset; // @[RegFile.scala 78:19:@128236.4]
  assign regs_231_io_enable = 1'h1; // @[RegFile.scala 74:20:@128230.4]
  assign regs_232_clock = clock; // @[:@128239.4]
  assign regs_232_reset = io_reset; // @[:@128240.4 RegFile.scala 76:16:@128247.4]
  assign regs_232_io_in = 64'h0; // @[RegFile.scala 75:16:@128246.4]
  assign regs_232_io_reset = reset; // @[RegFile.scala 78:19:@128250.4]
  assign regs_232_io_enable = 1'h1; // @[RegFile.scala 74:20:@128244.4]
  assign regs_233_clock = clock; // @[:@128253.4]
  assign regs_233_reset = io_reset; // @[:@128254.4 RegFile.scala 76:16:@128261.4]
  assign regs_233_io_in = 64'h0; // @[RegFile.scala 75:16:@128260.4]
  assign regs_233_io_reset = reset; // @[RegFile.scala 78:19:@128264.4]
  assign regs_233_io_enable = 1'h1; // @[RegFile.scala 74:20:@128258.4]
  assign regs_234_clock = clock; // @[:@128267.4]
  assign regs_234_reset = io_reset; // @[:@128268.4 RegFile.scala 76:16:@128275.4]
  assign regs_234_io_in = 64'h0; // @[RegFile.scala 75:16:@128274.4]
  assign regs_234_io_reset = reset; // @[RegFile.scala 78:19:@128278.4]
  assign regs_234_io_enable = 1'h1; // @[RegFile.scala 74:20:@128272.4]
  assign regs_235_clock = clock; // @[:@128281.4]
  assign regs_235_reset = io_reset; // @[:@128282.4 RegFile.scala 76:16:@128289.4]
  assign regs_235_io_in = 64'h0; // @[RegFile.scala 75:16:@128288.4]
  assign regs_235_io_reset = reset; // @[RegFile.scala 78:19:@128292.4]
  assign regs_235_io_enable = 1'h1; // @[RegFile.scala 74:20:@128286.4]
  assign regs_236_clock = clock; // @[:@128295.4]
  assign regs_236_reset = io_reset; // @[:@128296.4 RegFile.scala 76:16:@128303.4]
  assign regs_236_io_in = 64'h0; // @[RegFile.scala 75:16:@128302.4]
  assign regs_236_io_reset = reset; // @[RegFile.scala 78:19:@128306.4]
  assign regs_236_io_enable = 1'h1; // @[RegFile.scala 74:20:@128300.4]
  assign regs_237_clock = clock; // @[:@128309.4]
  assign regs_237_reset = io_reset; // @[:@128310.4 RegFile.scala 76:16:@128317.4]
  assign regs_237_io_in = 64'h0; // @[RegFile.scala 75:16:@128316.4]
  assign regs_237_io_reset = reset; // @[RegFile.scala 78:19:@128320.4]
  assign regs_237_io_enable = 1'h1; // @[RegFile.scala 74:20:@128314.4]
  assign regs_238_clock = clock; // @[:@128323.4]
  assign regs_238_reset = io_reset; // @[:@128324.4 RegFile.scala 76:16:@128331.4]
  assign regs_238_io_in = 64'h0; // @[RegFile.scala 75:16:@128330.4]
  assign regs_238_io_reset = reset; // @[RegFile.scala 78:19:@128334.4]
  assign regs_238_io_enable = 1'h1; // @[RegFile.scala 74:20:@128328.4]
  assign regs_239_clock = clock; // @[:@128337.4]
  assign regs_239_reset = io_reset; // @[:@128338.4 RegFile.scala 76:16:@128345.4]
  assign regs_239_io_in = 64'h0; // @[RegFile.scala 75:16:@128344.4]
  assign regs_239_io_reset = reset; // @[RegFile.scala 78:19:@128348.4]
  assign regs_239_io_enable = 1'h1; // @[RegFile.scala 74:20:@128342.4]
  assign regs_240_clock = clock; // @[:@128351.4]
  assign regs_240_reset = io_reset; // @[:@128352.4 RegFile.scala 76:16:@128359.4]
  assign regs_240_io_in = 64'h0; // @[RegFile.scala 75:16:@128358.4]
  assign regs_240_io_reset = reset; // @[RegFile.scala 78:19:@128362.4]
  assign regs_240_io_enable = 1'h1; // @[RegFile.scala 74:20:@128356.4]
  assign regs_241_clock = clock; // @[:@128365.4]
  assign regs_241_reset = io_reset; // @[:@128366.4 RegFile.scala 76:16:@128373.4]
  assign regs_241_io_in = 64'h0; // @[RegFile.scala 75:16:@128372.4]
  assign regs_241_io_reset = reset; // @[RegFile.scala 78:19:@128376.4]
  assign regs_241_io_enable = 1'h1; // @[RegFile.scala 74:20:@128370.4]
  assign regs_242_clock = clock; // @[:@128379.4]
  assign regs_242_reset = io_reset; // @[:@128380.4 RegFile.scala 76:16:@128387.4]
  assign regs_242_io_in = 64'h0; // @[RegFile.scala 75:16:@128386.4]
  assign regs_242_io_reset = reset; // @[RegFile.scala 78:19:@128390.4]
  assign regs_242_io_enable = 1'h1; // @[RegFile.scala 74:20:@128384.4]
  assign regs_243_clock = clock; // @[:@128393.4]
  assign regs_243_reset = io_reset; // @[:@128394.4 RegFile.scala 76:16:@128401.4]
  assign regs_243_io_in = 64'h0; // @[RegFile.scala 75:16:@128400.4]
  assign regs_243_io_reset = reset; // @[RegFile.scala 78:19:@128404.4]
  assign regs_243_io_enable = 1'h1; // @[RegFile.scala 74:20:@128398.4]
  assign regs_244_clock = clock; // @[:@128407.4]
  assign regs_244_reset = io_reset; // @[:@128408.4 RegFile.scala 76:16:@128415.4]
  assign regs_244_io_in = 64'h0; // @[RegFile.scala 75:16:@128414.4]
  assign regs_244_io_reset = reset; // @[RegFile.scala 78:19:@128418.4]
  assign regs_244_io_enable = 1'h1; // @[RegFile.scala 74:20:@128412.4]
  assign regs_245_clock = clock; // @[:@128421.4]
  assign regs_245_reset = io_reset; // @[:@128422.4 RegFile.scala 76:16:@128429.4]
  assign regs_245_io_in = 64'h0; // @[RegFile.scala 75:16:@128428.4]
  assign regs_245_io_reset = reset; // @[RegFile.scala 78:19:@128432.4]
  assign regs_245_io_enable = 1'h1; // @[RegFile.scala 74:20:@128426.4]
  assign regs_246_clock = clock; // @[:@128435.4]
  assign regs_246_reset = io_reset; // @[:@128436.4 RegFile.scala 76:16:@128443.4]
  assign regs_246_io_in = 64'h0; // @[RegFile.scala 75:16:@128442.4]
  assign regs_246_io_reset = reset; // @[RegFile.scala 78:19:@128446.4]
  assign regs_246_io_enable = 1'h1; // @[RegFile.scala 74:20:@128440.4]
  assign regs_247_clock = clock; // @[:@128449.4]
  assign regs_247_reset = io_reset; // @[:@128450.4 RegFile.scala 76:16:@128457.4]
  assign regs_247_io_in = 64'h0; // @[RegFile.scala 75:16:@128456.4]
  assign regs_247_io_reset = reset; // @[RegFile.scala 78:19:@128460.4]
  assign regs_247_io_enable = 1'h1; // @[RegFile.scala 74:20:@128454.4]
  assign regs_248_clock = clock; // @[:@128463.4]
  assign regs_248_reset = io_reset; // @[:@128464.4 RegFile.scala 76:16:@128471.4]
  assign regs_248_io_in = 64'h0; // @[RegFile.scala 75:16:@128470.4]
  assign regs_248_io_reset = reset; // @[RegFile.scala 78:19:@128474.4]
  assign regs_248_io_enable = 1'h1; // @[RegFile.scala 74:20:@128468.4]
  assign regs_249_clock = clock; // @[:@128477.4]
  assign regs_249_reset = io_reset; // @[:@128478.4 RegFile.scala 76:16:@128485.4]
  assign regs_249_io_in = 64'h0; // @[RegFile.scala 75:16:@128484.4]
  assign regs_249_io_reset = reset; // @[RegFile.scala 78:19:@128488.4]
  assign regs_249_io_enable = 1'h1; // @[RegFile.scala 74:20:@128482.4]
  assign regs_250_clock = clock; // @[:@128491.4]
  assign regs_250_reset = io_reset; // @[:@128492.4 RegFile.scala 76:16:@128499.4]
  assign regs_250_io_in = 64'h0; // @[RegFile.scala 75:16:@128498.4]
  assign regs_250_io_reset = reset; // @[RegFile.scala 78:19:@128502.4]
  assign regs_250_io_enable = 1'h1; // @[RegFile.scala 74:20:@128496.4]
  assign regs_251_clock = clock; // @[:@128505.4]
  assign regs_251_reset = io_reset; // @[:@128506.4 RegFile.scala 76:16:@128513.4]
  assign regs_251_io_in = 64'h0; // @[RegFile.scala 75:16:@128512.4]
  assign regs_251_io_reset = reset; // @[RegFile.scala 78:19:@128516.4]
  assign regs_251_io_enable = 1'h1; // @[RegFile.scala 74:20:@128510.4]
  assign regs_252_clock = clock; // @[:@128519.4]
  assign regs_252_reset = io_reset; // @[:@128520.4 RegFile.scala 76:16:@128527.4]
  assign regs_252_io_in = 64'h0; // @[RegFile.scala 75:16:@128526.4]
  assign regs_252_io_reset = reset; // @[RegFile.scala 78:19:@128530.4]
  assign regs_252_io_enable = 1'h1; // @[RegFile.scala 74:20:@128524.4]
  assign regs_253_clock = clock; // @[:@128533.4]
  assign regs_253_reset = io_reset; // @[:@128534.4 RegFile.scala 76:16:@128541.4]
  assign regs_253_io_in = 64'h0; // @[RegFile.scala 75:16:@128540.4]
  assign regs_253_io_reset = reset; // @[RegFile.scala 78:19:@128544.4]
  assign regs_253_io_enable = 1'h1; // @[RegFile.scala 74:20:@128538.4]
  assign regs_254_clock = clock; // @[:@128547.4]
  assign regs_254_reset = io_reset; // @[:@128548.4 RegFile.scala 76:16:@128555.4]
  assign regs_254_io_in = 64'h0; // @[RegFile.scala 75:16:@128554.4]
  assign regs_254_io_reset = reset; // @[RegFile.scala 78:19:@128558.4]
  assign regs_254_io_enable = 1'h1; // @[RegFile.scala 74:20:@128552.4]
  assign regs_255_clock = clock; // @[:@128561.4]
  assign regs_255_reset = io_reset; // @[:@128562.4 RegFile.scala 76:16:@128569.4]
  assign regs_255_io_in = 64'h0; // @[RegFile.scala 75:16:@128568.4]
  assign regs_255_io_reset = reset; // @[RegFile.scala 78:19:@128572.4]
  assign regs_255_io_enable = 1'h1; // @[RegFile.scala 74:20:@128566.4]
  assign regs_256_clock = clock; // @[:@128575.4]
  assign regs_256_reset = io_reset; // @[:@128576.4 RegFile.scala 76:16:@128583.4]
  assign regs_256_io_in = 64'h0; // @[RegFile.scala 75:16:@128582.4]
  assign regs_256_io_reset = reset; // @[RegFile.scala 78:19:@128586.4]
  assign regs_256_io_enable = 1'h1; // @[RegFile.scala 74:20:@128580.4]
  assign regs_257_clock = clock; // @[:@128589.4]
  assign regs_257_reset = io_reset; // @[:@128590.4 RegFile.scala 76:16:@128597.4]
  assign regs_257_io_in = 64'h0; // @[RegFile.scala 75:16:@128596.4]
  assign regs_257_io_reset = reset; // @[RegFile.scala 78:19:@128600.4]
  assign regs_257_io_enable = 1'h1; // @[RegFile.scala 74:20:@128594.4]
  assign regs_258_clock = clock; // @[:@128603.4]
  assign regs_258_reset = io_reset; // @[:@128604.4 RegFile.scala 76:16:@128611.4]
  assign regs_258_io_in = 64'h0; // @[RegFile.scala 75:16:@128610.4]
  assign regs_258_io_reset = reset; // @[RegFile.scala 78:19:@128614.4]
  assign regs_258_io_enable = 1'h1; // @[RegFile.scala 74:20:@128608.4]
  assign regs_259_clock = clock; // @[:@128617.4]
  assign regs_259_reset = io_reset; // @[:@128618.4 RegFile.scala 76:16:@128625.4]
  assign regs_259_io_in = 64'h0; // @[RegFile.scala 75:16:@128624.4]
  assign regs_259_io_reset = reset; // @[RegFile.scala 78:19:@128628.4]
  assign regs_259_io_enable = 1'h1; // @[RegFile.scala 74:20:@128622.4]
  assign regs_260_clock = clock; // @[:@128631.4]
  assign regs_260_reset = io_reset; // @[:@128632.4 RegFile.scala 76:16:@128639.4]
  assign regs_260_io_in = 64'h0; // @[RegFile.scala 75:16:@128638.4]
  assign regs_260_io_reset = reset; // @[RegFile.scala 78:19:@128642.4]
  assign regs_260_io_enable = 1'h1; // @[RegFile.scala 74:20:@128636.4]
  assign regs_261_clock = clock; // @[:@128645.4]
  assign regs_261_reset = io_reset; // @[:@128646.4 RegFile.scala 76:16:@128653.4]
  assign regs_261_io_in = 64'h0; // @[RegFile.scala 75:16:@128652.4]
  assign regs_261_io_reset = reset; // @[RegFile.scala 78:19:@128656.4]
  assign regs_261_io_enable = 1'h1; // @[RegFile.scala 74:20:@128650.4]
  assign regs_262_clock = clock; // @[:@128659.4]
  assign regs_262_reset = io_reset; // @[:@128660.4 RegFile.scala 76:16:@128667.4]
  assign regs_262_io_in = 64'h0; // @[RegFile.scala 75:16:@128666.4]
  assign regs_262_io_reset = reset; // @[RegFile.scala 78:19:@128670.4]
  assign regs_262_io_enable = 1'h1; // @[RegFile.scala 74:20:@128664.4]
  assign regs_263_clock = clock; // @[:@128673.4]
  assign regs_263_reset = io_reset; // @[:@128674.4 RegFile.scala 76:16:@128681.4]
  assign regs_263_io_in = 64'h0; // @[RegFile.scala 75:16:@128680.4]
  assign regs_263_io_reset = reset; // @[RegFile.scala 78:19:@128684.4]
  assign regs_263_io_enable = 1'h1; // @[RegFile.scala 74:20:@128678.4]
  assign regs_264_clock = clock; // @[:@128687.4]
  assign regs_264_reset = io_reset; // @[:@128688.4 RegFile.scala 76:16:@128695.4]
  assign regs_264_io_in = 64'h0; // @[RegFile.scala 75:16:@128694.4]
  assign regs_264_io_reset = reset; // @[RegFile.scala 78:19:@128698.4]
  assign regs_264_io_enable = 1'h1; // @[RegFile.scala 74:20:@128692.4]
  assign regs_265_clock = clock; // @[:@128701.4]
  assign regs_265_reset = io_reset; // @[:@128702.4 RegFile.scala 76:16:@128709.4]
  assign regs_265_io_in = 64'h0; // @[RegFile.scala 75:16:@128708.4]
  assign regs_265_io_reset = reset; // @[RegFile.scala 78:19:@128712.4]
  assign regs_265_io_enable = 1'h1; // @[RegFile.scala 74:20:@128706.4]
  assign regs_266_clock = clock; // @[:@128715.4]
  assign regs_266_reset = io_reset; // @[:@128716.4 RegFile.scala 76:16:@128723.4]
  assign regs_266_io_in = 64'h0; // @[RegFile.scala 75:16:@128722.4]
  assign regs_266_io_reset = reset; // @[RegFile.scala 78:19:@128726.4]
  assign regs_266_io_enable = 1'h1; // @[RegFile.scala 74:20:@128720.4]
  assign regs_267_clock = clock; // @[:@128729.4]
  assign regs_267_reset = io_reset; // @[:@128730.4 RegFile.scala 76:16:@128737.4]
  assign regs_267_io_in = 64'h0; // @[RegFile.scala 75:16:@128736.4]
  assign regs_267_io_reset = reset; // @[RegFile.scala 78:19:@128740.4]
  assign regs_267_io_enable = 1'h1; // @[RegFile.scala 74:20:@128734.4]
  assign regs_268_clock = clock; // @[:@128743.4]
  assign regs_268_reset = io_reset; // @[:@128744.4 RegFile.scala 76:16:@128751.4]
  assign regs_268_io_in = 64'h0; // @[RegFile.scala 75:16:@128750.4]
  assign regs_268_io_reset = reset; // @[RegFile.scala 78:19:@128754.4]
  assign regs_268_io_enable = 1'h1; // @[RegFile.scala 74:20:@128748.4]
  assign regs_269_clock = clock; // @[:@128757.4]
  assign regs_269_reset = io_reset; // @[:@128758.4 RegFile.scala 76:16:@128765.4]
  assign regs_269_io_in = 64'h0; // @[RegFile.scala 75:16:@128764.4]
  assign regs_269_io_reset = reset; // @[RegFile.scala 78:19:@128768.4]
  assign regs_269_io_enable = 1'h1; // @[RegFile.scala 74:20:@128762.4]
  assign regs_270_clock = clock; // @[:@128771.4]
  assign regs_270_reset = io_reset; // @[:@128772.4 RegFile.scala 76:16:@128779.4]
  assign regs_270_io_in = 64'h0; // @[RegFile.scala 75:16:@128778.4]
  assign regs_270_io_reset = reset; // @[RegFile.scala 78:19:@128782.4]
  assign regs_270_io_enable = 1'h1; // @[RegFile.scala 74:20:@128776.4]
  assign regs_271_clock = clock; // @[:@128785.4]
  assign regs_271_reset = io_reset; // @[:@128786.4 RegFile.scala 76:16:@128793.4]
  assign regs_271_io_in = 64'h0; // @[RegFile.scala 75:16:@128792.4]
  assign regs_271_io_reset = reset; // @[RegFile.scala 78:19:@128796.4]
  assign regs_271_io_enable = 1'h1; // @[RegFile.scala 74:20:@128790.4]
  assign regs_272_clock = clock; // @[:@128799.4]
  assign regs_272_reset = io_reset; // @[:@128800.4 RegFile.scala 76:16:@128807.4]
  assign regs_272_io_in = 64'h0; // @[RegFile.scala 75:16:@128806.4]
  assign regs_272_io_reset = reset; // @[RegFile.scala 78:19:@128810.4]
  assign regs_272_io_enable = 1'h1; // @[RegFile.scala 74:20:@128804.4]
  assign regs_273_clock = clock; // @[:@128813.4]
  assign regs_273_reset = io_reset; // @[:@128814.4 RegFile.scala 76:16:@128821.4]
  assign regs_273_io_in = 64'h0; // @[RegFile.scala 75:16:@128820.4]
  assign regs_273_io_reset = reset; // @[RegFile.scala 78:19:@128824.4]
  assign regs_273_io_enable = 1'h1; // @[RegFile.scala 74:20:@128818.4]
  assign regs_274_clock = clock; // @[:@128827.4]
  assign regs_274_reset = io_reset; // @[:@128828.4 RegFile.scala 76:16:@128835.4]
  assign regs_274_io_in = 64'h0; // @[RegFile.scala 75:16:@128834.4]
  assign regs_274_io_reset = reset; // @[RegFile.scala 78:19:@128838.4]
  assign regs_274_io_enable = 1'h1; // @[RegFile.scala 74:20:@128832.4]
  assign regs_275_clock = clock; // @[:@128841.4]
  assign regs_275_reset = io_reset; // @[:@128842.4 RegFile.scala 76:16:@128849.4]
  assign regs_275_io_in = 64'h0; // @[RegFile.scala 75:16:@128848.4]
  assign regs_275_io_reset = reset; // @[RegFile.scala 78:19:@128852.4]
  assign regs_275_io_enable = 1'h1; // @[RegFile.scala 74:20:@128846.4]
  assign regs_276_clock = clock; // @[:@128855.4]
  assign regs_276_reset = io_reset; // @[:@128856.4 RegFile.scala 76:16:@128863.4]
  assign regs_276_io_in = 64'h0; // @[RegFile.scala 75:16:@128862.4]
  assign regs_276_io_reset = reset; // @[RegFile.scala 78:19:@128866.4]
  assign regs_276_io_enable = 1'h1; // @[RegFile.scala 74:20:@128860.4]
  assign regs_277_clock = clock; // @[:@128869.4]
  assign regs_277_reset = io_reset; // @[:@128870.4 RegFile.scala 76:16:@128877.4]
  assign regs_277_io_in = 64'h0; // @[RegFile.scala 75:16:@128876.4]
  assign regs_277_io_reset = reset; // @[RegFile.scala 78:19:@128880.4]
  assign regs_277_io_enable = 1'h1; // @[RegFile.scala 74:20:@128874.4]
  assign regs_278_clock = clock; // @[:@128883.4]
  assign regs_278_reset = io_reset; // @[:@128884.4 RegFile.scala 76:16:@128891.4]
  assign regs_278_io_in = 64'h0; // @[RegFile.scala 75:16:@128890.4]
  assign regs_278_io_reset = reset; // @[RegFile.scala 78:19:@128894.4]
  assign regs_278_io_enable = 1'h1; // @[RegFile.scala 74:20:@128888.4]
  assign regs_279_clock = clock; // @[:@128897.4]
  assign regs_279_reset = io_reset; // @[:@128898.4 RegFile.scala 76:16:@128905.4]
  assign regs_279_io_in = 64'h0; // @[RegFile.scala 75:16:@128904.4]
  assign regs_279_io_reset = reset; // @[RegFile.scala 78:19:@128908.4]
  assign regs_279_io_enable = 1'h1; // @[RegFile.scala 74:20:@128902.4]
  assign regs_280_clock = clock; // @[:@128911.4]
  assign regs_280_reset = io_reset; // @[:@128912.4 RegFile.scala 76:16:@128919.4]
  assign regs_280_io_in = 64'h0; // @[RegFile.scala 75:16:@128918.4]
  assign regs_280_io_reset = reset; // @[RegFile.scala 78:19:@128922.4]
  assign regs_280_io_enable = 1'h1; // @[RegFile.scala 74:20:@128916.4]
  assign regs_281_clock = clock; // @[:@128925.4]
  assign regs_281_reset = io_reset; // @[:@128926.4 RegFile.scala 76:16:@128933.4]
  assign regs_281_io_in = 64'h0; // @[RegFile.scala 75:16:@128932.4]
  assign regs_281_io_reset = reset; // @[RegFile.scala 78:19:@128936.4]
  assign regs_281_io_enable = 1'h1; // @[RegFile.scala 74:20:@128930.4]
  assign regs_282_clock = clock; // @[:@128939.4]
  assign regs_282_reset = io_reset; // @[:@128940.4 RegFile.scala 76:16:@128947.4]
  assign regs_282_io_in = 64'h0; // @[RegFile.scala 75:16:@128946.4]
  assign regs_282_io_reset = reset; // @[RegFile.scala 78:19:@128950.4]
  assign regs_282_io_enable = 1'h1; // @[RegFile.scala 74:20:@128944.4]
  assign regs_283_clock = clock; // @[:@128953.4]
  assign regs_283_reset = io_reset; // @[:@128954.4 RegFile.scala 76:16:@128961.4]
  assign regs_283_io_in = 64'h0; // @[RegFile.scala 75:16:@128960.4]
  assign regs_283_io_reset = reset; // @[RegFile.scala 78:19:@128964.4]
  assign regs_283_io_enable = 1'h1; // @[RegFile.scala 74:20:@128958.4]
  assign regs_284_clock = clock; // @[:@128967.4]
  assign regs_284_reset = io_reset; // @[:@128968.4 RegFile.scala 76:16:@128975.4]
  assign regs_284_io_in = 64'h0; // @[RegFile.scala 75:16:@128974.4]
  assign regs_284_io_reset = reset; // @[RegFile.scala 78:19:@128978.4]
  assign regs_284_io_enable = 1'h1; // @[RegFile.scala 74:20:@128972.4]
  assign regs_285_clock = clock; // @[:@128981.4]
  assign regs_285_reset = io_reset; // @[:@128982.4 RegFile.scala 76:16:@128989.4]
  assign regs_285_io_in = 64'h0; // @[RegFile.scala 75:16:@128988.4]
  assign regs_285_io_reset = reset; // @[RegFile.scala 78:19:@128992.4]
  assign regs_285_io_enable = 1'h1; // @[RegFile.scala 74:20:@128986.4]
  assign regs_286_clock = clock; // @[:@128995.4]
  assign regs_286_reset = io_reset; // @[:@128996.4 RegFile.scala 76:16:@129003.4]
  assign regs_286_io_in = 64'h0; // @[RegFile.scala 75:16:@129002.4]
  assign regs_286_io_reset = reset; // @[RegFile.scala 78:19:@129006.4]
  assign regs_286_io_enable = 1'h1; // @[RegFile.scala 74:20:@129000.4]
  assign regs_287_clock = clock; // @[:@129009.4]
  assign regs_287_reset = io_reset; // @[:@129010.4 RegFile.scala 76:16:@129017.4]
  assign regs_287_io_in = 64'h0; // @[RegFile.scala 75:16:@129016.4]
  assign regs_287_io_reset = reset; // @[RegFile.scala 78:19:@129020.4]
  assign regs_287_io_enable = 1'h1; // @[RegFile.scala 74:20:@129014.4]
  assign regs_288_clock = clock; // @[:@129023.4]
  assign regs_288_reset = io_reset; // @[:@129024.4 RegFile.scala 76:16:@129031.4]
  assign regs_288_io_in = 64'h0; // @[RegFile.scala 75:16:@129030.4]
  assign regs_288_io_reset = reset; // @[RegFile.scala 78:19:@129034.4]
  assign regs_288_io_enable = 1'h1; // @[RegFile.scala 74:20:@129028.4]
  assign regs_289_clock = clock; // @[:@129037.4]
  assign regs_289_reset = io_reset; // @[:@129038.4 RegFile.scala 76:16:@129045.4]
  assign regs_289_io_in = 64'h0; // @[RegFile.scala 75:16:@129044.4]
  assign regs_289_io_reset = reset; // @[RegFile.scala 78:19:@129048.4]
  assign regs_289_io_enable = 1'h1; // @[RegFile.scala 74:20:@129042.4]
  assign regs_290_clock = clock; // @[:@129051.4]
  assign regs_290_reset = io_reset; // @[:@129052.4 RegFile.scala 76:16:@129059.4]
  assign regs_290_io_in = 64'h0; // @[RegFile.scala 75:16:@129058.4]
  assign regs_290_io_reset = reset; // @[RegFile.scala 78:19:@129062.4]
  assign regs_290_io_enable = 1'h1; // @[RegFile.scala 74:20:@129056.4]
  assign regs_291_clock = clock; // @[:@129065.4]
  assign regs_291_reset = io_reset; // @[:@129066.4 RegFile.scala 76:16:@129073.4]
  assign regs_291_io_in = 64'h0; // @[RegFile.scala 75:16:@129072.4]
  assign regs_291_io_reset = reset; // @[RegFile.scala 78:19:@129076.4]
  assign regs_291_io_enable = 1'h1; // @[RegFile.scala 74:20:@129070.4]
  assign regs_292_clock = clock; // @[:@129079.4]
  assign regs_292_reset = io_reset; // @[:@129080.4 RegFile.scala 76:16:@129087.4]
  assign regs_292_io_in = 64'h0; // @[RegFile.scala 75:16:@129086.4]
  assign regs_292_io_reset = reset; // @[RegFile.scala 78:19:@129090.4]
  assign regs_292_io_enable = 1'h1; // @[RegFile.scala 74:20:@129084.4]
  assign regs_293_clock = clock; // @[:@129093.4]
  assign regs_293_reset = io_reset; // @[:@129094.4 RegFile.scala 76:16:@129101.4]
  assign regs_293_io_in = 64'h0; // @[RegFile.scala 75:16:@129100.4]
  assign regs_293_io_reset = reset; // @[RegFile.scala 78:19:@129104.4]
  assign regs_293_io_enable = 1'h1; // @[RegFile.scala 74:20:@129098.4]
  assign regs_294_clock = clock; // @[:@129107.4]
  assign regs_294_reset = io_reset; // @[:@129108.4 RegFile.scala 76:16:@129115.4]
  assign regs_294_io_in = 64'h0; // @[RegFile.scala 75:16:@129114.4]
  assign regs_294_io_reset = reset; // @[RegFile.scala 78:19:@129118.4]
  assign regs_294_io_enable = 1'h1; // @[RegFile.scala 74:20:@129112.4]
  assign regs_295_clock = clock; // @[:@129121.4]
  assign regs_295_reset = io_reset; // @[:@129122.4 RegFile.scala 76:16:@129129.4]
  assign regs_295_io_in = 64'h0; // @[RegFile.scala 75:16:@129128.4]
  assign regs_295_io_reset = reset; // @[RegFile.scala 78:19:@129132.4]
  assign regs_295_io_enable = 1'h1; // @[RegFile.scala 74:20:@129126.4]
  assign regs_296_clock = clock; // @[:@129135.4]
  assign regs_296_reset = io_reset; // @[:@129136.4 RegFile.scala 76:16:@129143.4]
  assign regs_296_io_in = 64'h0; // @[RegFile.scala 75:16:@129142.4]
  assign regs_296_io_reset = reset; // @[RegFile.scala 78:19:@129146.4]
  assign regs_296_io_enable = 1'h1; // @[RegFile.scala 74:20:@129140.4]
  assign regs_297_clock = clock; // @[:@129149.4]
  assign regs_297_reset = io_reset; // @[:@129150.4 RegFile.scala 76:16:@129157.4]
  assign regs_297_io_in = 64'h0; // @[RegFile.scala 75:16:@129156.4]
  assign regs_297_io_reset = reset; // @[RegFile.scala 78:19:@129160.4]
  assign regs_297_io_enable = 1'h1; // @[RegFile.scala 74:20:@129154.4]
  assign regs_298_clock = clock; // @[:@129163.4]
  assign regs_298_reset = io_reset; // @[:@129164.4 RegFile.scala 76:16:@129171.4]
  assign regs_298_io_in = 64'h0; // @[RegFile.scala 75:16:@129170.4]
  assign regs_298_io_reset = reset; // @[RegFile.scala 78:19:@129174.4]
  assign regs_298_io_enable = 1'h1; // @[RegFile.scala 74:20:@129168.4]
  assign regs_299_clock = clock; // @[:@129177.4]
  assign regs_299_reset = io_reset; // @[:@129178.4 RegFile.scala 76:16:@129185.4]
  assign regs_299_io_in = 64'h0; // @[RegFile.scala 75:16:@129184.4]
  assign regs_299_io_reset = reset; // @[RegFile.scala 78:19:@129188.4]
  assign regs_299_io_enable = 1'h1; // @[RegFile.scala 74:20:@129182.4]
  assign regs_300_clock = clock; // @[:@129191.4]
  assign regs_300_reset = io_reset; // @[:@129192.4 RegFile.scala 76:16:@129199.4]
  assign regs_300_io_in = 64'h0; // @[RegFile.scala 75:16:@129198.4]
  assign regs_300_io_reset = reset; // @[RegFile.scala 78:19:@129202.4]
  assign regs_300_io_enable = 1'h1; // @[RegFile.scala 74:20:@129196.4]
  assign regs_301_clock = clock; // @[:@129205.4]
  assign regs_301_reset = io_reset; // @[:@129206.4 RegFile.scala 76:16:@129213.4]
  assign regs_301_io_in = 64'h0; // @[RegFile.scala 75:16:@129212.4]
  assign regs_301_io_reset = reset; // @[RegFile.scala 78:19:@129216.4]
  assign regs_301_io_enable = 1'h1; // @[RegFile.scala 74:20:@129210.4]
  assign regs_302_clock = clock; // @[:@129219.4]
  assign regs_302_reset = io_reset; // @[:@129220.4 RegFile.scala 76:16:@129227.4]
  assign regs_302_io_in = 64'h0; // @[RegFile.scala 75:16:@129226.4]
  assign regs_302_io_reset = reset; // @[RegFile.scala 78:19:@129230.4]
  assign regs_302_io_enable = 1'h1; // @[RegFile.scala 74:20:@129224.4]
  assign regs_303_clock = clock; // @[:@129233.4]
  assign regs_303_reset = io_reset; // @[:@129234.4 RegFile.scala 76:16:@129241.4]
  assign regs_303_io_in = 64'h0; // @[RegFile.scala 75:16:@129240.4]
  assign regs_303_io_reset = reset; // @[RegFile.scala 78:19:@129244.4]
  assign regs_303_io_enable = 1'h1; // @[RegFile.scala 74:20:@129238.4]
  assign regs_304_clock = clock; // @[:@129247.4]
  assign regs_304_reset = io_reset; // @[:@129248.4 RegFile.scala 76:16:@129255.4]
  assign regs_304_io_in = 64'h0; // @[RegFile.scala 75:16:@129254.4]
  assign regs_304_io_reset = reset; // @[RegFile.scala 78:19:@129258.4]
  assign regs_304_io_enable = 1'h1; // @[RegFile.scala 74:20:@129252.4]
  assign regs_305_clock = clock; // @[:@129261.4]
  assign regs_305_reset = io_reset; // @[:@129262.4 RegFile.scala 76:16:@129269.4]
  assign regs_305_io_in = 64'h0; // @[RegFile.scala 75:16:@129268.4]
  assign regs_305_io_reset = reset; // @[RegFile.scala 78:19:@129272.4]
  assign regs_305_io_enable = 1'h1; // @[RegFile.scala 74:20:@129266.4]
  assign regs_306_clock = clock; // @[:@129275.4]
  assign regs_306_reset = io_reset; // @[:@129276.4 RegFile.scala 76:16:@129283.4]
  assign regs_306_io_in = 64'h0; // @[RegFile.scala 75:16:@129282.4]
  assign regs_306_io_reset = reset; // @[RegFile.scala 78:19:@129286.4]
  assign regs_306_io_enable = 1'h1; // @[RegFile.scala 74:20:@129280.4]
  assign regs_307_clock = clock; // @[:@129289.4]
  assign regs_307_reset = io_reset; // @[:@129290.4 RegFile.scala 76:16:@129297.4]
  assign regs_307_io_in = 64'h0; // @[RegFile.scala 75:16:@129296.4]
  assign regs_307_io_reset = reset; // @[RegFile.scala 78:19:@129300.4]
  assign regs_307_io_enable = 1'h1; // @[RegFile.scala 74:20:@129294.4]
  assign regs_308_clock = clock; // @[:@129303.4]
  assign regs_308_reset = io_reset; // @[:@129304.4 RegFile.scala 76:16:@129311.4]
  assign regs_308_io_in = 64'h0; // @[RegFile.scala 75:16:@129310.4]
  assign regs_308_io_reset = reset; // @[RegFile.scala 78:19:@129314.4]
  assign regs_308_io_enable = 1'h1; // @[RegFile.scala 74:20:@129308.4]
  assign regs_309_clock = clock; // @[:@129317.4]
  assign regs_309_reset = io_reset; // @[:@129318.4 RegFile.scala 76:16:@129325.4]
  assign regs_309_io_in = 64'h0; // @[RegFile.scala 75:16:@129324.4]
  assign regs_309_io_reset = reset; // @[RegFile.scala 78:19:@129328.4]
  assign regs_309_io_enable = 1'h1; // @[RegFile.scala 74:20:@129322.4]
  assign regs_310_clock = clock; // @[:@129331.4]
  assign regs_310_reset = io_reset; // @[:@129332.4 RegFile.scala 76:16:@129339.4]
  assign regs_310_io_in = 64'h0; // @[RegFile.scala 75:16:@129338.4]
  assign regs_310_io_reset = reset; // @[RegFile.scala 78:19:@129342.4]
  assign regs_310_io_enable = 1'h1; // @[RegFile.scala 74:20:@129336.4]
  assign regs_311_clock = clock; // @[:@129345.4]
  assign regs_311_reset = io_reset; // @[:@129346.4 RegFile.scala 76:16:@129353.4]
  assign regs_311_io_in = 64'h0; // @[RegFile.scala 75:16:@129352.4]
  assign regs_311_io_reset = reset; // @[RegFile.scala 78:19:@129356.4]
  assign regs_311_io_enable = 1'h1; // @[RegFile.scala 74:20:@129350.4]
  assign regs_312_clock = clock; // @[:@129359.4]
  assign regs_312_reset = io_reset; // @[:@129360.4 RegFile.scala 76:16:@129367.4]
  assign regs_312_io_in = 64'h0; // @[RegFile.scala 75:16:@129366.4]
  assign regs_312_io_reset = reset; // @[RegFile.scala 78:19:@129370.4]
  assign regs_312_io_enable = 1'h1; // @[RegFile.scala 74:20:@129364.4]
  assign regs_313_clock = clock; // @[:@129373.4]
  assign regs_313_reset = io_reset; // @[:@129374.4 RegFile.scala 76:16:@129381.4]
  assign regs_313_io_in = 64'h0; // @[RegFile.scala 75:16:@129380.4]
  assign regs_313_io_reset = reset; // @[RegFile.scala 78:19:@129384.4]
  assign regs_313_io_enable = 1'h1; // @[RegFile.scala 74:20:@129378.4]
  assign regs_314_clock = clock; // @[:@129387.4]
  assign regs_314_reset = io_reset; // @[:@129388.4 RegFile.scala 76:16:@129395.4]
  assign regs_314_io_in = 64'h0; // @[RegFile.scala 75:16:@129394.4]
  assign regs_314_io_reset = reset; // @[RegFile.scala 78:19:@129398.4]
  assign regs_314_io_enable = 1'h1; // @[RegFile.scala 74:20:@129392.4]
  assign regs_315_clock = clock; // @[:@129401.4]
  assign regs_315_reset = io_reset; // @[:@129402.4 RegFile.scala 76:16:@129409.4]
  assign regs_315_io_in = 64'h0; // @[RegFile.scala 75:16:@129408.4]
  assign regs_315_io_reset = reset; // @[RegFile.scala 78:19:@129412.4]
  assign regs_315_io_enable = 1'h1; // @[RegFile.scala 74:20:@129406.4]
  assign regs_316_clock = clock; // @[:@129415.4]
  assign regs_316_reset = io_reset; // @[:@129416.4 RegFile.scala 76:16:@129423.4]
  assign regs_316_io_in = 64'h0; // @[RegFile.scala 75:16:@129422.4]
  assign regs_316_io_reset = reset; // @[RegFile.scala 78:19:@129426.4]
  assign regs_316_io_enable = 1'h1; // @[RegFile.scala 74:20:@129420.4]
  assign regs_317_clock = clock; // @[:@129429.4]
  assign regs_317_reset = io_reset; // @[:@129430.4 RegFile.scala 76:16:@129437.4]
  assign regs_317_io_in = 64'h0; // @[RegFile.scala 75:16:@129436.4]
  assign regs_317_io_reset = reset; // @[RegFile.scala 78:19:@129440.4]
  assign regs_317_io_enable = 1'h1; // @[RegFile.scala 74:20:@129434.4]
  assign regs_318_clock = clock; // @[:@129443.4]
  assign regs_318_reset = io_reset; // @[:@129444.4 RegFile.scala 76:16:@129451.4]
  assign regs_318_io_in = 64'h0; // @[RegFile.scala 75:16:@129450.4]
  assign regs_318_io_reset = reset; // @[RegFile.scala 78:19:@129454.4]
  assign regs_318_io_enable = 1'h1; // @[RegFile.scala 74:20:@129448.4]
  assign regs_319_clock = clock; // @[:@129457.4]
  assign regs_319_reset = io_reset; // @[:@129458.4 RegFile.scala 76:16:@129465.4]
  assign regs_319_io_in = 64'h0; // @[RegFile.scala 75:16:@129464.4]
  assign regs_319_io_reset = reset; // @[RegFile.scala 78:19:@129468.4]
  assign regs_319_io_enable = 1'h1; // @[RegFile.scala 74:20:@129462.4]
  assign regs_320_clock = clock; // @[:@129471.4]
  assign regs_320_reset = io_reset; // @[:@129472.4 RegFile.scala 76:16:@129479.4]
  assign regs_320_io_in = 64'h0; // @[RegFile.scala 75:16:@129478.4]
  assign regs_320_io_reset = reset; // @[RegFile.scala 78:19:@129482.4]
  assign regs_320_io_enable = 1'h1; // @[RegFile.scala 74:20:@129476.4]
  assign regs_321_clock = clock; // @[:@129485.4]
  assign regs_321_reset = io_reset; // @[:@129486.4 RegFile.scala 76:16:@129493.4]
  assign regs_321_io_in = 64'h0; // @[RegFile.scala 75:16:@129492.4]
  assign regs_321_io_reset = reset; // @[RegFile.scala 78:19:@129496.4]
  assign regs_321_io_enable = 1'h1; // @[RegFile.scala 74:20:@129490.4]
  assign regs_322_clock = clock; // @[:@129499.4]
  assign regs_322_reset = io_reset; // @[:@129500.4 RegFile.scala 76:16:@129507.4]
  assign regs_322_io_in = 64'h0; // @[RegFile.scala 75:16:@129506.4]
  assign regs_322_io_reset = reset; // @[RegFile.scala 78:19:@129510.4]
  assign regs_322_io_enable = 1'h1; // @[RegFile.scala 74:20:@129504.4]
  assign regs_323_clock = clock; // @[:@129513.4]
  assign regs_323_reset = io_reset; // @[:@129514.4 RegFile.scala 76:16:@129521.4]
  assign regs_323_io_in = 64'h0; // @[RegFile.scala 75:16:@129520.4]
  assign regs_323_io_reset = reset; // @[RegFile.scala 78:19:@129524.4]
  assign regs_323_io_enable = 1'h1; // @[RegFile.scala 74:20:@129518.4]
  assign regs_324_clock = clock; // @[:@129527.4]
  assign regs_324_reset = io_reset; // @[:@129528.4 RegFile.scala 76:16:@129535.4]
  assign regs_324_io_in = 64'h0; // @[RegFile.scala 75:16:@129534.4]
  assign regs_324_io_reset = reset; // @[RegFile.scala 78:19:@129538.4]
  assign regs_324_io_enable = 1'h1; // @[RegFile.scala 74:20:@129532.4]
  assign regs_325_clock = clock; // @[:@129541.4]
  assign regs_325_reset = io_reset; // @[:@129542.4 RegFile.scala 76:16:@129549.4]
  assign regs_325_io_in = 64'h0; // @[RegFile.scala 75:16:@129548.4]
  assign regs_325_io_reset = reset; // @[RegFile.scala 78:19:@129552.4]
  assign regs_325_io_enable = 1'h1; // @[RegFile.scala 74:20:@129546.4]
  assign regs_326_clock = clock; // @[:@129555.4]
  assign regs_326_reset = io_reset; // @[:@129556.4 RegFile.scala 76:16:@129563.4]
  assign regs_326_io_in = 64'h0; // @[RegFile.scala 75:16:@129562.4]
  assign regs_326_io_reset = reset; // @[RegFile.scala 78:19:@129566.4]
  assign regs_326_io_enable = 1'h1; // @[RegFile.scala 74:20:@129560.4]
  assign regs_327_clock = clock; // @[:@129569.4]
  assign regs_327_reset = io_reset; // @[:@129570.4 RegFile.scala 76:16:@129577.4]
  assign regs_327_io_in = 64'h0; // @[RegFile.scala 75:16:@129576.4]
  assign regs_327_io_reset = reset; // @[RegFile.scala 78:19:@129580.4]
  assign regs_327_io_enable = 1'h1; // @[RegFile.scala 74:20:@129574.4]
  assign regs_328_clock = clock; // @[:@129583.4]
  assign regs_328_reset = io_reset; // @[:@129584.4 RegFile.scala 76:16:@129591.4]
  assign regs_328_io_in = 64'h0; // @[RegFile.scala 75:16:@129590.4]
  assign regs_328_io_reset = reset; // @[RegFile.scala 78:19:@129594.4]
  assign regs_328_io_enable = 1'h1; // @[RegFile.scala 74:20:@129588.4]
  assign regs_329_clock = clock; // @[:@129597.4]
  assign regs_329_reset = io_reset; // @[:@129598.4 RegFile.scala 76:16:@129605.4]
  assign regs_329_io_in = 64'h0; // @[RegFile.scala 75:16:@129604.4]
  assign regs_329_io_reset = reset; // @[RegFile.scala 78:19:@129608.4]
  assign regs_329_io_enable = 1'h1; // @[RegFile.scala 74:20:@129602.4]
  assign regs_330_clock = clock; // @[:@129611.4]
  assign regs_330_reset = io_reset; // @[:@129612.4 RegFile.scala 76:16:@129619.4]
  assign regs_330_io_in = 64'h0; // @[RegFile.scala 75:16:@129618.4]
  assign regs_330_io_reset = reset; // @[RegFile.scala 78:19:@129622.4]
  assign regs_330_io_enable = 1'h1; // @[RegFile.scala 74:20:@129616.4]
  assign regs_331_clock = clock; // @[:@129625.4]
  assign regs_331_reset = io_reset; // @[:@129626.4 RegFile.scala 76:16:@129633.4]
  assign regs_331_io_in = 64'h0; // @[RegFile.scala 75:16:@129632.4]
  assign regs_331_io_reset = reset; // @[RegFile.scala 78:19:@129636.4]
  assign regs_331_io_enable = 1'h1; // @[RegFile.scala 74:20:@129630.4]
  assign regs_332_clock = clock; // @[:@129639.4]
  assign regs_332_reset = io_reset; // @[:@129640.4 RegFile.scala 76:16:@129647.4]
  assign regs_332_io_in = 64'h0; // @[RegFile.scala 75:16:@129646.4]
  assign regs_332_io_reset = reset; // @[RegFile.scala 78:19:@129650.4]
  assign regs_332_io_enable = 1'h1; // @[RegFile.scala 74:20:@129644.4]
  assign regs_333_clock = clock; // @[:@129653.4]
  assign regs_333_reset = io_reset; // @[:@129654.4 RegFile.scala 76:16:@129661.4]
  assign regs_333_io_in = 64'h0; // @[RegFile.scala 75:16:@129660.4]
  assign regs_333_io_reset = reset; // @[RegFile.scala 78:19:@129664.4]
  assign regs_333_io_enable = 1'h1; // @[RegFile.scala 74:20:@129658.4]
  assign regs_334_clock = clock; // @[:@129667.4]
  assign regs_334_reset = io_reset; // @[:@129668.4 RegFile.scala 76:16:@129675.4]
  assign regs_334_io_in = 64'h0; // @[RegFile.scala 75:16:@129674.4]
  assign regs_334_io_reset = reset; // @[RegFile.scala 78:19:@129678.4]
  assign regs_334_io_enable = 1'h1; // @[RegFile.scala 74:20:@129672.4]
  assign regs_335_clock = clock; // @[:@129681.4]
  assign regs_335_reset = io_reset; // @[:@129682.4 RegFile.scala 76:16:@129689.4]
  assign regs_335_io_in = 64'h0; // @[RegFile.scala 75:16:@129688.4]
  assign regs_335_io_reset = reset; // @[RegFile.scala 78:19:@129692.4]
  assign regs_335_io_enable = 1'h1; // @[RegFile.scala 74:20:@129686.4]
  assign regs_336_clock = clock; // @[:@129695.4]
  assign regs_336_reset = io_reset; // @[:@129696.4 RegFile.scala 76:16:@129703.4]
  assign regs_336_io_in = 64'h0; // @[RegFile.scala 75:16:@129702.4]
  assign regs_336_io_reset = reset; // @[RegFile.scala 78:19:@129706.4]
  assign regs_336_io_enable = 1'h1; // @[RegFile.scala 74:20:@129700.4]
  assign regs_337_clock = clock; // @[:@129709.4]
  assign regs_337_reset = io_reset; // @[:@129710.4 RegFile.scala 76:16:@129717.4]
  assign regs_337_io_in = 64'h0; // @[RegFile.scala 75:16:@129716.4]
  assign regs_337_io_reset = reset; // @[RegFile.scala 78:19:@129720.4]
  assign regs_337_io_enable = 1'h1; // @[RegFile.scala 74:20:@129714.4]
  assign regs_338_clock = clock; // @[:@129723.4]
  assign regs_338_reset = io_reset; // @[:@129724.4 RegFile.scala 76:16:@129731.4]
  assign regs_338_io_in = 64'h0; // @[RegFile.scala 75:16:@129730.4]
  assign regs_338_io_reset = reset; // @[RegFile.scala 78:19:@129734.4]
  assign regs_338_io_enable = 1'h1; // @[RegFile.scala 74:20:@129728.4]
  assign regs_339_clock = clock; // @[:@129737.4]
  assign regs_339_reset = io_reset; // @[:@129738.4 RegFile.scala 76:16:@129745.4]
  assign regs_339_io_in = 64'h0; // @[RegFile.scala 75:16:@129744.4]
  assign regs_339_io_reset = reset; // @[RegFile.scala 78:19:@129748.4]
  assign regs_339_io_enable = 1'h1; // @[RegFile.scala 74:20:@129742.4]
  assign regs_340_clock = clock; // @[:@129751.4]
  assign regs_340_reset = io_reset; // @[:@129752.4 RegFile.scala 76:16:@129759.4]
  assign regs_340_io_in = 64'h0; // @[RegFile.scala 75:16:@129758.4]
  assign regs_340_io_reset = reset; // @[RegFile.scala 78:19:@129762.4]
  assign regs_340_io_enable = 1'h1; // @[RegFile.scala 74:20:@129756.4]
  assign regs_341_clock = clock; // @[:@129765.4]
  assign regs_341_reset = io_reset; // @[:@129766.4 RegFile.scala 76:16:@129773.4]
  assign regs_341_io_in = 64'h0; // @[RegFile.scala 75:16:@129772.4]
  assign regs_341_io_reset = reset; // @[RegFile.scala 78:19:@129776.4]
  assign regs_341_io_enable = 1'h1; // @[RegFile.scala 74:20:@129770.4]
  assign regs_342_clock = clock; // @[:@129779.4]
  assign regs_342_reset = io_reset; // @[:@129780.4 RegFile.scala 76:16:@129787.4]
  assign regs_342_io_in = 64'h0; // @[RegFile.scala 75:16:@129786.4]
  assign regs_342_io_reset = reset; // @[RegFile.scala 78:19:@129790.4]
  assign regs_342_io_enable = 1'h1; // @[RegFile.scala 74:20:@129784.4]
  assign regs_343_clock = clock; // @[:@129793.4]
  assign regs_343_reset = io_reset; // @[:@129794.4 RegFile.scala 76:16:@129801.4]
  assign regs_343_io_in = 64'h0; // @[RegFile.scala 75:16:@129800.4]
  assign regs_343_io_reset = reset; // @[RegFile.scala 78:19:@129804.4]
  assign regs_343_io_enable = 1'h1; // @[RegFile.scala 74:20:@129798.4]
  assign regs_344_clock = clock; // @[:@129807.4]
  assign regs_344_reset = io_reset; // @[:@129808.4 RegFile.scala 76:16:@129815.4]
  assign regs_344_io_in = 64'h0; // @[RegFile.scala 75:16:@129814.4]
  assign regs_344_io_reset = reset; // @[RegFile.scala 78:19:@129818.4]
  assign regs_344_io_enable = 1'h1; // @[RegFile.scala 74:20:@129812.4]
  assign regs_345_clock = clock; // @[:@129821.4]
  assign regs_345_reset = io_reset; // @[:@129822.4 RegFile.scala 76:16:@129829.4]
  assign regs_345_io_in = 64'h0; // @[RegFile.scala 75:16:@129828.4]
  assign regs_345_io_reset = reset; // @[RegFile.scala 78:19:@129832.4]
  assign regs_345_io_enable = 1'h1; // @[RegFile.scala 74:20:@129826.4]
  assign regs_346_clock = clock; // @[:@129835.4]
  assign regs_346_reset = io_reset; // @[:@129836.4 RegFile.scala 76:16:@129843.4]
  assign regs_346_io_in = 64'h0; // @[RegFile.scala 75:16:@129842.4]
  assign regs_346_io_reset = reset; // @[RegFile.scala 78:19:@129846.4]
  assign regs_346_io_enable = 1'h1; // @[RegFile.scala 74:20:@129840.4]
  assign regs_347_clock = clock; // @[:@129849.4]
  assign regs_347_reset = io_reset; // @[:@129850.4 RegFile.scala 76:16:@129857.4]
  assign regs_347_io_in = 64'h0; // @[RegFile.scala 75:16:@129856.4]
  assign regs_347_io_reset = reset; // @[RegFile.scala 78:19:@129860.4]
  assign regs_347_io_enable = 1'h1; // @[RegFile.scala 74:20:@129854.4]
  assign regs_348_clock = clock; // @[:@129863.4]
  assign regs_348_reset = io_reset; // @[:@129864.4 RegFile.scala 76:16:@129871.4]
  assign regs_348_io_in = 64'h0; // @[RegFile.scala 75:16:@129870.4]
  assign regs_348_io_reset = reset; // @[RegFile.scala 78:19:@129874.4]
  assign regs_348_io_enable = 1'h1; // @[RegFile.scala 74:20:@129868.4]
  assign regs_349_clock = clock; // @[:@129877.4]
  assign regs_349_reset = io_reset; // @[:@129878.4 RegFile.scala 76:16:@129885.4]
  assign regs_349_io_in = 64'h0; // @[RegFile.scala 75:16:@129884.4]
  assign regs_349_io_reset = reset; // @[RegFile.scala 78:19:@129888.4]
  assign regs_349_io_enable = 1'h1; // @[RegFile.scala 74:20:@129882.4]
  assign regs_350_clock = clock; // @[:@129891.4]
  assign regs_350_reset = io_reset; // @[:@129892.4 RegFile.scala 76:16:@129899.4]
  assign regs_350_io_in = 64'h0; // @[RegFile.scala 75:16:@129898.4]
  assign regs_350_io_reset = reset; // @[RegFile.scala 78:19:@129902.4]
  assign regs_350_io_enable = 1'h1; // @[RegFile.scala 74:20:@129896.4]
  assign regs_351_clock = clock; // @[:@129905.4]
  assign regs_351_reset = io_reset; // @[:@129906.4 RegFile.scala 76:16:@129913.4]
  assign regs_351_io_in = 64'h0; // @[RegFile.scala 75:16:@129912.4]
  assign regs_351_io_reset = reset; // @[RegFile.scala 78:19:@129916.4]
  assign regs_351_io_enable = 1'h1; // @[RegFile.scala 74:20:@129910.4]
  assign regs_352_clock = clock; // @[:@129919.4]
  assign regs_352_reset = io_reset; // @[:@129920.4 RegFile.scala 76:16:@129927.4]
  assign regs_352_io_in = 64'h0; // @[RegFile.scala 75:16:@129926.4]
  assign regs_352_io_reset = reset; // @[RegFile.scala 78:19:@129930.4]
  assign regs_352_io_enable = 1'h1; // @[RegFile.scala 74:20:@129924.4]
  assign regs_353_clock = clock; // @[:@129933.4]
  assign regs_353_reset = io_reset; // @[:@129934.4 RegFile.scala 76:16:@129941.4]
  assign regs_353_io_in = 64'h0; // @[RegFile.scala 75:16:@129940.4]
  assign regs_353_io_reset = reset; // @[RegFile.scala 78:19:@129944.4]
  assign regs_353_io_enable = 1'h1; // @[RegFile.scala 74:20:@129938.4]
  assign regs_354_clock = clock; // @[:@129947.4]
  assign regs_354_reset = io_reset; // @[:@129948.4 RegFile.scala 76:16:@129955.4]
  assign regs_354_io_in = 64'h0; // @[RegFile.scala 75:16:@129954.4]
  assign regs_354_io_reset = reset; // @[RegFile.scala 78:19:@129958.4]
  assign regs_354_io_enable = 1'h1; // @[RegFile.scala 74:20:@129952.4]
  assign regs_355_clock = clock; // @[:@129961.4]
  assign regs_355_reset = io_reset; // @[:@129962.4 RegFile.scala 76:16:@129969.4]
  assign regs_355_io_in = 64'h0; // @[RegFile.scala 75:16:@129968.4]
  assign regs_355_io_reset = reset; // @[RegFile.scala 78:19:@129972.4]
  assign regs_355_io_enable = 1'h1; // @[RegFile.scala 74:20:@129966.4]
  assign regs_356_clock = clock; // @[:@129975.4]
  assign regs_356_reset = io_reset; // @[:@129976.4 RegFile.scala 76:16:@129983.4]
  assign regs_356_io_in = 64'h0; // @[RegFile.scala 75:16:@129982.4]
  assign regs_356_io_reset = reset; // @[RegFile.scala 78:19:@129986.4]
  assign regs_356_io_enable = 1'h1; // @[RegFile.scala 74:20:@129980.4]
  assign regs_357_clock = clock; // @[:@129989.4]
  assign regs_357_reset = io_reset; // @[:@129990.4 RegFile.scala 76:16:@129997.4]
  assign regs_357_io_in = 64'h0; // @[RegFile.scala 75:16:@129996.4]
  assign regs_357_io_reset = reset; // @[RegFile.scala 78:19:@130000.4]
  assign regs_357_io_enable = 1'h1; // @[RegFile.scala 74:20:@129994.4]
  assign regs_358_clock = clock; // @[:@130003.4]
  assign regs_358_reset = io_reset; // @[:@130004.4 RegFile.scala 76:16:@130011.4]
  assign regs_358_io_in = 64'h0; // @[RegFile.scala 75:16:@130010.4]
  assign regs_358_io_reset = reset; // @[RegFile.scala 78:19:@130014.4]
  assign regs_358_io_enable = 1'h1; // @[RegFile.scala 74:20:@130008.4]
  assign regs_359_clock = clock; // @[:@130017.4]
  assign regs_359_reset = io_reset; // @[:@130018.4 RegFile.scala 76:16:@130025.4]
  assign regs_359_io_in = 64'h0; // @[RegFile.scala 75:16:@130024.4]
  assign regs_359_io_reset = reset; // @[RegFile.scala 78:19:@130028.4]
  assign regs_359_io_enable = 1'h1; // @[RegFile.scala 74:20:@130022.4]
  assign regs_360_clock = clock; // @[:@130031.4]
  assign regs_360_reset = io_reset; // @[:@130032.4 RegFile.scala 76:16:@130039.4]
  assign regs_360_io_in = 64'h0; // @[RegFile.scala 75:16:@130038.4]
  assign regs_360_io_reset = reset; // @[RegFile.scala 78:19:@130042.4]
  assign regs_360_io_enable = 1'h1; // @[RegFile.scala 74:20:@130036.4]
  assign regs_361_clock = clock; // @[:@130045.4]
  assign regs_361_reset = io_reset; // @[:@130046.4 RegFile.scala 76:16:@130053.4]
  assign regs_361_io_in = 64'h0; // @[RegFile.scala 75:16:@130052.4]
  assign regs_361_io_reset = reset; // @[RegFile.scala 78:19:@130056.4]
  assign regs_361_io_enable = 1'h1; // @[RegFile.scala 74:20:@130050.4]
  assign regs_362_clock = clock; // @[:@130059.4]
  assign regs_362_reset = io_reset; // @[:@130060.4 RegFile.scala 76:16:@130067.4]
  assign regs_362_io_in = 64'h0; // @[RegFile.scala 75:16:@130066.4]
  assign regs_362_io_reset = reset; // @[RegFile.scala 78:19:@130070.4]
  assign regs_362_io_enable = 1'h1; // @[RegFile.scala 74:20:@130064.4]
  assign regs_363_clock = clock; // @[:@130073.4]
  assign regs_363_reset = io_reset; // @[:@130074.4 RegFile.scala 76:16:@130081.4]
  assign regs_363_io_in = 64'h0; // @[RegFile.scala 75:16:@130080.4]
  assign regs_363_io_reset = reset; // @[RegFile.scala 78:19:@130084.4]
  assign regs_363_io_enable = 1'h1; // @[RegFile.scala 74:20:@130078.4]
  assign regs_364_clock = clock; // @[:@130087.4]
  assign regs_364_reset = io_reset; // @[:@130088.4 RegFile.scala 76:16:@130095.4]
  assign regs_364_io_in = 64'h0; // @[RegFile.scala 75:16:@130094.4]
  assign regs_364_io_reset = reset; // @[RegFile.scala 78:19:@130098.4]
  assign regs_364_io_enable = 1'h1; // @[RegFile.scala 74:20:@130092.4]
  assign regs_365_clock = clock; // @[:@130101.4]
  assign regs_365_reset = io_reset; // @[:@130102.4 RegFile.scala 76:16:@130109.4]
  assign regs_365_io_in = 64'h0; // @[RegFile.scala 75:16:@130108.4]
  assign regs_365_io_reset = reset; // @[RegFile.scala 78:19:@130112.4]
  assign regs_365_io_enable = 1'h1; // @[RegFile.scala 74:20:@130106.4]
  assign regs_366_clock = clock; // @[:@130115.4]
  assign regs_366_reset = io_reset; // @[:@130116.4 RegFile.scala 76:16:@130123.4]
  assign regs_366_io_in = 64'h0; // @[RegFile.scala 75:16:@130122.4]
  assign regs_366_io_reset = reset; // @[RegFile.scala 78:19:@130126.4]
  assign regs_366_io_enable = 1'h1; // @[RegFile.scala 74:20:@130120.4]
  assign regs_367_clock = clock; // @[:@130129.4]
  assign regs_367_reset = io_reset; // @[:@130130.4 RegFile.scala 76:16:@130137.4]
  assign regs_367_io_in = 64'h0; // @[RegFile.scala 75:16:@130136.4]
  assign regs_367_io_reset = reset; // @[RegFile.scala 78:19:@130140.4]
  assign regs_367_io_enable = 1'h1; // @[RegFile.scala 74:20:@130134.4]
  assign regs_368_clock = clock; // @[:@130143.4]
  assign regs_368_reset = io_reset; // @[:@130144.4 RegFile.scala 76:16:@130151.4]
  assign regs_368_io_in = 64'h0; // @[RegFile.scala 75:16:@130150.4]
  assign regs_368_io_reset = reset; // @[RegFile.scala 78:19:@130154.4]
  assign regs_368_io_enable = 1'h1; // @[RegFile.scala 74:20:@130148.4]
  assign regs_369_clock = clock; // @[:@130157.4]
  assign regs_369_reset = io_reset; // @[:@130158.4 RegFile.scala 76:16:@130165.4]
  assign regs_369_io_in = 64'h0; // @[RegFile.scala 75:16:@130164.4]
  assign regs_369_io_reset = reset; // @[RegFile.scala 78:19:@130168.4]
  assign regs_369_io_enable = 1'h1; // @[RegFile.scala 74:20:@130162.4]
  assign regs_370_clock = clock; // @[:@130171.4]
  assign regs_370_reset = io_reset; // @[:@130172.4 RegFile.scala 76:16:@130179.4]
  assign regs_370_io_in = 64'h0; // @[RegFile.scala 75:16:@130178.4]
  assign regs_370_io_reset = reset; // @[RegFile.scala 78:19:@130182.4]
  assign regs_370_io_enable = 1'h1; // @[RegFile.scala 74:20:@130176.4]
  assign regs_371_clock = clock; // @[:@130185.4]
  assign regs_371_reset = io_reset; // @[:@130186.4 RegFile.scala 76:16:@130193.4]
  assign regs_371_io_in = 64'h0; // @[RegFile.scala 75:16:@130192.4]
  assign regs_371_io_reset = reset; // @[RegFile.scala 78:19:@130196.4]
  assign regs_371_io_enable = 1'h1; // @[RegFile.scala 74:20:@130190.4]
  assign regs_372_clock = clock; // @[:@130199.4]
  assign regs_372_reset = io_reset; // @[:@130200.4 RegFile.scala 76:16:@130207.4]
  assign regs_372_io_in = 64'h0; // @[RegFile.scala 75:16:@130206.4]
  assign regs_372_io_reset = reset; // @[RegFile.scala 78:19:@130210.4]
  assign regs_372_io_enable = 1'h1; // @[RegFile.scala 74:20:@130204.4]
  assign regs_373_clock = clock; // @[:@130213.4]
  assign regs_373_reset = io_reset; // @[:@130214.4 RegFile.scala 76:16:@130221.4]
  assign regs_373_io_in = 64'h0; // @[RegFile.scala 75:16:@130220.4]
  assign regs_373_io_reset = reset; // @[RegFile.scala 78:19:@130224.4]
  assign regs_373_io_enable = 1'h1; // @[RegFile.scala 74:20:@130218.4]
  assign regs_374_clock = clock; // @[:@130227.4]
  assign regs_374_reset = io_reset; // @[:@130228.4 RegFile.scala 76:16:@130235.4]
  assign regs_374_io_in = 64'h0; // @[RegFile.scala 75:16:@130234.4]
  assign regs_374_io_reset = reset; // @[RegFile.scala 78:19:@130238.4]
  assign regs_374_io_enable = 1'h1; // @[RegFile.scala 74:20:@130232.4]
  assign regs_375_clock = clock; // @[:@130241.4]
  assign regs_375_reset = io_reset; // @[:@130242.4 RegFile.scala 76:16:@130249.4]
  assign regs_375_io_in = 64'h0; // @[RegFile.scala 75:16:@130248.4]
  assign regs_375_io_reset = reset; // @[RegFile.scala 78:19:@130252.4]
  assign regs_375_io_enable = 1'h1; // @[RegFile.scala 74:20:@130246.4]
  assign regs_376_clock = clock; // @[:@130255.4]
  assign regs_376_reset = io_reset; // @[:@130256.4 RegFile.scala 76:16:@130263.4]
  assign regs_376_io_in = 64'h0; // @[RegFile.scala 75:16:@130262.4]
  assign regs_376_io_reset = reset; // @[RegFile.scala 78:19:@130266.4]
  assign regs_376_io_enable = 1'h1; // @[RegFile.scala 74:20:@130260.4]
  assign regs_377_clock = clock; // @[:@130269.4]
  assign regs_377_reset = io_reset; // @[:@130270.4 RegFile.scala 76:16:@130277.4]
  assign regs_377_io_in = 64'h0; // @[RegFile.scala 75:16:@130276.4]
  assign regs_377_io_reset = reset; // @[RegFile.scala 78:19:@130280.4]
  assign regs_377_io_enable = 1'h1; // @[RegFile.scala 74:20:@130274.4]
  assign regs_378_clock = clock; // @[:@130283.4]
  assign regs_378_reset = io_reset; // @[:@130284.4 RegFile.scala 76:16:@130291.4]
  assign regs_378_io_in = 64'h0; // @[RegFile.scala 75:16:@130290.4]
  assign regs_378_io_reset = reset; // @[RegFile.scala 78:19:@130294.4]
  assign regs_378_io_enable = 1'h1; // @[RegFile.scala 74:20:@130288.4]
  assign regs_379_clock = clock; // @[:@130297.4]
  assign regs_379_reset = io_reset; // @[:@130298.4 RegFile.scala 76:16:@130305.4]
  assign regs_379_io_in = 64'h0; // @[RegFile.scala 75:16:@130304.4]
  assign regs_379_io_reset = reset; // @[RegFile.scala 78:19:@130308.4]
  assign regs_379_io_enable = 1'h1; // @[RegFile.scala 74:20:@130302.4]
  assign regs_380_clock = clock; // @[:@130311.4]
  assign regs_380_reset = io_reset; // @[:@130312.4 RegFile.scala 76:16:@130319.4]
  assign regs_380_io_in = 64'h0; // @[RegFile.scala 75:16:@130318.4]
  assign regs_380_io_reset = reset; // @[RegFile.scala 78:19:@130322.4]
  assign regs_380_io_enable = 1'h1; // @[RegFile.scala 74:20:@130316.4]
  assign regs_381_clock = clock; // @[:@130325.4]
  assign regs_381_reset = io_reset; // @[:@130326.4 RegFile.scala 76:16:@130333.4]
  assign regs_381_io_in = 64'h0; // @[RegFile.scala 75:16:@130332.4]
  assign regs_381_io_reset = reset; // @[RegFile.scala 78:19:@130336.4]
  assign regs_381_io_enable = 1'h1; // @[RegFile.scala 74:20:@130330.4]
  assign regs_382_clock = clock; // @[:@130339.4]
  assign regs_382_reset = io_reset; // @[:@130340.4 RegFile.scala 76:16:@130347.4]
  assign regs_382_io_in = 64'h0; // @[RegFile.scala 75:16:@130346.4]
  assign regs_382_io_reset = reset; // @[RegFile.scala 78:19:@130350.4]
  assign regs_382_io_enable = 1'h1; // @[RegFile.scala 74:20:@130344.4]
  assign regs_383_clock = clock; // @[:@130353.4]
  assign regs_383_reset = io_reset; // @[:@130354.4 RegFile.scala 76:16:@130361.4]
  assign regs_383_io_in = 64'h0; // @[RegFile.scala 75:16:@130360.4]
  assign regs_383_io_reset = reset; // @[RegFile.scala 78:19:@130364.4]
  assign regs_383_io_enable = 1'h1; // @[RegFile.scala 74:20:@130358.4]
  assign regs_384_clock = clock; // @[:@130367.4]
  assign regs_384_reset = io_reset; // @[:@130368.4 RegFile.scala 76:16:@130375.4]
  assign regs_384_io_in = 64'h0; // @[RegFile.scala 75:16:@130374.4]
  assign regs_384_io_reset = reset; // @[RegFile.scala 78:19:@130378.4]
  assign regs_384_io_enable = 1'h1; // @[RegFile.scala 74:20:@130372.4]
  assign regs_385_clock = clock; // @[:@130381.4]
  assign regs_385_reset = io_reset; // @[:@130382.4 RegFile.scala 76:16:@130389.4]
  assign regs_385_io_in = 64'h0; // @[RegFile.scala 75:16:@130388.4]
  assign regs_385_io_reset = reset; // @[RegFile.scala 78:19:@130392.4]
  assign regs_385_io_enable = 1'h1; // @[RegFile.scala 74:20:@130386.4]
  assign regs_386_clock = clock; // @[:@130395.4]
  assign regs_386_reset = io_reset; // @[:@130396.4 RegFile.scala 76:16:@130403.4]
  assign regs_386_io_in = 64'h0; // @[RegFile.scala 75:16:@130402.4]
  assign regs_386_io_reset = reset; // @[RegFile.scala 78:19:@130406.4]
  assign regs_386_io_enable = 1'h1; // @[RegFile.scala 74:20:@130400.4]
  assign regs_387_clock = clock; // @[:@130409.4]
  assign regs_387_reset = io_reset; // @[:@130410.4 RegFile.scala 76:16:@130417.4]
  assign regs_387_io_in = 64'h0; // @[RegFile.scala 75:16:@130416.4]
  assign regs_387_io_reset = reset; // @[RegFile.scala 78:19:@130420.4]
  assign regs_387_io_enable = 1'h1; // @[RegFile.scala 74:20:@130414.4]
  assign regs_388_clock = clock; // @[:@130423.4]
  assign regs_388_reset = io_reset; // @[:@130424.4 RegFile.scala 76:16:@130431.4]
  assign regs_388_io_in = 64'h0; // @[RegFile.scala 75:16:@130430.4]
  assign regs_388_io_reset = reset; // @[RegFile.scala 78:19:@130434.4]
  assign regs_388_io_enable = 1'h1; // @[RegFile.scala 74:20:@130428.4]
  assign regs_389_clock = clock; // @[:@130437.4]
  assign regs_389_reset = io_reset; // @[:@130438.4 RegFile.scala 76:16:@130445.4]
  assign regs_389_io_in = 64'h0; // @[RegFile.scala 75:16:@130444.4]
  assign regs_389_io_reset = reset; // @[RegFile.scala 78:19:@130448.4]
  assign regs_389_io_enable = 1'h1; // @[RegFile.scala 74:20:@130442.4]
  assign regs_390_clock = clock; // @[:@130451.4]
  assign regs_390_reset = io_reset; // @[:@130452.4 RegFile.scala 76:16:@130459.4]
  assign regs_390_io_in = 64'h0; // @[RegFile.scala 75:16:@130458.4]
  assign regs_390_io_reset = reset; // @[RegFile.scala 78:19:@130462.4]
  assign regs_390_io_enable = 1'h1; // @[RegFile.scala 74:20:@130456.4]
  assign regs_391_clock = clock; // @[:@130465.4]
  assign regs_391_reset = io_reset; // @[:@130466.4 RegFile.scala 76:16:@130473.4]
  assign regs_391_io_in = 64'h0; // @[RegFile.scala 75:16:@130472.4]
  assign regs_391_io_reset = reset; // @[RegFile.scala 78:19:@130476.4]
  assign regs_391_io_enable = 1'h1; // @[RegFile.scala 74:20:@130470.4]
  assign regs_392_clock = clock; // @[:@130479.4]
  assign regs_392_reset = io_reset; // @[:@130480.4 RegFile.scala 76:16:@130487.4]
  assign regs_392_io_in = 64'h0; // @[RegFile.scala 75:16:@130486.4]
  assign regs_392_io_reset = reset; // @[RegFile.scala 78:19:@130490.4]
  assign regs_392_io_enable = 1'h1; // @[RegFile.scala 74:20:@130484.4]
  assign regs_393_clock = clock; // @[:@130493.4]
  assign regs_393_reset = io_reset; // @[:@130494.4 RegFile.scala 76:16:@130501.4]
  assign regs_393_io_in = 64'h0; // @[RegFile.scala 75:16:@130500.4]
  assign regs_393_io_reset = reset; // @[RegFile.scala 78:19:@130504.4]
  assign regs_393_io_enable = 1'h1; // @[RegFile.scala 74:20:@130498.4]
  assign regs_394_clock = clock; // @[:@130507.4]
  assign regs_394_reset = io_reset; // @[:@130508.4 RegFile.scala 76:16:@130515.4]
  assign regs_394_io_in = 64'h0; // @[RegFile.scala 75:16:@130514.4]
  assign regs_394_io_reset = reset; // @[RegFile.scala 78:19:@130518.4]
  assign regs_394_io_enable = 1'h1; // @[RegFile.scala 74:20:@130512.4]
  assign regs_395_clock = clock; // @[:@130521.4]
  assign regs_395_reset = io_reset; // @[:@130522.4 RegFile.scala 76:16:@130529.4]
  assign regs_395_io_in = 64'h0; // @[RegFile.scala 75:16:@130528.4]
  assign regs_395_io_reset = reset; // @[RegFile.scala 78:19:@130532.4]
  assign regs_395_io_enable = 1'h1; // @[RegFile.scala 74:20:@130526.4]
  assign regs_396_clock = clock; // @[:@130535.4]
  assign regs_396_reset = io_reset; // @[:@130536.4 RegFile.scala 76:16:@130543.4]
  assign regs_396_io_in = 64'h0; // @[RegFile.scala 75:16:@130542.4]
  assign regs_396_io_reset = reset; // @[RegFile.scala 78:19:@130546.4]
  assign regs_396_io_enable = 1'h1; // @[RegFile.scala 74:20:@130540.4]
  assign regs_397_clock = clock; // @[:@130549.4]
  assign regs_397_reset = io_reset; // @[:@130550.4 RegFile.scala 76:16:@130557.4]
  assign regs_397_io_in = 64'h0; // @[RegFile.scala 75:16:@130556.4]
  assign regs_397_io_reset = reset; // @[RegFile.scala 78:19:@130560.4]
  assign regs_397_io_enable = 1'h1; // @[RegFile.scala 74:20:@130554.4]
  assign regs_398_clock = clock; // @[:@130563.4]
  assign regs_398_reset = io_reset; // @[:@130564.4 RegFile.scala 76:16:@130571.4]
  assign regs_398_io_in = 64'h0; // @[RegFile.scala 75:16:@130570.4]
  assign regs_398_io_reset = reset; // @[RegFile.scala 78:19:@130574.4]
  assign regs_398_io_enable = 1'h1; // @[RegFile.scala 74:20:@130568.4]
  assign regs_399_clock = clock; // @[:@130577.4]
  assign regs_399_reset = io_reset; // @[:@130578.4 RegFile.scala 76:16:@130585.4]
  assign regs_399_io_in = 64'h0; // @[RegFile.scala 75:16:@130584.4]
  assign regs_399_io_reset = reset; // @[RegFile.scala 78:19:@130588.4]
  assign regs_399_io_enable = 1'h1; // @[RegFile.scala 74:20:@130582.4]
  assign regs_400_clock = clock; // @[:@130591.4]
  assign regs_400_reset = io_reset; // @[:@130592.4 RegFile.scala 76:16:@130599.4]
  assign regs_400_io_in = 64'h0; // @[RegFile.scala 75:16:@130598.4]
  assign regs_400_io_reset = reset; // @[RegFile.scala 78:19:@130602.4]
  assign regs_400_io_enable = 1'h1; // @[RegFile.scala 74:20:@130596.4]
  assign regs_401_clock = clock; // @[:@130605.4]
  assign regs_401_reset = io_reset; // @[:@130606.4 RegFile.scala 76:16:@130613.4]
  assign regs_401_io_in = 64'h0; // @[RegFile.scala 75:16:@130612.4]
  assign regs_401_io_reset = reset; // @[RegFile.scala 78:19:@130616.4]
  assign regs_401_io_enable = 1'h1; // @[RegFile.scala 74:20:@130610.4]
  assign regs_402_clock = clock; // @[:@130619.4]
  assign regs_402_reset = io_reset; // @[:@130620.4 RegFile.scala 76:16:@130627.4]
  assign regs_402_io_in = 64'h0; // @[RegFile.scala 75:16:@130626.4]
  assign regs_402_io_reset = reset; // @[RegFile.scala 78:19:@130630.4]
  assign regs_402_io_enable = 1'h1; // @[RegFile.scala 74:20:@130624.4]
  assign regs_403_clock = clock; // @[:@130633.4]
  assign regs_403_reset = io_reset; // @[:@130634.4 RegFile.scala 76:16:@130641.4]
  assign regs_403_io_in = 64'h0; // @[RegFile.scala 75:16:@130640.4]
  assign regs_403_io_reset = reset; // @[RegFile.scala 78:19:@130644.4]
  assign regs_403_io_enable = 1'h1; // @[RegFile.scala 74:20:@130638.4]
  assign regs_404_clock = clock; // @[:@130647.4]
  assign regs_404_reset = io_reset; // @[:@130648.4 RegFile.scala 76:16:@130655.4]
  assign regs_404_io_in = 64'h0; // @[RegFile.scala 75:16:@130654.4]
  assign regs_404_io_reset = reset; // @[RegFile.scala 78:19:@130658.4]
  assign regs_404_io_enable = 1'h1; // @[RegFile.scala 74:20:@130652.4]
  assign regs_405_clock = clock; // @[:@130661.4]
  assign regs_405_reset = io_reset; // @[:@130662.4 RegFile.scala 76:16:@130669.4]
  assign regs_405_io_in = 64'h0; // @[RegFile.scala 75:16:@130668.4]
  assign regs_405_io_reset = reset; // @[RegFile.scala 78:19:@130672.4]
  assign regs_405_io_enable = 1'h1; // @[RegFile.scala 74:20:@130666.4]
  assign regs_406_clock = clock; // @[:@130675.4]
  assign regs_406_reset = io_reset; // @[:@130676.4 RegFile.scala 76:16:@130683.4]
  assign regs_406_io_in = 64'h0; // @[RegFile.scala 75:16:@130682.4]
  assign regs_406_io_reset = reset; // @[RegFile.scala 78:19:@130686.4]
  assign regs_406_io_enable = 1'h1; // @[RegFile.scala 74:20:@130680.4]
  assign regs_407_clock = clock; // @[:@130689.4]
  assign regs_407_reset = io_reset; // @[:@130690.4 RegFile.scala 76:16:@130697.4]
  assign regs_407_io_in = 64'h0; // @[RegFile.scala 75:16:@130696.4]
  assign regs_407_io_reset = reset; // @[RegFile.scala 78:19:@130700.4]
  assign regs_407_io_enable = 1'h1; // @[RegFile.scala 74:20:@130694.4]
  assign regs_408_clock = clock; // @[:@130703.4]
  assign regs_408_reset = io_reset; // @[:@130704.4 RegFile.scala 76:16:@130711.4]
  assign regs_408_io_in = 64'h0; // @[RegFile.scala 75:16:@130710.4]
  assign regs_408_io_reset = reset; // @[RegFile.scala 78:19:@130714.4]
  assign regs_408_io_enable = 1'h1; // @[RegFile.scala 74:20:@130708.4]
  assign regs_409_clock = clock; // @[:@130717.4]
  assign regs_409_reset = io_reset; // @[:@130718.4 RegFile.scala 76:16:@130725.4]
  assign regs_409_io_in = 64'h0; // @[RegFile.scala 75:16:@130724.4]
  assign regs_409_io_reset = reset; // @[RegFile.scala 78:19:@130728.4]
  assign regs_409_io_enable = 1'h1; // @[RegFile.scala 74:20:@130722.4]
  assign regs_410_clock = clock; // @[:@130731.4]
  assign regs_410_reset = io_reset; // @[:@130732.4 RegFile.scala 76:16:@130739.4]
  assign regs_410_io_in = 64'h0; // @[RegFile.scala 75:16:@130738.4]
  assign regs_410_io_reset = reset; // @[RegFile.scala 78:19:@130742.4]
  assign regs_410_io_enable = 1'h1; // @[RegFile.scala 74:20:@130736.4]
  assign regs_411_clock = clock; // @[:@130745.4]
  assign regs_411_reset = io_reset; // @[:@130746.4 RegFile.scala 76:16:@130753.4]
  assign regs_411_io_in = 64'h0; // @[RegFile.scala 75:16:@130752.4]
  assign regs_411_io_reset = reset; // @[RegFile.scala 78:19:@130756.4]
  assign regs_411_io_enable = 1'h1; // @[RegFile.scala 74:20:@130750.4]
  assign regs_412_clock = clock; // @[:@130759.4]
  assign regs_412_reset = io_reset; // @[:@130760.4 RegFile.scala 76:16:@130767.4]
  assign regs_412_io_in = 64'h0; // @[RegFile.scala 75:16:@130766.4]
  assign regs_412_io_reset = reset; // @[RegFile.scala 78:19:@130770.4]
  assign regs_412_io_enable = 1'h1; // @[RegFile.scala 74:20:@130764.4]
  assign regs_413_clock = clock; // @[:@130773.4]
  assign regs_413_reset = io_reset; // @[:@130774.4 RegFile.scala 76:16:@130781.4]
  assign regs_413_io_in = 64'h0; // @[RegFile.scala 75:16:@130780.4]
  assign regs_413_io_reset = reset; // @[RegFile.scala 78:19:@130784.4]
  assign regs_413_io_enable = 1'h1; // @[RegFile.scala 74:20:@130778.4]
  assign regs_414_clock = clock; // @[:@130787.4]
  assign regs_414_reset = io_reset; // @[:@130788.4 RegFile.scala 76:16:@130795.4]
  assign regs_414_io_in = 64'h0; // @[RegFile.scala 75:16:@130794.4]
  assign regs_414_io_reset = reset; // @[RegFile.scala 78:19:@130798.4]
  assign regs_414_io_enable = 1'h1; // @[RegFile.scala 74:20:@130792.4]
  assign regs_415_clock = clock; // @[:@130801.4]
  assign regs_415_reset = io_reset; // @[:@130802.4 RegFile.scala 76:16:@130809.4]
  assign regs_415_io_in = 64'h0; // @[RegFile.scala 75:16:@130808.4]
  assign regs_415_io_reset = reset; // @[RegFile.scala 78:19:@130812.4]
  assign regs_415_io_enable = 1'h1; // @[RegFile.scala 74:20:@130806.4]
  assign regs_416_clock = clock; // @[:@130815.4]
  assign regs_416_reset = io_reset; // @[:@130816.4 RegFile.scala 76:16:@130823.4]
  assign regs_416_io_in = 64'h0; // @[RegFile.scala 75:16:@130822.4]
  assign regs_416_io_reset = reset; // @[RegFile.scala 78:19:@130826.4]
  assign regs_416_io_enable = 1'h1; // @[RegFile.scala 74:20:@130820.4]
  assign regs_417_clock = clock; // @[:@130829.4]
  assign regs_417_reset = io_reset; // @[:@130830.4 RegFile.scala 76:16:@130837.4]
  assign regs_417_io_in = 64'h0; // @[RegFile.scala 75:16:@130836.4]
  assign regs_417_io_reset = reset; // @[RegFile.scala 78:19:@130840.4]
  assign regs_417_io_enable = 1'h1; // @[RegFile.scala 74:20:@130834.4]
  assign regs_418_clock = clock; // @[:@130843.4]
  assign regs_418_reset = io_reset; // @[:@130844.4 RegFile.scala 76:16:@130851.4]
  assign regs_418_io_in = 64'h0; // @[RegFile.scala 75:16:@130850.4]
  assign regs_418_io_reset = reset; // @[RegFile.scala 78:19:@130854.4]
  assign regs_418_io_enable = 1'h1; // @[RegFile.scala 74:20:@130848.4]
  assign regs_419_clock = clock; // @[:@130857.4]
  assign regs_419_reset = io_reset; // @[:@130858.4 RegFile.scala 76:16:@130865.4]
  assign regs_419_io_in = 64'h0; // @[RegFile.scala 75:16:@130864.4]
  assign regs_419_io_reset = reset; // @[RegFile.scala 78:19:@130868.4]
  assign regs_419_io_enable = 1'h1; // @[RegFile.scala 74:20:@130862.4]
  assign regs_420_clock = clock; // @[:@130871.4]
  assign regs_420_reset = io_reset; // @[:@130872.4 RegFile.scala 76:16:@130879.4]
  assign regs_420_io_in = 64'h0; // @[RegFile.scala 75:16:@130878.4]
  assign regs_420_io_reset = reset; // @[RegFile.scala 78:19:@130882.4]
  assign regs_420_io_enable = 1'h1; // @[RegFile.scala 74:20:@130876.4]
  assign regs_421_clock = clock; // @[:@130885.4]
  assign regs_421_reset = io_reset; // @[:@130886.4 RegFile.scala 76:16:@130893.4]
  assign regs_421_io_in = 64'h0; // @[RegFile.scala 75:16:@130892.4]
  assign regs_421_io_reset = reset; // @[RegFile.scala 78:19:@130896.4]
  assign regs_421_io_enable = 1'h1; // @[RegFile.scala 74:20:@130890.4]
  assign regs_422_clock = clock; // @[:@130899.4]
  assign regs_422_reset = io_reset; // @[:@130900.4 RegFile.scala 76:16:@130907.4]
  assign regs_422_io_in = 64'h0; // @[RegFile.scala 75:16:@130906.4]
  assign regs_422_io_reset = reset; // @[RegFile.scala 78:19:@130910.4]
  assign regs_422_io_enable = 1'h1; // @[RegFile.scala 74:20:@130904.4]
  assign regs_423_clock = clock; // @[:@130913.4]
  assign regs_423_reset = io_reset; // @[:@130914.4 RegFile.scala 76:16:@130921.4]
  assign regs_423_io_in = 64'h0; // @[RegFile.scala 75:16:@130920.4]
  assign regs_423_io_reset = reset; // @[RegFile.scala 78:19:@130924.4]
  assign regs_423_io_enable = 1'h1; // @[RegFile.scala 74:20:@130918.4]
  assign regs_424_clock = clock; // @[:@130927.4]
  assign regs_424_reset = io_reset; // @[:@130928.4 RegFile.scala 76:16:@130935.4]
  assign regs_424_io_in = 64'h0; // @[RegFile.scala 75:16:@130934.4]
  assign regs_424_io_reset = reset; // @[RegFile.scala 78:19:@130938.4]
  assign regs_424_io_enable = 1'h1; // @[RegFile.scala 74:20:@130932.4]
  assign regs_425_clock = clock; // @[:@130941.4]
  assign regs_425_reset = io_reset; // @[:@130942.4 RegFile.scala 76:16:@130949.4]
  assign regs_425_io_in = 64'h0; // @[RegFile.scala 75:16:@130948.4]
  assign regs_425_io_reset = reset; // @[RegFile.scala 78:19:@130952.4]
  assign regs_425_io_enable = 1'h1; // @[RegFile.scala 74:20:@130946.4]
  assign regs_426_clock = clock; // @[:@130955.4]
  assign regs_426_reset = io_reset; // @[:@130956.4 RegFile.scala 76:16:@130963.4]
  assign regs_426_io_in = 64'h0; // @[RegFile.scala 75:16:@130962.4]
  assign regs_426_io_reset = reset; // @[RegFile.scala 78:19:@130966.4]
  assign regs_426_io_enable = 1'h1; // @[RegFile.scala 74:20:@130960.4]
  assign regs_427_clock = clock; // @[:@130969.4]
  assign regs_427_reset = io_reset; // @[:@130970.4 RegFile.scala 76:16:@130977.4]
  assign regs_427_io_in = 64'h0; // @[RegFile.scala 75:16:@130976.4]
  assign regs_427_io_reset = reset; // @[RegFile.scala 78:19:@130980.4]
  assign regs_427_io_enable = 1'h1; // @[RegFile.scala 74:20:@130974.4]
  assign regs_428_clock = clock; // @[:@130983.4]
  assign regs_428_reset = io_reset; // @[:@130984.4 RegFile.scala 76:16:@130991.4]
  assign regs_428_io_in = 64'h0; // @[RegFile.scala 75:16:@130990.4]
  assign regs_428_io_reset = reset; // @[RegFile.scala 78:19:@130994.4]
  assign regs_428_io_enable = 1'h1; // @[RegFile.scala 74:20:@130988.4]
  assign regs_429_clock = clock; // @[:@130997.4]
  assign regs_429_reset = io_reset; // @[:@130998.4 RegFile.scala 76:16:@131005.4]
  assign regs_429_io_in = 64'h0; // @[RegFile.scala 75:16:@131004.4]
  assign regs_429_io_reset = reset; // @[RegFile.scala 78:19:@131008.4]
  assign regs_429_io_enable = 1'h1; // @[RegFile.scala 74:20:@131002.4]
  assign regs_430_clock = clock; // @[:@131011.4]
  assign regs_430_reset = io_reset; // @[:@131012.4 RegFile.scala 76:16:@131019.4]
  assign regs_430_io_in = 64'h0; // @[RegFile.scala 75:16:@131018.4]
  assign regs_430_io_reset = reset; // @[RegFile.scala 78:19:@131022.4]
  assign regs_430_io_enable = 1'h1; // @[RegFile.scala 74:20:@131016.4]
  assign regs_431_clock = clock; // @[:@131025.4]
  assign regs_431_reset = io_reset; // @[:@131026.4 RegFile.scala 76:16:@131033.4]
  assign regs_431_io_in = 64'h0; // @[RegFile.scala 75:16:@131032.4]
  assign regs_431_io_reset = reset; // @[RegFile.scala 78:19:@131036.4]
  assign regs_431_io_enable = 1'h1; // @[RegFile.scala 74:20:@131030.4]
  assign regs_432_clock = clock; // @[:@131039.4]
  assign regs_432_reset = io_reset; // @[:@131040.4 RegFile.scala 76:16:@131047.4]
  assign regs_432_io_in = 64'h0; // @[RegFile.scala 75:16:@131046.4]
  assign regs_432_io_reset = reset; // @[RegFile.scala 78:19:@131050.4]
  assign regs_432_io_enable = 1'h1; // @[RegFile.scala 74:20:@131044.4]
  assign regs_433_clock = clock; // @[:@131053.4]
  assign regs_433_reset = io_reset; // @[:@131054.4 RegFile.scala 76:16:@131061.4]
  assign regs_433_io_in = 64'h0; // @[RegFile.scala 75:16:@131060.4]
  assign regs_433_io_reset = reset; // @[RegFile.scala 78:19:@131064.4]
  assign regs_433_io_enable = 1'h1; // @[RegFile.scala 74:20:@131058.4]
  assign regs_434_clock = clock; // @[:@131067.4]
  assign regs_434_reset = io_reset; // @[:@131068.4 RegFile.scala 76:16:@131075.4]
  assign regs_434_io_in = 64'h0; // @[RegFile.scala 75:16:@131074.4]
  assign regs_434_io_reset = reset; // @[RegFile.scala 78:19:@131078.4]
  assign regs_434_io_enable = 1'h1; // @[RegFile.scala 74:20:@131072.4]
  assign regs_435_clock = clock; // @[:@131081.4]
  assign regs_435_reset = io_reset; // @[:@131082.4 RegFile.scala 76:16:@131089.4]
  assign regs_435_io_in = 64'h0; // @[RegFile.scala 75:16:@131088.4]
  assign regs_435_io_reset = reset; // @[RegFile.scala 78:19:@131092.4]
  assign regs_435_io_enable = 1'h1; // @[RegFile.scala 74:20:@131086.4]
  assign regs_436_clock = clock; // @[:@131095.4]
  assign regs_436_reset = io_reset; // @[:@131096.4 RegFile.scala 76:16:@131103.4]
  assign regs_436_io_in = 64'h0; // @[RegFile.scala 75:16:@131102.4]
  assign regs_436_io_reset = reset; // @[RegFile.scala 78:19:@131106.4]
  assign regs_436_io_enable = 1'h1; // @[RegFile.scala 74:20:@131100.4]
  assign regs_437_clock = clock; // @[:@131109.4]
  assign regs_437_reset = io_reset; // @[:@131110.4 RegFile.scala 76:16:@131117.4]
  assign regs_437_io_in = 64'h0; // @[RegFile.scala 75:16:@131116.4]
  assign regs_437_io_reset = reset; // @[RegFile.scala 78:19:@131120.4]
  assign regs_437_io_enable = 1'h1; // @[RegFile.scala 74:20:@131114.4]
  assign regs_438_clock = clock; // @[:@131123.4]
  assign regs_438_reset = io_reset; // @[:@131124.4 RegFile.scala 76:16:@131131.4]
  assign regs_438_io_in = 64'h0; // @[RegFile.scala 75:16:@131130.4]
  assign regs_438_io_reset = reset; // @[RegFile.scala 78:19:@131134.4]
  assign regs_438_io_enable = 1'h1; // @[RegFile.scala 74:20:@131128.4]
  assign regs_439_clock = clock; // @[:@131137.4]
  assign regs_439_reset = io_reset; // @[:@131138.4 RegFile.scala 76:16:@131145.4]
  assign regs_439_io_in = 64'h0; // @[RegFile.scala 75:16:@131144.4]
  assign regs_439_io_reset = reset; // @[RegFile.scala 78:19:@131148.4]
  assign regs_439_io_enable = 1'h1; // @[RegFile.scala 74:20:@131142.4]
  assign regs_440_clock = clock; // @[:@131151.4]
  assign regs_440_reset = io_reset; // @[:@131152.4 RegFile.scala 76:16:@131159.4]
  assign regs_440_io_in = 64'h0; // @[RegFile.scala 75:16:@131158.4]
  assign regs_440_io_reset = reset; // @[RegFile.scala 78:19:@131162.4]
  assign regs_440_io_enable = 1'h1; // @[RegFile.scala 74:20:@131156.4]
  assign regs_441_clock = clock; // @[:@131165.4]
  assign regs_441_reset = io_reset; // @[:@131166.4 RegFile.scala 76:16:@131173.4]
  assign regs_441_io_in = 64'h0; // @[RegFile.scala 75:16:@131172.4]
  assign regs_441_io_reset = reset; // @[RegFile.scala 78:19:@131176.4]
  assign regs_441_io_enable = 1'h1; // @[RegFile.scala 74:20:@131170.4]
  assign regs_442_clock = clock; // @[:@131179.4]
  assign regs_442_reset = io_reset; // @[:@131180.4 RegFile.scala 76:16:@131187.4]
  assign regs_442_io_in = 64'h0; // @[RegFile.scala 75:16:@131186.4]
  assign regs_442_io_reset = reset; // @[RegFile.scala 78:19:@131190.4]
  assign regs_442_io_enable = 1'h1; // @[RegFile.scala 74:20:@131184.4]
  assign regs_443_clock = clock; // @[:@131193.4]
  assign regs_443_reset = io_reset; // @[:@131194.4 RegFile.scala 76:16:@131201.4]
  assign regs_443_io_in = 64'h0; // @[RegFile.scala 75:16:@131200.4]
  assign regs_443_io_reset = reset; // @[RegFile.scala 78:19:@131204.4]
  assign regs_443_io_enable = 1'h1; // @[RegFile.scala 74:20:@131198.4]
  assign regs_444_clock = clock; // @[:@131207.4]
  assign regs_444_reset = io_reset; // @[:@131208.4 RegFile.scala 76:16:@131215.4]
  assign regs_444_io_in = 64'h0; // @[RegFile.scala 75:16:@131214.4]
  assign regs_444_io_reset = reset; // @[RegFile.scala 78:19:@131218.4]
  assign regs_444_io_enable = 1'h1; // @[RegFile.scala 74:20:@131212.4]
  assign regs_445_clock = clock; // @[:@131221.4]
  assign regs_445_reset = io_reset; // @[:@131222.4 RegFile.scala 76:16:@131229.4]
  assign regs_445_io_in = 64'h0; // @[RegFile.scala 75:16:@131228.4]
  assign regs_445_io_reset = reset; // @[RegFile.scala 78:19:@131232.4]
  assign regs_445_io_enable = 1'h1; // @[RegFile.scala 74:20:@131226.4]
  assign regs_446_clock = clock; // @[:@131235.4]
  assign regs_446_reset = io_reset; // @[:@131236.4 RegFile.scala 76:16:@131243.4]
  assign regs_446_io_in = 64'h0; // @[RegFile.scala 75:16:@131242.4]
  assign regs_446_io_reset = reset; // @[RegFile.scala 78:19:@131246.4]
  assign regs_446_io_enable = 1'h1; // @[RegFile.scala 74:20:@131240.4]
  assign regs_447_clock = clock; // @[:@131249.4]
  assign regs_447_reset = io_reset; // @[:@131250.4 RegFile.scala 76:16:@131257.4]
  assign regs_447_io_in = 64'h0; // @[RegFile.scala 75:16:@131256.4]
  assign regs_447_io_reset = reset; // @[RegFile.scala 78:19:@131260.4]
  assign regs_447_io_enable = 1'h1; // @[RegFile.scala 74:20:@131254.4]
  assign regs_448_clock = clock; // @[:@131263.4]
  assign regs_448_reset = io_reset; // @[:@131264.4 RegFile.scala 76:16:@131271.4]
  assign regs_448_io_in = 64'h0; // @[RegFile.scala 75:16:@131270.4]
  assign regs_448_io_reset = reset; // @[RegFile.scala 78:19:@131274.4]
  assign regs_448_io_enable = 1'h1; // @[RegFile.scala 74:20:@131268.4]
  assign regs_449_clock = clock; // @[:@131277.4]
  assign regs_449_reset = io_reset; // @[:@131278.4 RegFile.scala 76:16:@131285.4]
  assign regs_449_io_in = 64'h0; // @[RegFile.scala 75:16:@131284.4]
  assign regs_449_io_reset = reset; // @[RegFile.scala 78:19:@131288.4]
  assign regs_449_io_enable = 1'h1; // @[RegFile.scala 74:20:@131282.4]
  assign regs_450_clock = clock; // @[:@131291.4]
  assign regs_450_reset = io_reset; // @[:@131292.4 RegFile.scala 76:16:@131299.4]
  assign regs_450_io_in = 64'h0; // @[RegFile.scala 75:16:@131298.4]
  assign regs_450_io_reset = reset; // @[RegFile.scala 78:19:@131302.4]
  assign regs_450_io_enable = 1'h1; // @[RegFile.scala 74:20:@131296.4]
  assign regs_451_clock = clock; // @[:@131305.4]
  assign regs_451_reset = io_reset; // @[:@131306.4 RegFile.scala 76:16:@131313.4]
  assign regs_451_io_in = 64'h0; // @[RegFile.scala 75:16:@131312.4]
  assign regs_451_io_reset = reset; // @[RegFile.scala 78:19:@131316.4]
  assign regs_451_io_enable = 1'h1; // @[RegFile.scala 74:20:@131310.4]
  assign regs_452_clock = clock; // @[:@131319.4]
  assign regs_452_reset = io_reset; // @[:@131320.4 RegFile.scala 76:16:@131327.4]
  assign regs_452_io_in = 64'h0; // @[RegFile.scala 75:16:@131326.4]
  assign regs_452_io_reset = reset; // @[RegFile.scala 78:19:@131330.4]
  assign regs_452_io_enable = 1'h1; // @[RegFile.scala 74:20:@131324.4]
  assign regs_453_clock = clock; // @[:@131333.4]
  assign regs_453_reset = io_reset; // @[:@131334.4 RegFile.scala 76:16:@131341.4]
  assign regs_453_io_in = 64'h0; // @[RegFile.scala 75:16:@131340.4]
  assign regs_453_io_reset = reset; // @[RegFile.scala 78:19:@131344.4]
  assign regs_453_io_enable = 1'h1; // @[RegFile.scala 74:20:@131338.4]
  assign regs_454_clock = clock; // @[:@131347.4]
  assign regs_454_reset = io_reset; // @[:@131348.4 RegFile.scala 76:16:@131355.4]
  assign regs_454_io_in = 64'h0; // @[RegFile.scala 75:16:@131354.4]
  assign regs_454_io_reset = reset; // @[RegFile.scala 78:19:@131358.4]
  assign regs_454_io_enable = 1'h1; // @[RegFile.scala 74:20:@131352.4]
  assign regs_455_clock = clock; // @[:@131361.4]
  assign regs_455_reset = io_reset; // @[:@131362.4 RegFile.scala 76:16:@131369.4]
  assign regs_455_io_in = 64'h0; // @[RegFile.scala 75:16:@131368.4]
  assign regs_455_io_reset = reset; // @[RegFile.scala 78:19:@131372.4]
  assign regs_455_io_enable = 1'h1; // @[RegFile.scala 74:20:@131366.4]
  assign regs_456_clock = clock; // @[:@131375.4]
  assign regs_456_reset = io_reset; // @[:@131376.4 RegFile.scala 76:16:@131383.4]
  assign regs_456_io_in = 64'h0; // @[RegFile.scala 75:16:@131382.4]
  assign regs_456_io_reset = reset; // @[RegFile.scala 78:19:@131386.4]
  assign regs_456_io_enable = 1'h1; // @[RegFile.scala 74:20:@131380.4]
  assign regs_457_clock = clock; // @[:@131389.4]
  assign regs_457_reset = io_reset; // @[:@131390.4 RegFile.scala 76:16:@131397.4]
  assign regs_457_io_in = 64'h0; // @[RegFile.scala 75:16:@131396.4]
  assign regs_457_io_reset = reset; // @[RegFile.scala 78:19:@131400.4]
  assign regs_457_io_enable = 1'h1; // @[RegFile.scala 74:20:@131394.4]
  assign regs_458_clock = clock; // @[:@131403.4]
  assign regs_458_reset = io_reset; // @[:@131404.4 RegFile.scala 76:16:@131411.4]
  assign regs_458_io_in = 64'h0; // @[RegFile.scala 75:16:@131410.4]
  assign regs_458_io_reset = reset; // @[RegFile.scala 78:19:@131414.4]
  assign regs_458_io_enable = 1'h1; // @[RegFile.scala 74:20:@131408.4]
  assign regs_459_clock = clock; // @[:@131417.4]
  assign regs_459_reset = io_reset; // @[:@131418.4 RegFile.scala 76:16:@131425.4]
  assign regs_459_io_in = 64'h0; // @[RegFile.scala 75:16:@131424.4]
  assign regs_459_io_reset = reset; // @[RegFile.scala 78:19:@131428.4]
  assign regs_459_io_enable = 1'h1; // @[RegFile.scala 74:20:@131422.4]
  assign regs_460_clock = clock; // @[:@131431.4]
  assign regs_460_reset = io_reset; // @[:@131432.4 RegFile.scala 76:16:@131439.4]
  assign regs_460_io_in = 64'h0; // @[RegFile.scala 75:16:@131438.4]
  assign regs_460_io_reset = reset; // @[RegFile.scala 78:19:@131442.4]
  assign regs_460_io_enable = 1'h1; // @[RegFile.scala 74:20:@131436.4]
  assign regs_461_clock = clock; // @[:@131445.4]
  assign regs_461_reset = io_reset; // @[:@131446.4 RegFile.scala 76:16:@131453.4]
  assign regs_461_io_in = 64'h0; // @[RegFile.scala 75:16:@131452.4]
  assign regs_461_io_reset = reset; // @[RegFile.scala 78:19:@131456.4]
  assign regs_461_io_enable = 1'h1; // @[RegFile.scala 74:20:@131450.4]
  assign regs_462_clock = clock; // @[:@131459.4]
  assign regs_462_reset = io_reset; // @[:@131460.4 RegFile.scala 76:16:@131467.4]
  assign regs_462_io_in = 64'h0; // @[RegFile.scala 75:16:@131466.4]
  assign regs_462_io_reset = reset; // @[RegFile.scala 78:19:@131470.4]
  assign regs_462_io_enable = 1'h1; // @[RegFile.scala 74:20:@131464.4]
  assign regs_463_clock = clock; // @[:@131473.4]
  assign regs_463_reset = io_reset; // @[:@131474.4 RegFile.scala 76:16:@131481.4]
  assign regs_463_io_in = 64'h0; // @[RegFile.scala 75:16:@131480.4]
  assign regs_463_io_reset = reset; // @[RegFile.scala 78:19:@131484.4]
  assign regs_463_io_enable = 1'h1; // @[RegFile.scala 74:20:@131478.4]
  assign regs_464_clock = clock; // @[:@131487.4]
  assign regs_464_reset = io_reset; // @[:@131488.4 RegFile.scala 76:16:@131495.4]
  assign regs_464_io_in = 64'h0; // @[RegFile.scala 75:16:@131494.4]
  assign regs_464_io_reset = reset; // @[RegFile.scala 78:19:@131498.4]
  assign regs_464_io_enable = 1'h1; // @[RegFile.scala 74:20:@131492.4]
  assign regs_465_clock = clock; // @[:@131501.4]
  assign regs_465_reset = io_reset; // @[:@131502.4 RegFile.scala 76:16:@131509.4]
  assign regs_465_io_in = 64'h0; // @[RegFile.scala 75:16:@131508.4]
  assign regs_465_io_reset = reset; // @[RegFile.scala 78:19:@131512.4]
  assign regs_465_io_enable = 1'h1; // @[RegFile.scala 74:20:@131506.4]
  assign regs_466_clock = clock; // @[:@131515.4]
  assign regs_466_reset = io_reset; // @[:@131516.4 RegFile.scala 76:16:@131523.4]
  assign regs_466_io_in = 64'h0; // @[RegFile.scala 75:16:@131522.4]
  assign regs_466_io_reset = reset; // @[RegFile.scala 78:19:@131526.4]
  assign regs_466_io_enable = 1'h1; // @[RegFile.scala 74:20:@131520.4]
  assign regs_467_clock = clock; // @[:@131529.4]
  assign regs_467_reset = io_reset; // @[:@131530.4 RegFile.scala 76:16:@131537.4]
  assign regs_467_io_in = 64'h0; // @[RegFile.scala 75:16:@131536.4]
  assign regs_467_io_reset = reset; // @[RegFile.scala 78:19:@131540.4]
  assign regs_467_io_enable = 1'h1; // @[RegFile.scala 74:20:@131534.4]
  assign regs_468_clock = clock; // @[:@131543.4]
  assign regs_468_reset = io_reset; // @[:@131544.4 RegFile.scala 76:16:@131551.4]
  assign regs_468_io_in = 64'h0; // @[RegFile.scala 75:16:@131550.4]
  assign regs_468_io_reset = reset; // @[RegFile.scala 78:19:@131554.4]
  assign regs_468_io_enable = 1'h1; // @[RegFile.scala 74:20:@131548.4]
  assign regs_469_clock = clock; // @[:@131557.4]
  assign regs_469_reset = io_reset; // @[:@131558.4 RegFile.scala 76:16:@131565.4]
  assign regs_469_io_in = 64'h0; // @[RegFile.scala 75:16:@131564.4]
  assign regs_469_io_reset = reset; // @[RegFile.scala 78:19:@131568.4]
  assign regs_469_io_enable = 1'h1; // @[RegFile.scala 74:20:@131562.4]
  assign regs_470_clock = clock; // @[:@131571.4]
  assign regs_470_reset = io_reset; // @[:@131572.4 RegFile.scala 76:16:@131579.4]
  assign regs_470_io_in = 64'h0; // @[RegFile.scala 75:16:@131578.4]
  assign regs_470_io_reset = reset; // @[RegFile.scala 78:19:@131582.4]
  assign regs_470_io_enable = 1'h1; // @[RegFile.scala 74:20:@131576.4]
  assign regs_471_clock = clock; // @[:@131585.4]
  assign regs_471_reset = io_reset; // @[:@131586.4 RegFile.scala 76:16:@131593.4]
  assign regs_471_io_in = 64'h0; // @[RegFile.scala 75:16:@131592.4]
  assign regs_471_io_reset = reset; // @[RegFile.scala 78:19:@131596.4]
  assign regs_471_io_enable = 1'h1; // @[RegFile.scala 74:20:@131590.4]
  assign regs_472_clock = clock; // @[:@131599.4]
  assign regs_472_reset = io_reset; // @[:@131600.4 RegFile.scala 76:16:@131607.4]
  assign regs_472_io_in = 64'h0; // @[RegFile.scala 75:16:@131606.4]
  assign regs_472_io_reset = reset; // @[RegFile.scala 78:19:@131610.4]
  assign regs_472_io_enable = 1'h1; // @[RegFile.scala 74:20:@131604.4]
  assign regs_473_clock = clock; // @[:@131613.4]
  assign regs_473_reset = io_reset; // @[:@131614.4 RegFile.scala 76:16:@131621.4]
  assign regs_473_io_in = 64'h0; // @[RegFile.scala 75:16:@131620.4]
  assign regs_473_io_reset = reset; // @[RegFile.scala 78:19:@131624.4]
  assign regs_473_io_enable = 1'h1; // @[RegFile.scala 74:20:@131618.4]
  assign regs_474_clock = clock; // @[:@131627.4]
  assign regs_474_reset = io_reset; // @[:@131628.4 RegFile.scala 76:16:@131635.4]
  assign regs_474_io_in = 64'h0; // @[RegFile.scala 75:16:@131634.4]
  assign regs_474_io_reset = reset; // @[RegFile.scala 78:19:@131638.4]
  assign regs_474_io_enable = 1'h1; // @[RegFile.scala 74:20:@131632.4]
  assign regs_475_clock = clock; // @[:@131641.4]
  assign regs_475_reset = io_reset; // @[:@131642.4 RegFile.scala 76:16:@131649.4]
  assign regs_475_io_in = 64'h0; // @[RegFile.scala 75:16:@131648.4]
  assign regs_475_io_reset = reset; // @[RegFile.scala 78:19:@131652.4]
  assign regs_475_io_enable = 1'h1; // @[RegFile.scala 74:20:@131646.4]
  assign regs_476_clock = clock; // @[:@131655.4]
  assign regs_476_reset = io_reset; // @[:@131656.4 RegFile.scala 76:16:@131663.4]
  assign regs_476_io_in = 64'h0; // @[RegFile.scala 75:16:@131662.4]
  assign regs_476_io_reset = reset; // @[RegFile.scala 78:19:@131666.4]
  assign regs_476_io_enable = 1'h1; // @[RegFile.scala 74:20:@131660.4]
  assign regs_477_clock = clock; // @[:@131669.4]
  assign regs_477_reset = io_reset; // @[:@131670.4 RegFile.scala 76:16:@131677.4]
  assign regs_477_io_in = 64'h0; // @[RegFile.scala 75:16:@131676.4]
  assign regs_477_io_reset = reset; // @[RegFile.scala 78:19:@131680.4]
  assign regs_477_io_enable = 1'h1; // @[RegFile.scala 74:20:@131674.4]
  assign regs_478_clock = clock; // @[:@131683.4]
  assign regs_478_reset = io_reset; // @[:@131684.4 RegFile.scala 76:16:@131691.4]
  assign regs_478_io_in = 64'h0; // @[RegFile.scala 75:16:@131690.4]
  assign regs_478_io_reset = reset; // @[RegFile.scala 78:19:@131694.4]
  assign regs_478_io_enable = 1'h1; // @[RegFile.scala 74:20:@131688.4]
  assign regs_479_clock = clock; // @[:@131697.4]
  assign regs_479_reset = io_reset; // @[:@131698.4 RegFile.scala 76:16:@131705.4]
  assign regs_479_io_in = 64'h0; // @[RegFile.scala 75:16:@131704.4]
  assign regs_479_io_reset = reset; // @[RegFile.scala 78:19:@131708.4]
  assign regs_479_io_enable = 1'h1; // @[RegFile.scala 74:20:@131702.4]
  assign regs_480_clock = clock; // @[:@131711.4]
  assign regs_480_reset = io_reset; // @[:@131712.4 RegFile.scala 76:16:@131719.4]
  assign regs_480_io_in = 64'h0; // @[RegFile.scala 75:16:@131718.4]
  assign regs_480_io_reset = reset; // @[RegFile.scala 78:19:@131722.4]
  assign regs_480_io_enable = 1'h1; // @[RegFile.scala 74:20:@131716.4]
  assign regs_481_clock = clock; // @[:@131725.4]
  assign regs_481_reset = io_reset; // @[:@131726.4 RegFile.scala 76:16:@131733.4]
  assign regs_481_io_in = 64'h0; // @[RegFile.scala 75:16:@131732.4]
  assign regs_481_io_reset = reset; // @[RegFile.scala 78:19:@131736.4]
  assign regs_481_io_enable = 1'h1; // @[RegFile.scala 74:20:@131730.4]
  assign regs_482_clock = clock; // @[:@131739.4]
  assign regs_482_reset = io_reset; // @[:@131740.4 RegFile.scala 76:16:@131747.4]
  assign regs_482_io_in = 64'h0; // @[RegFile.scala 75:16:@131746.4]
  assign regs_482_io_reset = reset; // @[RegFile.scala 78:19:@131750.4]
  assign regs_482_io_enable = 1'h1; // @[RegFile.scala 74:20:@131744.4]
  assign regs_483_clock = clock; // @[:@131753.4]
  assign regs_483_reset = io_reset; // @[:@131754.4 RegFile.scala 76:16:@131761.4]
  assign regs_483_io_in = 64'h0; // @[RegFile.scala 75:16:@131760.4]
  assign regs_483_io_reset = reset; // @[RegFile.scala 78:19:@131764.4]
  assign regs_483_io_enable = 1'h1; // @[RegFile.scala 74:20:@131758.4]
  assign regs_484_clock = clock; // @[:@131767.4]
  assign regs_484_reset = io_reset; // @[:@131768.4 RegFile.scala 76:16:@131775.4]
  assign regs_484_io_in = 64'h0; // @[RegFile.scala 75:16:@131774.4]
  assign regs_484_io_reset = reset; // @[RegFile.scala 78:19:@131778.4]
  assign regs_484_io_enable = 1'h1; // @[RegFile.scala 74:20:@131772.4]
  assign regs_485_clock = clock; // @[:@131781.4]
  assign regs_485_reset = io_reset; // @[:@131782.4 RegFile.scala 76:16:@131789.4]
  assign regs_485_io_in = 64'h0; // @[RegFile.scala 75:16:@131788.4]
  assign regs_485_io_reset = reset; // @[RegFile.scala 78:19:@131792.4]
  assign regs_485_io_enable = 1'h1; // @[RegFile.scala 74:20:@131786.4]
  assign regs_486_clock = clock; // @[:@131795.4]
  assign regs_486_reset = io_reset; // @[:@131796.4 RegFile.scala 76:16:@131803.4]
  assign regs_486_io_in = 64'h0; // @[RegFile.scala 75:16:@131802.4]
  assign regs_486_io_reset = reset; // @[RegFile.scala 78:19:@131806.4]
  assign regs_486_io_enable = 1'h1; // @[RegFile.scala 74:20:@131800.4]
  assign regs_487_clock = clock; // @[:@131809.4]
  assign regs_487_reset = io_reset; // @[:@131810.4 RegFile.scala 76:16:@131817.4]
  assign regs_487_io_in = 64'h0; // @[RegFile.scala 75:16:@131816.4]
  assign regs_487_io_reset = reset; // @[RegFile.scala 78:19:@131820.4]
  assign regs_487_io_enable = 1'h1; // @[RegFile.scala 74:20:@131814.4]
  assign regs_488_clock = clock; // @[:@131823.4]
  assign regs_488_reset = io_reset; // @[:@131824.4 RegFile.scala 76:16:@131831.4]
  assign regs_488_io_in = 64'h0; // @[RegFile.scala 75:16:@131830.4]
  assign regs_488_io_reset = reset; // @[RegFile.scala 78:19:@131834.4]
  assign regs_488_io_enable = 1'h1; // @[RegFile.scala 74:20:@131828.4]
  assign regs_489_clock = clock; // @[:@131837.4]
  assign regs_489_reset = io_reset; // @[:@131838.4 RegFile.scala 76:16:@131845.4]
  assign regs_489_io_in = 64'h0; // @[RegFile.scala 75:16:@131844.4]
  assign regs_489_io_reset = reset; // @[RegFile.scala 78:19:@131848.4]
  assign regs_489_io_enable = 1'h1; // @[RegFile.scala 74:20:@131842.4]
  assign regs_490_clock = clock; // @[:@131851.4]
  assign regs_490_reset = io_reset; // @[:@131852.4 RegFile.scala 76:16:@131859.4]
  assign regs_490_io_in = 64'h0; // @[RegFile.scala 75:16:@131858.4]
  assign regs_490_io_reset = reset; // @[RegFile.scala 78:19:@131862.4]
  assign regs_490_io_enable = 1'h1; // @[RegFile.scala 74:20:@131856.4]
  assign regs_491_clock = clock; // @[:@131865.4]
  assign regs_491_reset = io_reset; // @[:@131866.4 RegFile.scala 76:16:@131873.4]
  assign regs_491_io_in = 64'h0; // @[RegFile.scala 75:16:@131872.4]
  assign regs_491_io_reset = reset; // @[RegFile.scala 78:19:@131876.4]
  assign regs_491_io_enable = 1'h1; // @[RegFile.scala 74:20:@131870.4]
  assign regs_492_clock = clock; // @[:@131879.4]
  assign regs_492_reset = io_reset; // @[:@131880.4 RegFile.scala 76:16:@131887.4]
  assign regs_492_io_in = 64'h0; // @[RegFile.scala 75:16:@131886.4]
  assign regs_492_io_reset = reset; // @[RegFile.scala 78:19:@131890.4]
  assign regs_492_io_enable = 1'h1; // @[RegFile.scala 74:20:@131884.4]
  assign regs_493_clock = clock; // @[:@131893.4]
  assign regs_493_reset = io_reset; // @[:@131894.4 RegFile.scala 76:16:@131901.4]
  assign regs_493_io_in = 64'h0; // @[RegFile.scala 75:16:@131900.4]
  assign regs_493_io_reset = reset; // @[RegFile.scala 78:19:@131904.4]
  assign regs_493_io_enable = 1'h1; // @[RegFile.scala 74:20:@131898.4]
  assign regs_494_clock = clock; // @[:@131907.4]
  assign regs_494_reset = io_reset; // @[:@131908.4 RegFile.scala 76:16:@131915.4]
  assign regs_494_io_in = 64'h0; // @[RegFile.scala 75:16:@131914.4]
  assign regs_494_io_reset = reset; // @[RegFile.scala 78:19:@131918.4]
  assign regs_494_io_enable = 1'h1; // @[RegFile.scala 74:20:@131912.4]
  assign regs_495_clock = clock; // @[:@131921.4]
  assign regs_495_reset = io_reset; // @[:@131922.4 RegFile.scala 76:16:@131929.4]
  assign regs_495_io_in = 64'h0; // @[RegFile.scala 75:16:@131928.4]
  assign regs_495_io_reset = reset; // @[RegFile.scala 78:19:@131932.4]
  assign regs_495_io_enable = 1'h1; // @[RegFile.scala 74:20:@131926.4]
  assign regs_496_clock = clock; // @[:@131935.4]
  assign regs_496_reset = io_reset; // @[:@131936.4 RegFile.scala 76:16:@131943.4]
  assign regs_496_io_in = 64'h0; // @[RegFile.scala 75:16:@131942.4]
  assign regs_496_io_reset = reset; // @[RegFile.scala 78:19:@131946.4]
  assign regs_496_io_enable = 1'h1; // @[RegFile.scala 74:20:@131940.4]
  assign regs_497_clock = clock; // @[:@131949.4]
  assign regs_497_reset = io_reset; // @[:@131950.4 RegFile.scala 76:16:@131957.4]
  assign regs_497_io_in = 64'h0; // @[RegFile.scala 75:16:@131956.4]
  assign regs_497_io_reset = reset; // @[RegFile.scala 78:19:@131960.4]
  assign regs_497_io_enable = 1'h1; // @[RegFile.scala 74:20:@131954.4]
  assign regs_498_clock = clock; // @[:@131963.4]
  assign regs_498_reset = io_reset; // @[:@131964.4 RegFile.scala 76:16:@131971.4]
  assign regs_498_io_in = 64'h0; // @[RegFile.scala 75:16:@131970.4]
  assign regs_498_io_reset = reset; // @[RegFile.scala 78:19:@131974.4]
  assign regs_498_io_enable = 1'h1; // @[RegFile.scala 74:20:@131968.4]
  assign regs_499_clock = clock; // @[:@131977.4]
  assign regs_499_reset = io_reset; // @[:@131978.4 RegFile.scala 76:16:@131985.4]
  assign regs_499_io_in = 64'h0; // @[RegFile.scala 75:16:@131984.4]
  assign regs_499_io_reset = reset; // @[RegFile.scala 78:19:@131988.4]
  assign regs_499_io_enable = 1'h1; // @[RegFile.scala 74:20:@131982.4]
  assign regs_500_clock = clock; // @[:@131991.4]
  assign regs_500_reset = io_reset; // @[:@131992.4 RegFile.scala 76:16:@131999.4]
  assign regs_500_io_in = 64'h0; // @[RegFile.scala 75:16:@131998.4]
  assign regs_500_io_reset = reset; // @[RegFile.scala 78:19:@132002.4]
  assign regs_500_io_enable = 1'h1; // @[RegFile.scala 74:20:@131996.4]
  assign regs_501_clock = clock; // @[:@132005.4]
  assign regs_501_reset = io_reset; // @[:@132006.4 RegFile.scala 76:16:@132013.4]
  assign regs_501_io_in = 64'h0; // @[RegFile.scala 75:16:@132012.4]
  assign regs_501_io_reset = reset; // @[RegFile.scala 78:19:@132016.4]
  assign regs_501_io_enable = 1'h1; // @[RegFile.scala 74:20:@132010.4]
  assign regs_502_clock = clock; // @[:@132019.4]
  assign regs_502_reset = io_reset; // @[:@132020.4 RegFile.scala 76:16:@132027.4]
  assign regs_502_io_in = 64'h0; // @[RegFile.scala 75:16:@132026.4]
  assign regs_502_io_reset = reset; // @[RegFile.scala 78:19:@132030.4]
  assign regs_502_io_enable = 1'h1; // @[RegFile.scala 74:20:@132024.4]
  assign rport_io_ins_0 = regs_0_io_out; // @[RegFile.scala 97:16:@132539.4]
  assign rport_io_ins_1 = regs_1_io_out; // @[RegFile.scala 97:16:@132540.4]
  assign rport_io_ins_2 = regs_2_io_out; // @[RegFile.scala 97:16:@132541.4]
  assign rport_io_ins_3 = regs_3_io_out; // @[RegFile.scala 97:16:@132542.4]
  assign rport_io_ins_4 = regs_4_io_out; // @[RegFile.scala 97:16:@132543.4]
  assign rport_io_ins_5 = regs_5_io_out; // @[RegFile.scala 97:16:@132544.4]
  assign rport_io_ins_6 = regs_6_io_out; // @[RegFile.scala 97:16:@132545.4]
  assign rport_io_ins_7 = regs_7_io_out; // @[RegFile.scala 97:16:@132546.4]
  assign rport_io_ins_8 = regs_8_io_out; // @[RegFile.scala 97:16:@132547.4]
  assign rport_io_ins_9 = regs_9_io_out; // @[RegFile.scala 97:16:@132548.4]
  assign rport_io_ins_10 = regs_10_io_out; // @[RegFile.scala 97:16:@132549.4]
  assign rport_io_ins_11 = regs_11_io_out; // @[RegFile.scala 97:16:@132550.4]
  assign rport_io_ins_12 = regs_12_io_out; // @[RegFile.scala 97:16:@132551.4]
  assign rport_io_ins_13 = regs_13_io_out; // @[RegFile.scala 97:16:@132552.4]
  assign rport_io_ins_14 = regs_14_io_out; // @[RegFile.scala 97:16:@132553.4]
  assign rport_io_ins_15 = regs_15_io_out; // @[RegFile.scala 97:16:@132554.4]
  assign rport_io_ins_16 = regs_16_io_out; // @[RegFile.scala 97:16:@132555.4]
  assign rport_io_ins_17 = regs_17_io_out; // @[RegFile.scala 97:16:@132556.4]
  assign rport_io_ins_18 = regs_18_io_out; // @[RegFile.scala 97:16:@132557.4]
  assign rport_io_ins_19 = regs_19_io_out; // @[RegFile.scala 97:16:@132558.4]
  assign rport_io_ins_20 = regs_20_io_out; // @[RegFile.scala 97:16:@132559.4]
  assign rport_io_ins_21 = regs_21_io_out; // @[RegFile.scala 97:16:@132560.4]
  assign rport_io_ins_22 = regs_22_io_out; // @[RegFile.scala 97:16:@132561.4]
  assign rport_io_ins_23 = regs_23_io_out; // @[RegFile.scala 97:16:@132562.4]
  assign rport_io_ins_24 = regs_24_io_out; // @[RegFile.scala 97:16:@132563.4]
  assign rport_io_ins_25 = regs_25_io_out; // @[RegFile.scala 97:16:@132564.4]
  assign rport_io_ins_26 = regs_26_io_out; // @[RegFile.scala 97:16:@132565.4]
  assign rport_io_ins_27 = regs_27_io_out; // @[RegFile.scala 97:16:@132566.4]
  assign rport_io_ins_28 = regs_28_io_out; // @[RegFile.scala 97:16:@132567.4]
  assign rport_io_ins_29 = regs_29_io_out; // @[RegFile.scala 97:16:@132568.4]
  assign rport_io_ins_30 = regs_30_io_out; // @[RegFile.scala 97:16:@132569.4]
  assign rport_io_ins_31 = regs_31_io_out; // @[RegFile.scala 97:16:@132570.4]
  assign rport_io_ins_32 = regs_32_io_out; // @[RegFile.scala 97:16:@132571.4]
  assign rport_io_ins_33 = regs_33_io_out; // @[RegFile.scala 97:16:@132572.4]
  assign rport_io_ins_34 = regs_34_io_out; // @[RegFile.scala 97:16:@132573.4]
  assign rport_io_ins_35 = regs_35_io_out; // @[RegFile.scala 97:16:@132574.4]
  assign rport_io_ins_36 = regs_36_io_out; // @[RegFile.scala 97:16:@132575.4]
  assign rport_io_ins_37 = regs_37_io_out; // @[RegFile.scala 97:16:@132576.4]
  assign rport_io_ins_38 = regs_38_io_out; // @[RegFile.scala 97:16:@132577.4]
  assign rport_io_ins_39 = regs_39_io_out; // @[RegFile.scala 97:16:@132578.4]
  assign rport_io_ins_40 = regs_40_io_out; // @[RegFile.scala 97:16:@132579.4]
  assign rport_io_ins_41 = regs_41_io_out; // @[RegFile.scala 97:16:@132580.4]
  assign rport_io_ins_42 = regs_42_io_out; // @[RegFile.scala 97:16:@132581.4]
  assign rport_io_ins_43 = regs_43_io_out; // @[RegFile.scala 97:16:@132582.4]
  assign rport_io_ins_44 = regs_44_io_out; // @[RegFile.scala 97:16:@132583.4]
  assign rport_io_ins_45 = regs_45_io_out; // @[RegFile.scala 97:16:@132584.4]
  assign rport_io_ins_46 = regs_46_io_out; // @[RegFile.scala 97:16:@132585.4]
  assign rport_io_ins_47 = regs_47_io_out; // @[RegFile.scala 97:16:@132586.4]
  assign rport_io_ins_48 = regs_48_io_out; // @[RegFile.scala 97:16:@132587.4]
  assign rport_io_ins_49 = regs_49_io_out; // @[RegFile.scala 97:16:@132588.4]
  assign rport_io_ins_50 = regs_50_io_out; // @[RegFile.scala 97:16:@132589.4]
  assign rport_io_ins_51 = regs_51_io_out; // @[RegFile.scala 97:16:@132590.4]
  assign rport_io_ins_52 = regs_52_io_out; // @[RegFile.scala 97:16:@132591.4]
  assign rport_io_ins_53 = regs_53_io_out; // @[RegFile.scala 97:16:@132592.4]
  assign rport_io_ins_54 = regs_54_io_out; // @[RegFile.scala 97:16:@132593.4]
  assign rport_io_ins_55 = regs_55_io_out; // @[RegFile.scala 97:16:@132594.4]
  assign rport_io_ins_56 = regs_56_io_out; // @[RegFile.scala 97:16:@132595.4]
  assign rport_io_ins_57 = regs_57_io_out; // @[RegFile.scala 97:16:@132596.4]
  assign rport_io_ins_58 = regs_58_io_out; // @[RegFile.scala 97:16:@132597.4]
  assign rport_io_ins_59 = regs_59_io_out; // @[RegFile.scala 97:16:@132598.4]
  assign rport_io_ins_60 = regs_60_io_out; // @[RegFile.scala 97:16:@132599.4]
  assign rport_io_ins_61 = regs_61_io_out; // @[RegFile.scala 97:16:@132600.4]
  assign rport_io_ins_62 = regs_62_io_out; // @[RegFile.scala 97:16:@132601.4]
  assign rport_io_ins_63 = regs_63_io_out; // @[RegFile.scala 97:16:@132602.4]
  assign rport_io_ins_64 = regs_64_io_out; // @[RegFile.scala 97:16:@132603.4]
  assign rport_io_ins_65 = regs_65_io_out; // @[RegFile.scala 97:16:@132604.4]
  assign rport_io_ins_66 = regs_66_io_out; // @[RegFile.scala 97:16:@132605.4]
  assign rport_io_ins_67 = regs_67_io_out; // @[RegFile.scala 97:16:@132606.4]
  assign rport_io_ins_68 = regs_68_io_out; // @[RegFile.scala 97:16:@132607.4]
  assign rport_io_ins_69 = regs_69_io_out; // @[RegFile.scala 97:16:@132608.4]
  assign rport_io_ins_70 = regs_70_io_out; // @[RegFile.scala 97:16:@132609.4]
  assign rport_io_ins_71 = regs_71_io_out; // @[RegFile.scala 97:16:@132610.4]
  assign rport_io_ins_72 = regs_72_io_out; // @[RegFile.scala 97:16:@132611.4]
  assign rport_io_ins_73 = regs_73_io_out; // @[RegFile.scala 97:16:@132612.4]
  assign rport_io_ins_74 = regs_74_io_out; // @[RegFile.scala 97:16:@132613.4]
  assign rport_io_ins_75 = regs_75_io_out; // @[RegFile.scala 97:16:@132614.4]
  assign rport_io_ins_76 = regs_76_io_out; // @[RegFile.scala 97:16:@132615.4]
  assign rport_io_ins_77 = regs_77_io_out; // @[RegFile.scala 97:16:@132616.4]
  assign rport_io_ins_78 = regs_78_io_out; // @[RegFile.scala 97:16:@132617.4]
  assign rport_io_ins_79 = regs_79_io_out; // @[RegFile.scala 97:16:@132618.4]
  assign rport_io_ins_80 = regs_80_io_out; // @[RegFile.scala 97:16:@132619.4]
  assign rport_io_ins_81 = regs_81_io_out; // @[RegFile.scala 97:16:@132620.4]
  assign rport_io_ins_82 = regs_82_io_out; // @[RegFile.scala 97:16:@132621.4]
  assign rport_io_ins_83 = regs_83_io_out; // @[RegFile.scala 97:16:@132622.4]
  assign rport_io_ins_84 = regs_84_io_out; // @[RegFile.scala 97:16:@132623.4]
  assign rport_io_ins_85 = regs_85_io_out; // @[RegFile.scala 97:16:@132624.4]
  assign rport_io_ins_86 = regs_86_io_out; // @[RegFile.scala 97:16:@132625.4]
  assign rport_io_ins_87 = regs_87_io_out; // @[RegFile.scala 97:16:@132626.4]
  assign rport_io_ins_88 = regs_88_io_out; // @[RegFile.scala 97:16:@132627.4]
  assign rport_io_ins_89 = regs_89_io_out; // @[RegFile.scala 97:16:@132628.4]
  assign rport_io_ins_90 = regs_90_io_out; // @[RegFile.scala 97:16:@132629.4]
  assign rport_io_ins_91 = regs_91_io_out; // @[RegFile.scala 97:16:@132630.4]
  assign rport_io_ins_92 = regs_92_io_out; // @[RegFile.scala 97:16:@132631.4]
  assign rport_io_ins_93 = regs_93_io_out; // @[RegFile.scala 97:16:@132632.4]
  assign rport_io_ins_94 = regs_94_io_out; // @[RegFile.scala 97:16:@132633.4]
  assign rport_io_ins_95 = regs_95_io_out; // @[RegFile.scala 97:16:@132634.4]
  assign rport_io_ins_96 = regs_96_io_out; // @[RegFile.scala 97:16:@132635.4]
  assign rport_io_ins_97 = regs_97_io_out; // @[RegFile.scala 97:16:@132636.4]
  assign rport_io_ins_98 = regs_98_io_out; // @[RegFile.scala 97:16:@132637.4]
  assign rport_io_ins_99 = regs_99_io_out; // @[RegFile.scala 97:16:@132638.4]
  assign rport_io_ins_100 = regs_100_io_out; // @[RegFile.scala 97:16:@132639.4]
  assign rport_io_ins_101 = regs_101_io_out; // @[RegFile.scala 97:16:@132640.4]
  assign rport_io_ins_102 = regs_102_io_out; // @[RegFile.scala 97:16:@132641.4]
  assign rport_io_ins_103 = regs_103_io_out; // @[RegFile.scala 97:16:@132642.4]
  assign rport_io_ins_104 = regs_104_io_out; // @[RegFile.scala 97:16:@132643.4]
  assign rport_io_ins_105 = regs_105_io_out; // @[RegFile.scala 97:16:@132644.4]
  assign rport_io_ins_106 = regs_106_io_out; // @[RegFile.scala 97:16:@132645.4]
  assign rport_io_ins_107 = regs_107_io_out; // @[RegFile.scala 97:16:@132646.4]
  assign rport_io_ins_108 = regs_108_io_out; // @[RegFile.scala 97:16:@132647.4]
  assign rport_io_ins_109 = regs_109_io_out; // @[RegFile.scala 97:16:@132648.4]
  assign rport_io_ins_110 = regs_110_io_out; // @[RegFile.scala 97:16:@132649.4]
  assign rport_io_ins_111 = regs_111_io_out; // @[RegFile.scala 97:16:@132650.4]
  assign rport_io_ins_112 = regs_112_io_out; // @[RegFile.scala 97:16:@132651.4]
  assign rport_io_ins_113 = regs_113_io_out; // @[RegFile.scala 97:16:@132652.4]
  assign rport_io_ins_114 = regs_114_io_out; // @[RegFile.scala 97:16:@132653.4]
  assign rport_io_ins_115 = regs_115_io_out; // @[RegFile.scala 97:16:@132654.4]
  assign rport_io_ins_116 = regs_116_io_out; // @[RegFile.scala 97:16:@132655.4]
  assign rport_io_ins_117 = regs_117_io_out; // @[RegFile.scala 97:16:@132656.4]
  assign rport_io_ins_118 = regs_118_io_out; // @[RegFile.scala 97:16:@132657.4]
  assign rport_io_ins_119 = regs_119_io_out; // @[RegFile.scala 97:16:@132658.4]
  assign rport_io_ins_120 = regs_120_io_out; // @[RegFile.scala 97:16:@132659.4]
  assign rport_io_ins_121 = regs_121_io_out; // @[RegFile.scala 97:16:@132660.4]
  assign rport_io_ins_122 = regs_122_io_out; // @[RegFile.scala 97:16:@132661.4]
  assign rport_io_ins_123 = regs_123_io_out; // @[RegFile.scala 97:16:@132662.4]
  assign rport_io_ins_124 = regs_124_io_out; // @[RegFile.scala 97:16:@132663.4]
  assign rport_io_ins_125 = regs_125_io_out; // @[RegFile.scala 97:16:@132664.4]
  assign rport_io_ins_126 = regs_126_io_out; // @[RegFile.scala 97:16:@132665.4]
  assign rport_io_ins_127 = regs_127_io_out; // @[RegFile.scala 97:16:@132666.4]
  assign rport_io_ins_128 = regs_128_io_out; // @[RegFile.scala 97:16:@132667.4]
  assign rport_io_ins_129 = regs_129_io_out; // @[RegFile.scala 97:16:@132668.4]
  assign rport_io_ins_130 = regs_130_io_out; // @[RegFile.scala 97:16:@132669.4]
  assign rport_io_ins_131 = regs_131_io_out; // @[RegFile.scala 97:16:@132670.4]
  assign rport_io_ins_132 = regs_132_io_out; // @[RegFile.scala 97:16:@132671.4]
  assign rport_io_ins_133 = regs_133_io_out; // @[RegFile.scala 97:16:@132672.4]
  assign rport_io_ins_134 = regs_134_io_out; // @[RegFile.scala 97:16:@132673.4]
  assign rport_io_ins_135 = regs_135_io_out; // @[RegFile.scala 97:16:@132674.4]
  assign rport_io_ins_136 = regs_136_io_out; // @[RegFile.scala 97:16:@132675.4]
  assign rport_io_ins_137 = regs_137_io_out; // @[RegFile.scala 97:16:@132676.4]
  assign rport_io_ins_138 = regs_138_io_out; // @[RegFile.scala 97:16:@132677.4]
  assign rport_io_ins_139 = regs_139_io_out; // @[RegFile.scala 97:16:@132678.4]
  assign rport_io_ins_140 = regs_140_io_out; // @[RegFile.scala 97:16:@132679.4]
  assign rport_io_ins_141 = regs_141_io_out; // @[RegFile.scala 97:16:@132680.4]
  assign rport_io_ins_142 = regs_142_io_out; // @[RegFile.scala 97:16:@132681.4]
  assign rport_io_ins_143 = regs_143_io_out; // @[RegFile.scala 97:16:@132682.4]
  assign rport_io_ins_144 = regs_144_io_out; // @[RegFile.scala 97:16:@132683.4]
  assign rport_io_ins_145 = regs_145_io_out; // @[RegFile.scala 97:16:@132684.4]
  assign rport_io_ins_146 = regs_146_io_out; // @[RegFile.scala 97:16:@132685.4]
  assign rport_io_ins_147 = regs_147_io_out; // @[RegFile.scala 97:16:@132686.4]
  assign rport_io_ins_148 = regs_148_io_out; // @[RegFile.scala 97:16:@132687.4]
  assign rport_io_ins_149 = regs_149_io_out; // @[RegFile.scala 97:16:@132688.4]
  assign rport_io_ins_150 = regs_150_io_out; // @[RegFile.scala 97:16:@132689.4]
  assign rport_io_ins_151 = regs_151_io_out; // @[RegFile.scala 97:16:@132690.4]
  assign rport_io_ins_152 = regs_152_io_out; // @[RegFile.scala 97:16:@132691.4]
  assign rport_io_ins_153 = regs_153_io_out; // @[RegFile.scala 97:16:@132692.4]
  assign rport_io_ins_154 = regs_154_io_out; // @[RegFile.scala 97:16:@132693.4]
  assign rport_io_ins_155 = regs_155_io_out; // @[RegFile.scala 97:16:@132694.4]
  assign rport_io_ins_156 = regs_156_io_out; // @[RegFile.scala 97:16:@132695.4]
  assign rport_io_ins_157 = regs_157_io_out; // @[RegFile.scala 97:16:@132696.4]
  assign rport_io_ins_158 = regs_158_io_out; // @[RegFile.scala 97:16:@132697.4]
  assign rport_io_ins_159 = regs_159_io_out; // @[RegFile.scala 97:16:@132698.4]
  assign rport_io_ins_160 = regs_160_io_out; // @[RegFile.scala 97:16:@132699.4]
  assign rport_io_ins_161 = regs_161_io_out; // @[RegFile.scala 97:16:@132700.4]
  assign rport_io_ins_162 = regs_162_io_out; // @[RegFile.scala 97:16:@132701.4]
  assign rport_io_ins_163 = regs_163_io_out; // @[RegFile.scala 97:16:@132702.4]
  assign rport_io_ins_164 = regs_164_io_out; // @[RegFile.scala 97:16:@132703.4]
  assign rport_io_ins_165 = regs_165_io_out; // @[RegFile.scala 97:16:@132704.4]
  assign rport_io_ins_166 = regs_166_io_out; // @[RegFile.scala 97:16:@132705.4]
  assign rport_io_ins_167 = regs_167_io_out; // @[RegFile.scala 97:16:@132706.4]
  assign rport_io_ins_168 = regs_168_io_out; // @[RegFile.scala 97:16:@132707.4]
  assign rport_io_ins_169 = regs_169_io_out; // @[RegFile.scala 97:16:@132708.4]
  assign rport_io_ins_170 = regs_170_io_out; // @[RegFile.scala 97:16:@132709.4]
  assign rport_io_ins_171 = regs_171_io_out; // @[RegFile.scala 97:16:@132710.4]
  assign rport_io_ins_172 = regs_172_io_out; // @[RegFile.scala 97:16:@132711.4]
  assign rport_io_ins_173 = regs_173_io_out; // @[RegFile.scala 97:16:@132712.4]
  assign rport_io_ins_174 = regs_174_io_out; // @[RegFile.scala 97:16:@132713.4]
  assign rport_io_ins_175 = regs_175_io_out; // @[RegFile.scala 97:16:@132714.4]
  assign rport_io_ins_176 = regs_176_io_out; // @[RegFile.scala 97:16:@132715.4]
  assign rport_io_ins_177 = regs_177_io_out; // @[RegFile.scala 97:16:@132716.4]
  assign rport_io_ins_178 = regs_178_io_out; // @[RegFile.scala 97:16:@132717.4]
  assign rport_io_ins_179 = regs_179_io_out; // @[RegFile.scala 97:16:@132718.4]
  assign rport_io_ins_180 = regs_180_io_out; // @[RegFile.scala 97:16:@132719.4]
  assign rport_io_ins_181 = regs_181_io_out; // @[RegFile.scala 97:16:@132720.4]
  assign rport_io_ins_182 = regs_182_io_out; // @[RegFile.scala 97:16:@132721.4]
  assign rport_io_ins_183 = regs_183_io_out; // @[RegFile.scala 97:16:@132722.4]
  assign rport_io_ins_184 = regs_184_io_out; // @[RegFile.scala 97:16:@132723.4]
  assign rport_io_ins_185 = regs_185_io_out; // @[RegFile.scala 97:16:@132724.4]
  assign rport_io_ins_186 = regs_186_io_out; // @[RegFile.scala 97:16:@132725.4]
  assign rport_io_ins_187 = regs_187_io_out; // @[RegFile.scala 97:16:@132726.4]
  assign rport_io_ins_188 = regs_188_io_out; // @[RegFile.scala 97:16:@132727.4]
  assign rport_io_ins_189 = regs_189_io_out; // @[RegFile.scala 97:16:@132728.4]
  assign rport_io_ins_190 = regs_190_io_out; // @[RegFile.scala 97:16:@132729.4]
  assign rport_io_ins_191 = regs_191_io_out; // @[RegFile.scala 97:16:@132730.4]
  assign rport_io_ins_192 = regs_192_io_out; // @[RegFile.scala 97:16:@132731.4]
  assign rport_io_ins_193 = regs_193_io_out; // @[RegFile.scala 97:16:@132732.4]
  assign rport_io_ins_194 = regs_194_io_out; // @[RegFile.scala 97:16:@132733.4]
  assign rport_io_ins_195 = regs_195_io_out; // @[RegFile.scala 97:16:@132734.4]
  assign rport_io_ins_196 = regs_196_io_out; // @[RegFile.scala 97:16:@132735.4]
  assign rport_io_ins_197 = regs_197_io_out; // @[RegFile.scala 97:16:@132736.4]
  assign rport_io_ins_198 = regs_198_io_out; // @[RegFile.scala 97:16:@132737.4]
  assign rport_io_ins_199 = regs_199_io_out; // @[RegFile.scala 97:16:@132738.4]
  assign rport_io_ins_200 = regs_200_io_out; // @[RegFile.scala 97:16:@132739.4]
  assign rport_io_ins_201 = regs_201_io_out; // @[RegFile.scala 97:16:@132740.4]
  assign rport_io_ins_202 = regs_202_io_out; // @[RegFile.scala 97:16:@132741.4]
  assign rport_io_ins_203 = regs_203_io_out; // @[RegFile.scala 97:16:@132742.4]
  assign rport_io_ins_204 = regs_204_io_out; // @[RegFile.scala 97:16:@132743.4]
  assign rport_io_ins_205 = regs_205_io_out; // @[RegFile.scala 97:16:@132744.4]
  assign rport_io_ins_206 = regs_206_io_out; // @[RegFile.scala 97:16:@132745.4]
  assign rport_io_ins_207 = regs_207_io_out; // @[RegFile.scala 97:16:@132746.4]
  assign rport_io_ins_208 = regs_208_io_out; // @[RegFile.scala 97:16:@132747.4]
  assign rport_io_ins_209 = regs_209_io_out; // @[RegFile.scala 97:16:@132748.4]
  assign rport_io_ins_210 = regs_210_io_out; // @[RegFile.scala 97:16:@132749.4]
  assign rport_io_ins_211 = regs_211_io_out; // @[RegFile.scala 97:16:@132750.4]
  assign rport_io_ins_212 = regs_212_io_out; // @[RegFile.scala 97:16:@132751.4]
  assign rport_io_ins_213 = regs_213_io_out; // @[RegFile.scala 97:16:@132752.4]
  assign rport_io_ins_214 = regs_214_io_out; // @[RegFile.scala 97:16:@132753.4]
  assign rport_io_ins_215 = regs_215_io_out; // @[RegFile.scala 97:16:@132754.4]
  assign rport_io_ins_216 = regs_216_io_out; // @[RegFile.scala 97:16:@132755.4]
  assign rport_io_ins_217 = regs_217_io_out; // @[RegFile.scala 97:16:@132756.4]
  assign rport_io_ins_218 = regs_218_io_out; // @[RegFile.scala 97:16:@132757.4]
  assign rport_io_ins_219 = regs_219_io_out; // @[RegFile.scala 97:16:@132758.4]
  assign rport_io_ins_220 = regs_220_io_out; // @[RegFile.scala 97:16:@132759.4]
  assign rport_io_ins_221 = regs_221_io_out; // @[RegFile.scala 97:16:@132760.4]
  assign rport_io_ins_222 = regs_222_io_out; // @[RegFile.scala 97:16:@132761.4]
  assign rport_io_ins_223 = regs_223_io_out; // @[RegFile.scala 97:16:@132762.4]
  assign rport_io_ins_224 = regs_224_io_out; // @[RegFile.scala 97:16:@132763.4]
  assign rport_io_ins_225 = regs_225_io_out; // @[RegFile.scala 97:16:@132764.4]
  assign rport_io_ins_226 = regs_226_io_out; // @[RegFile.scala 97:16:@132765.4]
  assign rport_io_ins_227 = regs_227_io_out; // @[RegFile.scala 97:16:@132766.4]
  assign rport_io_ins_228 = regs_228_io_out; // @[RegFile.scala 97:16:@132767.4]
  assign rport_io_ins_229 = regs_229_io_out; // @[RegFile.scala 97:16:@132768.4]
  assign rport_io_ins_230 = regs_230_io_out; // @[RegFile.scala 97:16:@132769.4]
  assign rport_io_ins_231 = regs_231_io_out; // @[RegFile.scala 97:16:@132770.4]
  assign rport_io_ins_232 = regs_232_io_out; // @[RegFile.scala 97:16:@132771.4]
  assign rport_io_ins_233 = regs_233_io_out; // @[RegFile.scala 97:16:@132772.4]
  assign rport_io_ins_234 = regs_234_io_out; // @[RegFile.scala 97:16:@132773.4]
  assign rport_io_ins_235 = regs_235_io_out; // @[RegFile.scala 97:16:@132774.4]
  assign rport_io_ins_236 = regs_236_io_out; // @[RegFile.scala 97:16:@132775.4]
  assign rport_io_ins_237 = regs_237_io_out; // @[RegFile.scala 97:16:@132776.4]
  assign rport_io_ins_238 = regs_238_io_out; // @[RegFile.scala 97:16:@132777.4]
  assign rport_io_ins_239 = regs_239_io_out; // @[RegFile.scala 97:16:@132778.4]
  assign rport_io_ins_240 = regs_240_io_out; // @[RegFile.scala 97:16:@132779.4]
  assign rport_io_ins_241 = regs_241_io_out; // @[RegFile.scala 97:16:@132780.4]
  assign rport_io_ins_242 = regs_242_io_out; // @[RegFile.scala 97:16:@132781.4]
  assign rport_io_ins_243 = regs_243_io_out; // @[RegFile.scala 97:16:@132782.4]
  assign rport_io_ins_244 = regs_244_io_out; // @[RegFile.scala 97:16:@132783.4]
  assign rport_io_ins_245 = regs_245_io_out; // @[RegFile.scala 97:16:@132784.4]
  assign rport_io_ins_246 = regs_246_io_out; // @[RegFile.scala 97:16:@132785.4]
  assign rport_io_ins_247 = regs_247_io_out; // @[RegFile.scala 97:16:@132786.4]
  assign rport_io_ins_248 = regs_248_io_out; // @[RegFile.scala 97:16:@132787.4]
  assign rport_io_ins_249 = regs_249_io_out; // @[RegFile.scala 97:16:@132788.4]
  assign rport_io_ins_250 = regs_250_io_out; // @[RegFile.scala 97:16:@132789.4]
  assign rport_io_ins_251 = regs_251_io_out; // @[RegFile.scala 97:16:@132790.4]
  assign rport_io_ins_252 = regs_252_io_out; // @[RegFile.scala 97:16:@132791.4]
  assign rport_io_ins_253 = regs_253_io_out; // @[RegFile.scala 97:16:@132792.4]
  assign rport_io_ins_254 = regs_254_io_out; // @[RegFile.scala 97:16:@132793.4]
  assign rport_io_ins_255 = regs_255_io_out; // @[RegFile.scala 97:16:@132794.4]
  assign rport_io_ins_256 = regs_256_io_out; // @[RegFile.scala 97:16:@132795.4]
  assign rport_io_ins_257 = regs_257_io_out; // @[RegFile.scala 97:16:@132796.4]
  assign rport_io_ins_258 = regs_258_io_out; // @[RegFile.scala 97:16:@132797.4]
  assign rport_io_ins_259 = regs_259_io_out; // @[RegFile.scala 97:16:@132798.4]
  assign rport_io_ins_260 = regs_260_io_out; // @[RegFile.scala 97:16:@132799.4]
  assign rport_io_ins_261 = regs_261_io_out; // @[RegFile.scala 97:16:@132800.4]
  assign rport_io_ins_262 = regs_262_io_out; // @[RegFile.scala 97:16:@132801.4]
  assign rport_io_ins_263 = regs_263_io_out; // @[RegFile.scala 97:16:@132802.4]
  assign rport_io_ins_264 = regs_264_io_out; // @[RegFile.scala 97:16:@132803.4]
  assign rport_io_ins_265 = regs_265_io_out; // @[RegFile.scala 97:16:@132804.4]
  assign rport_io_ins_266 = regs_266_io_out; // @[RegFile.scala 97:16:@132805.4]
  assign rport_io_ins_267 = regs_267_io_out; // @[RegFile.scala 97:16:@132806.4]
  assign rport_io_ins_268 = regs_268_io_out; // @[RegFile.scala 97:16:@132807.4]
  assign rport_io_ins_269 = regs_269_io_out; // @[RegFile.scala 97:16:@132808.4]
  assign rport_io_ins_270 = regs_270_io_out; // @[RegFile.scala 97:16:@132809.4]
  assign rport_io_ins_271 = regs_271_io_out; // @[RegFile.scala 97:16:@132810.4]
  assign rport_io_ins_272 = regs_272_io_out; // @[RegFile.scala 97:16:@132811.4]
  assign rport_io_ins_273 = regs_273_io_out; // @[RegFile.scala 97:16:@132812.4]
  assign rport_io_ins_274 = regs_274_io_out; // @[RegFile.scala 97:16:@132813.4]
  assign rport_io_ins_275 = regs_275_io_out; // @[RegFile.scala 97:16:@132814.4]
  assign rport_io_ins_276 = regs_276_io_out; // @[RegFile.scala 97:16:@132815.4]
  assign rport_io_ins_277 = regs_277_io_out; // @[RegFile.scala 97:16:@132816.4]
  assign rport_io_ins_278 = regs_278_io_out; // @[RegFile.scala 97:16:@132817.4]
  assign rport_io_ins_279 = regs_279_io_out; // @[RegFile.scala 97:16:@132818.4]
  assign rport_io_ins_280 = regs_280_io_out; // @[RegFile.scala 97:16:@132819.4]
  assign rport_io_ins_281 = regs_281_io_out; // @[RegFile.scala 97:16:@132820.4]
  assign rport_io_ins_282 = regs_282_io_out; // @[RegFile.scala 97:16:@132821.4]
  assign rport_io_ins_283 = regs_283_io_out; // @[RegFile.scala 97:16:@132822.4]
  assign rport_io_ins_284 = regs_284_io_out; // @[RegFile.scala 97:16:@132823.4]
  assign rport_io_ins_285 = regs_285_io_out; // @[RegFile.scala 97:16:@132824.4]
  assign rport_io_ins_286 = regs_286_io_out; // @[RegFile.scala 97:16:@132825.4]
  assign rport_io_ins_287 = regs_287_io_out; // @[RegFile.scala 97:16:@132826.4]
  assign rport_io_ins_288 = regs_288_io_out; // @[RegFile.scala 97:16:@132827.4]
  assign rport_io_ins_289 = regs_289_io_out; // @[RegFile.scala 97:16:@132828.4]
  assign rport_io_ins_290 = regs_290_io_out; // @[RegFile.scala 97:16:@132829.4]
  assign rport_io_ins_291 = regs_291_io_out; // @[RegFile.scala 97:16:@132830.4]
  assign rport_io_ins_292 = regs_292_io_out; // @[RegFile.scala 97:16:@132831.4]
  assign rport_io_ins_293 = regs_293_io_out; // @[RegFile.scala 97:16:@132832.4]
  assign rport_io_ins_294 = regs_294_io_out; // @[RegFile.scala 97:16:@132833.4]
  assign rport_io_ins_295 = regs_295_io_out; // @[RegFile.scala 97:16:@132834.4]
  assign rport_io_ins_296 = regs_296_io_out; // @[RegFile.scala 97:16:@132835.4]
  assign rport_io_ins_297 = regs_297_io_out; // @[RegFile.scala 97:16:@132836.4]
  assign rport_io_ins_298 = regs_298_io_out; // @[RegFile.scala 97:16:@132837.4]
  assign rport_io_ins_299 = regs_299_io_out; // @[RegFile.scala 97:16:@132838.4]
  assign rport_io_ins_300 = regs_300_io_out; // @[RegFile.scala 97:16:@132839.4]
  assign rport_io_ins_301 = regs_301_io_out; // @[RegFile.scala 97:16:@132840.4]
  assign rport_io_ins_302 = regs_302_io_out; // @[RegFile.scala 97:16:@132841.4]
  assign rport_io_ins_303 = regs_303_io_out; // @[RegFile.scala 97:16:@132842.4]
  assign rport_io_ins_304 = regs_304_io_out; // @[RegFile.scala 97:16:@132843.4]
  assign rport_io_ins_305 = regs_305_io_out; // @[RegFile.scala 97:16:@132844.4]
  assign rport_io_ins_306 = regs_306_io_out; // @[RegFile.scala 97:16:@132845.4]
  assign rport_io_ins_307 = regs_307_io_out; // @[RegFile.scala 97:16:@132846.4]
  assign rport_io_ins_308 = regs_308_io_out; // @[RegFile.scala 97:16:@132847.4]
  assign rport_io_ins_309 = regs_309_io_out; // @[RegFile.scala 97:16:@132848.4]
  assign rport_io_ins_310 = regs_310_io_out; // @[RegFile.scala 97:16:@132849.4]
  assign rport_io_ins_311 = regs_311_io_out; // @[RegFile.scala 97:16:@132850.4]
  assign rport_io_ins_312 = regs_312_io_out; // @[RegFile.scala 97:16:@132851.4]
  assign rport_io_ins_313 = regs_313_io_out; // @[RegFile.scala 97:16:@132852.4]
  assign rport_io_ins_314 = regs_314_io_out; // @[RegFile.scala 97:16:@132853.4]
  assign rport_io_ins_315 = regs_315_io_out; // @[RegFile.scala 97:16:@132854.4]
  assign rport_io_ins_316 = regs_316_io_out; // @[RegFile.scala 97:16:@132855.4]
  assign rport_io_ins_317 = regs_317_io_out; // @[RegFile.scala 97:16:@132856.4]
  assign rport_io_ins_318 = regs_318_io_out; // @[RegFile.scala 97:16:@132857.4]
  assign rport_io_ins_319 = regs_319_io_out; // @[RegFile.scala 97:16:@132858.4]
  assign rport_io_ins_320 = regs_320_io_out; // @[RegFile.scala 97:16:@132859.4]
  assign rport_io_ins_321 = regs_321_io_out; // @[RegFile.scala 97:16:@132860.4]
  assign rport_io_ins_322 = regs_322_io_out; // @[RegFile.scala 97:16:@132861.4]
  assign rport_io_ins_323 = regs_323_io_out; // @[RegFile.scala 97:16:@132862.4]
  assign rport_io_ins_324 = regs_324_io_out; // @[RegFile.scala 97:16:@132863.4]
  assign rport_io_ins_325 = regs_325_io_out; // @[RegFile.scala 97:16:@132864.4]
  assign rport_io_ins_326 = regs_326_io_out; // @[RegFile.scala 97:16:@132865.4]
  assign rport_io_ins_327 = regs_327_io_out; // @[RegFile.scala 97:16:@132866.4]
  assign rport_io_ins_328 = regs_328_io_out; // @[RegFile.scala 97:16:@132867.4]
  assign rport_io_ins_329 = regs_329_io_out; // @[RegFile.scala 97:16:@132868.4]
  assign rport_io_ins_330 = regs_330_io_out; // @[RegFile.scala 97:16:@132869.4]
  assign rport_io_ins_331 = regs_331_io_out; // @[RegFile.scala 97:16:@132870.4]
  assign rport_io_ins_332 = regs_332_io_out; // @[RegFile.scala 97:16:@132871.4]
  assign rport_io_ins_333 = regs_333_io_out; // @[RegFile.scala 97:16:@132872.4]
  assign rport_io_ins_334 = regs_334_io_out; // @[RegFile.scala 97:16:@132873.4]
  assign rport_io_ins_335 = regs_335_io_out; // @[RegFile.scala 97:16:@132874.4]
  assign rport_io_ins_336 = regs_336_io_out; // @[RegFile.scala 97:16:@132875.4]
  assign rport_io_ins_337 = regs_337_io_out; // @[RegFile.scala 97:16:@132876.4]
  assign rport_io_ins_338 = regs_338_io_out; // @[RegFile.scala 97:16:@132877.4]
  assign rport_io_ins_339 = regs_339_io_out; // @[RegFile.scala 97:16:@132878.4]
  assign rport_io_ins_340 = regs_340_io_out; // @[RegFile.scala 97:16:@132879.4]
  assign rport_io_ins_341 = regs_341_io_out; // @[RegFile.scala 97:16:@132880.4]
  assign rport_io_ins_342 = regs_342_io_out; // @[RegFile.scala 97:16:@132881.4]
  assign rport_io_ins_343 = regs_343_io_out; // @[RegFile.scala 97:16:@132882.4]
  assign rport_io_ins_344 = regs_344_io_out; // @[RegFile.scala 97:16:@132883.4]
  assign rport_io_ins_345 = regs_345_io_out; // @[RegFile.scala 97:16:@132884.4]
  assign rport_io_ins_346 = regs_346_io_out; // @[RegFile.scala 97:16:@132885.4]
  assign rport_io_ins_347 = regs_347_io_out; // @[RegFile.scala 97:16:@132886.4]
  assign rport_io_ins_348 = regs_348_io_out; // @[RegFile.scala 97:16:@132887.4]
  assign rport_io_ins_349 = regs_349_io_out; // @[RegFile.scala 97:16:@132888.4]
  assign rport_io_ins_350 = regs_350_io_out; // @[RegFile.scala 97:16:@132889.4]
  assign rport_io_ins_351 = regs_351_io_out; // @[RegFile.scala 97:16:@132890.4]
  assign rport_io_ins_352 = regs_352_io_out; // @[RegFile.scala 97:16:@132891.4]
  assign rport_io_ins_353 = regs_353_io_out; // @[RegFile.scala 97:16:@132892.4]
  assign rport_io_ins_354 = regs_354_io_out; // @[RegFile.scala 97:16:@132893.4]
  assign rport_io_ins_355 = regs_355_io_out; // @[RegFile.scala 97:16:@132894.4]
  assign rport_io_ins_356 = regs_356_io_out; // @[RegFile.scala 97:16:@132895.4]
  assign rport_io_ins_357 = regs_357_io_out; // @[RegFile.scala 97:16:@132896.4]
  assign rport_io_ins_358 = regs_358_io_out; // @[RegFile.scala 97:16:@132897.4]
  assign rport_io_ins_359 = regs_359_io_out; // @[RegFile.scala 97:16:@132898.4]
  assign rport_io_ins_360 = regs_360_io_out; // @[RegFile.scala 97:16:@132899.4]
  assign rport_io_ins_361 = regs_361_io_out; // @[RegFile.scala 97:16:@132900.4]
  assign rport_io_ins_362 = regs_362_io_out; // @[RegFile.scala 97:16:@132901.4]
  assign rport_io_ins_363 = regs_363_io_out; // @[RegFile.scala 97:16:@132902.4]
  assign rport_io_ins_364 = regs_364_io_out; // @[RegFile.scala 97:16:@132903.4]
  assign rport_io_ins_365 = regs_365_io_out; // @[RegFile.scala 97:16:@132904.4]
  assign rport_io_ins_366 = regs_366_io_out; // @[RegFile.scala 97:16:@132905.4]
  assign rport_io_ins_367 = regs_367_io_out; // @[RegFile.scala 97:16:@132906.4]
  assign rport_io_ins_368 = regs_368_io_out; // @[RegFile.scala 97:16:@132907.4]
  assign rport_io_ins_369 = regs_369_io_out; // @[RegFile.scala 97:16:@132908.4]
  assign rport_io_ins_370 = regs_370_io_out; // @[RegFile.scala 97:16:@132909.4]
  assign rport_io_ins_371 = regs_371_io_out; // @[RegFile.scala 97:16:@132910.4]
  assign rport_io_ins_372 = regs_372_io_out; // @[RegFile.scala 97:16:@132911.4]
  assign rport_io_ins_373 = regs_373_io_out; // @[RegFile.scala 97:16:@132912.4]
  assign rport_io_ins_374 = regs_374_io_out; // @[RegFile.scala 97:16:@132913.4]
  assign rport_io_ins_375 = regs_375_io_out; // @[RegFile.scala 97:16:@132914.4]
  assign rport_io_ins_376 = regs_376_io_out; // @[RegFile.scala 97:16:@132915.4]
  assign rport_io_ins_377 = regs_377_io_out; // @[RegFile.scala 97:16:@132916.4]
  assign rport_io_ins_378 = regs_378_io_out; // @[RegFile.scala 97:16:@132917.4]
  assign rport_io_ins_379 = regs_379_io_out; // @[RegFile.scala 97:16:@132918.4]
  assign rport_io_ins_380 = regs_380_io_out; // @[RegFile.scala 97:16:@132919.4]
  assign rport_io_ins_381 = regs_381_io_out; // @[RegFile.scala 97:16:@132920.4]
  assign rport_io_ins_382 = regs_382_io_out; // @[RegFile.scala 97:16:@132921.4]
  assign rport_io_ins_383 = regs_383_io_out; // @[RegFile.scala 97:16:@132922.4]
  assign rport_io_ins_384 = regs_384_io_out; // @[RegFile.scala 97:16:@132923.4]
  assign rport_io_ins_385 = regs_385_io_out; // @[RegFile.scala 97:16:@132924.4]
  assign rport_io_ins_386 = regs_386_io_out; // @[RegFile.scala 97:16:@132925.4]
  assign rport_io_ins_387 = regs_387_io_out; // @[RegFile.scala 97:16:@132926.4]
  assign rport_io_ins_388 = regs_388_io_out; // @[RegFile.scala 97:16:@132927.4]
  assign rport_io_ins_389 = regs_389_io_out; // @[RegFile.scala 97:16:@132928.4]
  assign rport_io_ins_390 = regs_390_io_out; // @[RegFile.scala 97:16:@132929.4]
  assign rport_io_ins_391 = regs_391_io_out; // @[RegFile.scala 97:16:@132930.4]
  assign rport_io_ins_392 = regs_392_io_out; // @[RegFile.scala 97:16:@132931.4]
  assign rport_io_ins_393 = regs_393_io_out; // @[RegFile.scala 97:16:@132932.4]
  assign rport_io_ins_394 = regs_394_io_out; // @[RegFile.scala 97:16:@132933.4]
  assign rport_io_ins_395 = regs_395_io_out; // @[RegFile.scala 97:16:@132934.4]
  assign rport_io_ins_396 = regs_396_io_out; // @[RegFile.scala 97:16:@132935.4]
  assign rport_io_ins_397 = regs_397_io_out; // @[RegFile.scala 97:16:@132936.4]
  assign rport_io_ins_398 = regs_398_io_out; // @[RegFile.scala 97:16:@132937.4]
  assign rport_io_ins_399 = regs_399_io_out; // @[RegFile.scala 97:16:@132938.4]
  assign rport_io_ins_400 = regs_400_io_out; // @[RegFile.scala 97:16:@132939.4]
  assign rport_io_ins_401 = regs_401_io_out; // @[RegFile.scala 97:16:@132940.4]
  assign rport_io_ins_402 = regs_402_io_out; // @[RegFile.scala 97:16:@132941.4]
  assign rport_io_ins_403 = regs_403_io_out; // @[RegFile.scala 97:16:@132942.4]
  assign rport_io_ins_404 = regs_404_io_out; // @[RegFile.scala 97:16:@132943.4]
  assign rport_io_ins_405 = regs_405_io_out; // @[RegFile.scala 97:16:@132944.4]
  assign rport_io_ins_406 = regs_406_io_out; // @[RegFile.scala 97:16:@132945.4]
  assign rport_io_ins_407 = regs_407_io_out; // @[RegFile.scala 97:16:@132946.4]
  assign rport_io_ins_408 = regs_408_io_out; // @[RegFile.scala 97:16:@132947.4]
  assign rport_io_ins_409 = regs_409_io_out; // @[RegFile.scala 97:16:@132948.4]
  assign rport_io_ins_410 = regs_410_io_out; // @[RegFile.scala 97:16:@132949.4]
  assign rport_io_ins_411 = regs_411_io_out; // @[RegFile.scala 97:16:@132950.4]
  assign rport_io_ins_412 = regs_412_io_out; // @[RegFile.scala 97:16:@132951.4]
  assign rport_io_ins_413 = regs_413_io_out; // @[RegFile.scala 97:16:@132952.4]
  assign rport_io_ins_414 = regs_414_io_out; // @[RegFile.scala 97:16:@132953.4]
  assign rport_io_ins_415 = regs_415_io_out; // @[RegFile.scala 97:16:@132954.4]
  assign rport_io_ins_416 = regs_416_io_out; // @[RegFile.scala 97:16:@132955.4]
  assign rport_io_ins_417 = regs_417_io_out; // @[RegFile.scala 97:16:@132956.4]
  assign rport_io_ins_418 = regs_418_io_out; // @[RegFile.scala 97:16:@132957.4]
  assign rport_io_ins_419 = regs_419_io_out; // @[RegFile.scala 97:16:@132958.4]
  assign rport_io_ins_420 = regs_420_io_out; // @[RegFile.scala 97:16:@132959.4]
  assign rport_io_ins_421 = regs_421_io_out; // @[RegFile.scala 97:16:@132960.4]
  assign rport_io_ins_422 = regs_422_io_out; // @[RegFile.scala 97:16:@132961.4]
  assign rport_io_ins_423 = regs_423_io_out; // @[RegFile.scala 97:16:@132962.4]
  assign rport_io_ins_424 = regs_424_io_out; // @[RegFile.scala 97:16:@132963.4]
  assign rport_io_ins_425 = regs_425_io_out; // @[RegFile.scala 97:16:@132964.4]
  assign rport_io_ins_426 = regs_426_io_out; // @[RegFile.scala 97:16:@132965.4]
  assign rport_io_ins_427 = regs_427_io_out; // @[RegFile.scala 97:16:@132966.4]
  assign rport_io_ins_428 = regs_428_io_out; // @[RegFile.scala 97:16:@132967.4]
  assign rport_io_ins_429 = regs_429_io_out; // @[RegFile.scala 97:16:@132968.4]
  assign rport_io_ins_430 = regs_430_io_out; // @[RegFile.scala 97:16:@132969.4]
  assign rport_io_ins_431 = regs_431_io_out; // @[RegFile.scala 97:16:@132970.4]
  assign rport_io_ins_432 = regs_432_io_out; // @[RegFile.scala 97:16:@132971.4]
  assign rport_io_ins_433 = regs_433_io_out; // @[RegFile.scala 97:16:@132972.4]
  assign rport_io_ins_434 = regs_434_io_out; // @[RegFile.scala 97:16:@132973.4]
  assign rport_io_ins_435 = regs_435_io_out; // @[RegFile.scala 97:16:@132974.4]
  assign rport_io_ins_436 = regs_436_io_out; // @[RegFile.scala 97:16:@132975.4]
  assign rport_io_ins_437 = regs_437_io_out; // @[RegFile.scala 97:16:@132976.4]
  assign rport_io_ins_438 = regs_438_io_out; // @[RegFile.scala 97:16:@132977.4]
  assign rport_io_ins_439 = regs_439_io_out; // @[RegFile.scala 97:16:@132978.4]
  assign rport_io_ins_440 = regs_440_io_out; // @[RegFile.scala 97:16:@132979.4]
  assign rport_io_ins_441 = regs_441_io_out; // @[RegFile.scala 97:16:@132980.4]
  assign rport_io_ins_442 = regs_442_io_out; // @[RegFile.scala 97:16:@132981.4]
  assign rport_io_ins_443 = regs_443_io_out; // @[RegFile.scala 97:16:@132982.4]
  assign rport_io_ins_444 = regs_444_io_out; // @[RegFile.scala 97:16:@132983.4]
  assign rport_io_ins_445 = regs_445_io_out; // @[RegFile.scala 97:16:@132984.4]
  assign rport_io_ins_446 = regs_446_io_out; // @[RegFile.scala 97:16:@132985.4]
  assign rport_io_ins_447 = regs_447_io_out; // @[RegFile.scala 97:16:@132986.4]
  assign rport_io_ins_448 = regs_448_io_out; // @[RegFile.scala 97:16:@132987.4]
  assign rport_io_ins_449 = regs_449_io_out; // @[RegFile.scala 97:16:@132988.4]
  assign rport_io_ins_450 = regs_450_io_out; // @[RegFile.scala 97:16:@132989.4]
  assign rport_io_ins_451 = regs_451_io_out; // @[RegFile.scala 97:16:@132990.4]
  assign rport_io_ins_452 = regs_452_io_out; // @[RegFile.scala 97:16:@132991.4]
  assign rport_io_ins_453 = regs_453_io_out; // @[RegFile.scala 97:16:@132992.4]
  assign rport_io_ins_454 = regs_454_io_out; // @[RegFile.scala 97:16:@132993.4]
  assign rport_io_ins_455 = regs_455_io_out; // @[RegFile.scala 97:16:@132994.4]
  assign rport_io_ins_456 = regs_456_io_out; // @[RegFile.scala 97:16:@132995.4]
  assign rport_io_ins_457 = regs_457_io_out; // @[RegFile.scala 97:16:@132996.4]
  assign rport_io_ins_458 = regs_458_io_out; // @[RegFile.scala 97:16:@132997.4]
  assign rport_io_ins_459 = regs_459_io_out; // @[RegFile.scala 97:16:@132998.4]
  assign rport_io_ins_460 = regs_460_io_out; // @[RegFile.scala 97:16:@132999.4]
  assign rport_io_ins_461 = regs_461_io_out; // @[RegFile.scala 97:16:@133000.4]
  assign rport_io_ins_462 = regs_462_io_out; // @[RegFile.scala 97:16:@133001.4]
  assign rport_io_ins_463 = regs_463_io_out; // @[RegFile.scala 97:16:@133002.4]
  assign rport_io_ins_464 = regs_464_io_out; // @[RegFile.scala 97:16:@133003.4]
  assign rport_io_ins_465 = regs_465_io_out; // @[RegFile.scala 97:16:@133004.4]
  assign rport_io_ins_466 = regs_466_io_out; // @[RegFile.scala 97:16:@133005.4]
  assign rport_io_ins_467 = regs_467_io_out; // @[RegFile.scala 97:16:@133006.4]
  assign rport_io_ins_468 = regs_468_io_out; // @[RegFile.scala 97:16:@133007.4]
  assign rport_io_ins_469 = regs_469_io_out; // @[RegFile.scala 97:16:@133008.4]
  assign rport_io_ins_470 = regs_470_io_out; // @[RegFile.scala 97:16:@133009.4]
  assign rport_io_ins_471 = regs_471_io_out; // @[RegFile.scala 97:16:@133010.4]
  assign rport_io_ins_472 = regs_472_io_out; // @[RegFile.scala 97:16:@133011.4]
  assign rport_io_ins_473 = regs_473_io_out; // @[RegFile.scala 97:16:@133012.4]
  assign rport_io_ins_474 = regs_474_io_out; // @[RegFile.scala 97:16:@133013.4]
  assign rport_io_ins_475 = regs_475_io_out; // @[RegFile.scala 97:16:@133014.4]
  assign rport_io_ins_476 = regs_476_io_out; // @[RegFile.scala 97:16:@133015.4]
  assign rport_io_ins_477 = regs_477_io_out; // @[RegFile.scala 97:16:@133016.4]
  assign rport_io_ins_478 = regs_478_io_out; // @[RegFile.scala 97:16:@133017.4]
  assign rport_io_ins_479 = regs_479_io_out; // @[RegFile.scala 97:16:@133018.4]
  assign rport_io_ins_480 = regs_480_io_out; // @[RegFile.scala 97:16:@133019.4]
  assign rport_io_ins_481 = regs_481_io_out; // @[RegFile.scala 97:16:@133020.4]
  assign rport_io_ins_482 = regs_482_io_out; // @[RegFile.scala 97:16:@133021.4]
  assign rport_io_ins_483 = regs_483_io_out; // @[RegFile.scala 97:16:@133022.4]
  assign rport_io_ins_484 = regs_484_io_out; // @[RegFile.scala 97:16:@133023.4]
  assign rport_io_ins_485 = regs_485_io_out; // @[RegFile.scala 97:16:@133024.4]
  assign rport_io_ins_486 = regs_486_io_out; // @[RegFile.scala 97:16:@133025.4]
  assign rport_io_ins_487 = regs_487_io_out; // @[RegFile.scala 97:16:@133026.4]
  assign rport_io_ins_488 = regs_488_io_out; // @[RegFile.scala 97:16:@133027.4]
  assign rport_io_ins_489 = regs_489_io_out; // @[RegFile.scala 97:16:@133028.4]
  assign rport_io_ins_490 = regs_490_io_out; // @[RegFile.scala 97:16:@133029.4]
  assign rport_io_ins_491 = regs_491_io_out; // @[RegFile.scala 97:16:@133030.4]
  assign rport_io_ins_492 = regs_492_io_out; // @[RegFile.scala 97:16:@133031.4]
  assign rport_io_ins_493 = regs_493_io_out; // @[RegFile.scala 97:16:@133032.4]
  assign rport_io_ins_494 = regs_494_io_out; // @[RegFile.scala 97:16:@133033.4]
  assign rport_io_ins_495 = regs_495_io_out; // @[RegFile.scala 97:16:@133034.4]
  assign rport_io_ins_496 = regs_496_io_out; // @[RegFile.scala 97:16:@133035.4]
  assign rport_io_ins_497 = regs_497_io_out; // @[RegFile.scala 97:16:@133036.4]
  assign rport_io_ins_498 = regs_498_io_out; // @[RegFile.scala 97:16:@133037.4]
  assign rport_io_ins_499 = regs_499_io_out; // @[RegFile.scala 97:16:@133038.4]
  assign rport_io_ins_500 = regs_500_io_out; // @[RegFile.scala 97:16:@133039.4]
  assign rport_io_ins_501 = regs_501_io_out; // @[RegFile.scala 97:16:@133040.4]
  assign rport_io_ins_502 = regs_502_io_out; // @[RegFile.scala 97:16:@133041.4]
  assign rport_io_sel = io_raddr[8:0]; // @[RegFile.scala 106:18:@133042.4]
endmodule
module RetimeWrapper_810( // @[:@133066.2]
  input         clock, // @[:@133067.4]
  input         reset, // @[:@133068.4]
  input  [39:0] io_in, // @[:@133069.4]
  output [39:0] io_out // @[:@133069.4]
);
  wire [39:0] sr_out; // @[RetimeShiftRegister.scala 15:20:@133071.4]
  wire [39:0] sr_in; // @[RetimeShiftRegister.scala 15:20:@133071.4]
  wire [39:0] sr_init; // @[RetimeShiftRegister.scala 15:20:@133071.4]
  wire  sr_flow; // @[RetimeShiftRegister.scala 15:20:@133071.4]
  wire  sr_reset; // @[RetimeShiftRegister.scala 15:20:@133071.4]
  wire  sr_clock; // @[RetimeShiftRegister.scala 15:20:@133071.4]
  RetimeShiftRegister #(.WIDTH(40), .STAGES(1)) sr ( // @[RetimeShiftRegister.scala 15:20:@133071.4]
    .out(sr_out),
    .in(sr_in),
    .init(sr_init),
    .flow(sr_flow),
    .reset(sr_reset),
    .clock(sr_clock)
  );
  assign io_out = sr_out; // @[RetimeShiftRegister.scala 21:12:@133084.4]
  assign sr_in = io_in; // @[RetimeShiftRegister.scala 20:14:@133083.4]
  assign sr_init = 40'h0; // @[RetimeShiftRegister.scala 19:16:@133082.4]
  assign sr_flow = 1'h1; // @[RetimeShiftRegister.scala 18:16:@133081.4]
  assign sr_reset = reset; // @[RetimeShiftRegister.scala 17:17:@133080.4]
  assign sr_clock = clock; // @[RetimeShiftRegister.scala 16:17:@133078.4]
endmodule
module FringeFF_503( // @[:@133086.2]
  input         clock, // @[:@133087.4]
  input         reset, // @[:@133088.4]
  input  [39:0] io_in, // @[:@133089.4]
  output [39:0] io_out, // @[:@133089.4]
  input         io_enable // @[:@133089.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@133092.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@133092.4]
  wire [39:0] RetimeWrapper_io_in; // @[package.scala 93:22:@133092.4]
  wire [39:0] RetimeWrapper_io_out; // @[package.scala 93:22:@133092.4]
  wire [39:0] _T_18; // @[package.scala 96:25:@133097.4 package.scala 96:25:@133098.4]
  RetimeWrapper_810 RetimeWrapper ( // @[package.scala 93:22:@133092.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@133097.4 package.scala 96:25:@133098.4]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@133109.4]
  assign RetimeWrapper_clock = clock; // @[:@133093.4]
  assign RetimeWrapper_reset = reset; // @[:@133094.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _T_18; // @[package.scala 94:16:@133095.4]
endmodule
module FringeCounter( // @[:@133111.2]
  input   clock, // @[:@133112.4]
  input   reset, // @[:@133113.4]
  input   io_enable, // @[:@133114.4]
  output  io_done // @[:@133114.4]
);
  wire  reg$_clock; // @[FringeCounter.scala 24:19:@133116.4]
  wire  reg$_reset; // @[FringeCounter.scala 24:19:@133116.4]
  wire [39:0] reg$_io_in; // @[FringeCounter.scala 24:19:@133116.4]
  wire [39:0] reg$_io_out; // @[FringeCounter.scala 24:19:@133116.4]
  wire  reg$_io_enable; // @[FringeCounter.scala 24:19:@133116.4]
  wire [40:0] count; // @[Cat.scala 30:58:@133123.4]
  wire [41:0] _T_25; // @[FringeCounter.scala 31:22:@133124.4]
  wire [40:0] newval; // @[FringeCounter.scala 31:22:@133125.4]
  wire  isMax; // @[FringeCounter.scala 32:22:@133126.4]
  wire [40:0] next; // @[FringeCounter.scala 33:17:@133128.4]
  FringeFF_503 reg$ ( // @[FringeCounter.scala 24:19:@133116.4]
    .clock(reg$_clock),
    .reset(reg$_reset),
    .io_in(reg$_io_in),
    .io_out(reg$_io_out),
    .io_enable(reg$_io_enable)
  );
  assign count = {1'h0,reg$_io_out}; // @[Cat.scala 30:58:@133123.4]
  assign _T_25 = count + 41'h1; // @[FringeCounter.scala 31:22:@133124.4]
  assign newval = count + 41'h1; // @[FringeCounter.scala 31:22:@133125.4]
  assign isMax = newval >= 41'h2cb417800; // @[FringeCounter.scala 32:22:@133126.4]
  assign next = isMax ? count : newval; // @[FringeCounter.scala 33:17:@133128.4]
  assign io_done = io_enable & isMax; // @[FringeCounter.scala 43:11:@133139.4]
  assign reg$_clock = clock; // @[:@133117.4]
  assign reg$_reset = reset; // @[:@133118.4]
  assign reg$_io_in = next[39:0]; // @[FringeCounter.scala 35:15:@133130.6 FringeCounter.scala 37:15:@133133.6]
  assign reg$_io_enable = io_enable; // @[FringeCounter.scala 27:17:@133121.4]
endmodule
module FringeFF_504( // @[:@133173.2]
  input   clock, // @[:@133174.4]
  input   reset, // @[:@133175.4]
  input   io_in, // @[:@133176.4]
  input   io_reset, // @[:@133176.4]
  output  io_out, // @[:@133176.4]
  input   io_enable // @[:@133176.4]
);
  wire  RetimeWrapper_clock; // @[package.scala 93:22:@133179.4]
  wire  RetimeWrapper_reset; // @[package.scala 93:22:@133179.4]
  wire  RetimeWrapper_io_flow; // @[package.scala 93:22:@133179.4]
  wire  RetimeWrapper_io_in; // @[package.scala 93:22:@133179.4]
  wire  RetimeWrapper_io_out; // @[package.scala 93:22:@133179.4]
  wire  _T_18; // @[package.scala 96:25:@133184.4 package.scala 96:25:@133185.4]
  wire  _GEN_0; // @[FringeFF.scala 21:27:@133190.6]
  RetimeWrapper RetimeWrapper ( // @[package.scala 93:22:@133179.4]
    .clock(RetimeWrapper_clock),
    .reset(RetimeWrapper_reset),
    .io_flow(RetimeWrapper_io_flow),
    .io_in(RetimeWrapper_io_in),
    .io_out(RetimeWrapper_io_out)
  );
  assign _T_18 = RetimeWrapper_io_out; // @[package.scala 96:25:@133184.4 package.scala 96:25:@133185.4]
  assign _GEN_0 = io_reset ? 1'h0 : _T_18; // @[FringeFF.scala 21:27:@133190.6]
  assign io_out = RetimeWrapper_io_out; // @[FringeFF.scala 26:12:@133196.4]
  assign RetimeWrapper_clock = clock; // @[:@133180.4]
  assign RetimeWrapper_reset = reset; // @[:@133181.4]
  assign RetimeWrapper_io_flow = 1'h1; // @[package.scala 95:18:@133183.4]
  assign RetimeWrapper_io_in = io_enable ? io_in : _GEN_0; // @[package.scala 94:16:@133182.4]
endmodule
module Depulser( // @[:@133198.2]
  input   clock, // @[:@133199.4]
  input   reset, // @[:@133200.4]
  input   io_in, // @[:@133201.4]
  input   io_rst, // @[:@133201.4]
  output  io_out // @[:@133201.4]
);
  wire  r_clock; // @[Depulser.scala 14:17:@133203.4]
  wire  r_reset; // @[Depulser.scala 14:17:@133203.4]
  wire  r_io_in; // @[Depulser.scala 14:17:@133203.4]
  wire  r_io_reset; // @[Depulser.scala 14:17:@133203.4]
  wire  r_io_out; // @[Depulser.scala 14:17:@133203.4]
  wire  r_io_enable; // @[Depulser.scala 14:17:@133203.4]
  FringeFF_504 r ( // @[Depulser.scala 14:17:@133203.4]
    .clock(r_clock),
    .reset(r_reset),
    .io_in(r_io_in),
    .io_reset(r_io_reset),
    .io_out(r_io_out),
    .io_enable(r_io_enable)
  );
  assign io_out = r_io_out; // @[Depulser.scala 19:10:@133212.4]
  assign r_clock = clock; // @[:@133204.4]
  assign r_reset = reset; // @[:@133205.4]
  assign r_io_in = io_rst ? 1'h0 : io_in; // @[Depulser.scala 15:11:@133207.4]
  assign r_io_reset = io_rst; // @[Depulser.scala 18:14:@133211.4]
  assign r_io_enable = io_in | io_rst; // @[Depulser.scala 17:15:@133210.4]
endmodule
module Fringe( // @[:@133214.2]
  input         clock, // @[:@133215.4]
  input         reset, // @[:@133216.4]
  input  [31:0] io_raddr, // @[:@133217.4]
  input         io_wen, // @[:@133217.4]
  input  [31:0] io_waddr, // @[:@133217.4]
  input  [63:0] io_wdata, // @[:@133217.4]
  output [63:0] io_rdata, // @[:@133217.4]
  output        io_enable, // @[:@133217.4]
  input         io_done, // @[:@133217.4]
  output        io_reset, // @[:@133217.4]
  output [63:0] io_argIns_0, // @[:@133217.4]
  output [63:0] io_argIns_1, // @[:@133217.4]
  input         io_argOuts_0_valid, // @[:@133217.4]
  input  [63:0] io_argOuts_0_bits, // @[:@133217.4]
  output        io_memStreams_stores_0_cmd_ready, // @[:@133217.4]
  input         io_memStreams_stores_0_cmd_valid, // @[:@133217.4]
  input  [63:0] io_memStreams_stores_0_cmd_bits_addr, // @[:@133217.4]
  input  [31:0] io_memStreams_stores_0_cmd_bits_size, // @[:@133217.4]
  output        io_memStreams_stores_0_data_ready, // @[:@133217.4]
  input         io_memStreams_stores_0_data_valid, // @[:@133217.4]
  input  [31:0] io_memStreams_stores_0_data_bits_wdata_0, // @[:@133217.4]
  input         io_memStreams_stores_0_data_bits_wstrb, // @[:@133217.4]
  input         io_memStreams_stores_0_wresp_ready, // @[:@133217.4]
  output        io_memStreams_stores_0_wresp_valid, // @[:@133217.4]
  output        io_memStreams_stores_0_wresp_bits, // @[:@133217.4]
  input         io_dram_0_cmd_ready, // @[:@133217.4]
  output        io_dram_0_cmd_valid, // @[:@133217.4]
  output [63:0] io_dram_0_cmd_bits_addr, // @[:@133217.4]
  output [31:0] io_dram_0_cmd_bits_size, // @[:@133217.4]
  output        io_dram_0_cmd_bits_isWr, // @[:@133217.4]
  output [31:0] io_dram_0_cmd_bits_tag, // @[:@133217.4]
  input         io_dram_0_wdata_ready, // @[:@133217.4]
  output        io_dram_0_wdata_valid, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_0, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_1, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_2, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_3, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_4, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_5, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_6, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_7, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_8, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_9, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_10, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_11, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_12, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_13, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_14, // @[:@133217.4]
  output [31:0] io_dram_0_wdata_bits_wdata_15, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_0, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_1, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_2, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_3, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_4, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_5, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_6, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_7, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_8, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_9, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_10, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_11, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_12, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_13, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_14, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_15, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_16, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_17, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_18, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_19, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_20, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_21, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_22, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_23, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_24, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_25, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_26, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_27, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_28, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_29, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_30, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_31, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_32, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_33, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_34, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_35, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_36, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_37, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_38, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_39, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_40, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_41, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_42, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_43, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_44, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_45, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_46, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_47, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_48, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_49, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_50, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_51, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_52, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_53, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_54, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_55, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_56, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_57, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_58, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_59, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_60, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_61, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_62, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wstrb_63, // @[:@133217.4]
  output        io_dram_0_wdata_bits_wlast, // @[:@133217.4]
  output        io_dram_0_rresp_ready, // @[:@133217.4]
  output        io_dram_0_wresp_ready, // @[:@133217.4]
  input         io_dram_0_wresp_valid, // @[:@133217.4]
  input  [31:0] io_dram_0_wresp_bits_tag, // @[:@133217.4]
  input         io_dram_1_cmd_ready, // @[:@133217.4]
  output        io_dram_1_cmd_valid, // @[:@133217.4]
  output [63:0] io_dram_1_cmd_bits_addr, // @[:@133217.4]
  output [31:0] io_dram_1_cmd_bits_size, // @[:@133217.4]
  output        io_dram_1_cmd_bits_isWr, // @[:@133217.4]
  output [31:0] io_dram_1_cmd_bits_tag, // @[:@133217.4]
  input         io_dram_1_wdata_ready, // @[:@133217.4]
  output        io_dram_1_wdata_valid, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_0, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_1, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_2, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_3, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_4, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_5, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_6, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_7, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_8, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_9, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_10, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_11, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_12, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_13, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_14, // @[:@133217.4]
  output [31:0] io_dram_1_wdata_bits_wdata_15, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_0, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_1, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_2, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_3, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_4, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_5, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_6, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_7, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_8, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_9, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_10, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_11, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_12, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_13, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_14, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_15, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_16, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_17, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_18, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_19, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_20, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_21, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_22, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_23, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_24, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_25, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_26, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_27, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_28, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_29, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_30, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_31, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_32, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_33, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_34, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_35, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_36, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_37, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_38, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_39, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_40, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_41, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_42, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_43, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_44, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_45, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_46, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_47, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_48, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_49, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_50, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_51, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_52, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_53, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_54, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_55, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_56, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_57, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_58, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_59, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_60, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_61, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_62, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wstrb_63, // @[:@133217.4]
  output        io_dram_1_wdata_bits_wlast, // @[:@133217.4]
  output        io_dram_1_rresp_ready, // @[:@133217.4]
  output        io_dram_1_wresp_ready, // @[:@133217.4]
  input         io_dram_1_wresp_valid, // @[:@133217.4]
  input  [31:0] io_dram_1_wresp_bits_tag, // @[:@133217.4]
  input         io_dram_2_cmd_ready, // @[:@133217.4]
  output        io_dram_2_cmd_valid, // @[:@133217.4]
  output [63:0] io_dram_2_cmd_bits_addr, // @[:@133217.4]
  output [31:0] io_dram_2_cmd_bits_size, // @[:@133217.4]
  output        io_dram_2_cmd_bits_isWr, // @[:@133217.4]
  output [31:0] io_dram_2_cmd_bits_tag, // @[:@133217.4]
  input         io_dram_2_wdata_ready, // @[:@133217.4]
  output        io_dram_2_wdata_valid, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_0, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_1, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_2, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_3, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_4, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_5, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_6, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_7, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_8, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_9, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_10, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_11, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_12, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_13, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_14, // @[:@133217.4]
  output [31:0] io_dram_2_wdata_bits_wdata_15, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_0, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_1, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_2, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_3, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_4, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_5, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_6, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_7, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_8, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_9, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_10, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_11, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_12, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_13, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_14, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_15, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_16, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_17, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_18, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_19, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_20, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_21, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_22, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_23, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_24, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_25, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_26, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_27, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_28, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_29, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_30, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_31, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_32, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_33, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_34, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_35, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_36, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_37, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_38, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_39, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_40, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_41, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_42, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_43, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_44, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_45, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_46, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_47, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_48, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_49, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_50, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_51, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_52, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_53, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_54, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_55, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_56, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_57, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_58, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_59, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_60, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_61, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_62, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wstrb_63, // @[:@133217.4]
  output        io_dram_2_wdata_bits_wlast, // @[:@133217.4]
  output        io_dram_2_rresp_ready, // @[:@133217.4]
  output        io_dram_2_wresp_ready, // @[:@133217.4]
  input         io_dram_2_wresp_valid, // @[:@133217.4]
  input  [31:0] io_dram_2_wresp_bits_tag, // @[:@133217.4]
  input         io_dram_3_cmd_ready, // @[:@133217.4]
  output        io_dram_3_cmd_valid, // @[:@133217.4]
  output [63:0] io_dram_3_cmd_bits_addr, // @[:@133217.4]
  output [31:0] io_dram_3_cmd_bits_size, // @[:@133217.4]
  output        io_dram_3_cmd_bits_isWr, // @[:@133217.4]
  output [31:0] io_dram_3_cmd_bits_tag, // @[:@133217.4]
  input         io_dram_3_wdata_ready, // @[:@133217.4]
  output        io_dram_3_wdata_valid, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_0, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_1, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_2, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_3, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_4, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_5, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_6, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_7, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_8, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_9, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_10, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_11, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_12, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_13, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_14, // @[:@133217.4]
  output [31:0] io_dram_3_wdata_bits_wdata_15, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_0, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_1, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_2, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_3, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_4, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_5, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_6, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_7, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_8, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_9, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_10, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_11, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_12, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_13, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_14, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_15, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_16, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_17, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_18, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_19, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_20, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_21, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_22, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_23, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_24, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_25, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_26, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_27, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_28, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_29, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_30, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_31, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_32, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_33, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_34, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_35, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_36, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_37, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_38, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_39, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_40, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_41, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_42, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_43, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_44, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_45, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_46, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_47, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_48, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_49, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_50, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_51, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_52, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_53, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_54, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_55, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_56, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_57, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_58, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_59, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_60, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_61, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_62, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wstrb_63, // @[:@133217.4]
  output        io_dram_3_wdata_bits_wlast, // @[:@133217.4]
  output        io_dram_3_rresp_ready, // @[:@133217.4]
  output        io_dram_3_wresp_ready, // @[:@133217.4]
  input         io_dram_3_wresp_valid, // @[:@133217.4]
  input  [31:0] io_dram_3_wresp_bits_tag, // @[:@133217.4]
  input         io_heap_0_req_valid, // @[:@133217.4]
  input         io_heap_0_req_bits_allocDealloc, // @[:@133217.4]
  input  [63:0] io_heap_0_req_bits_sizeAddr, // @[:@133217.4]
  output        io_heap_0_resp_valid, // @[:@133217.4]
  output        io_heap_0_resp_bits_allocDealloc, // @[:@133217.4]
  output [63:0] io_heap_0_resp_bits_sizeAddr // @[:@133217.4]
);
  wire  dramArbs_0_clock; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_reset; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_enable; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_app_stores_0_cmd_valid; // @[Fringe.scala 91:25:@133223.4]
  wire [63:0] dramArbs_0_io_app_stores_0_cmd_bits_addr; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_app_stores_0_cmd_bits_size; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_app_stores_0_data_valid; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_app_stores_0_data_bits_wdata_0; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_app_stores_0_data_bits_wstrb; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_app_stores_0_wresp_ready; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_cmd_ready; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 91:25:@133223.4]
  wire [63:0] dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_ready; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_0_io_dram_wresp_valid; // @[Fringe.scala 91:25:@133223.4]
  wire [31:0] dramArbs_0_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@133223.4]
  wire  dramArbs_1_clock; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_reset; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_enable; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_cmd_ready; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 91:25:@134216.4]
  wire [63:0] dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_ready; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_1_io_dram_wresp_valid; // @[Fringe.scala 91:25:@134216.4]
  wire [31:0] dramArbs_1_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@134216.4]
  wire  dramArbs_2_clock; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_reset; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_enable; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_cmd_ready; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 91:25:@135176.4]
  wire [63:0] dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_ready; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_2_io_dram_wresp_valid; // @[Fringe.scala 91:25:@135176.4]
  wire [31:0] dramArbs_2_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@135176.4]
  wire  dramArbs_3_clock; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_reset; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_enable; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_cmd_ready; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 91:25:@136136.4]
  wire [63:0] dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_ready; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 91:25:@136136.4]
  wire  dramArbs_3_io_dram_wresp_valid; // @[Fringe.scala 91:25:@136136.4]
  wire [31:0] dramArbs_3_io_dram_wresp_bits_tag; // @[Fringe.scala 91:25:@136136.4]
  wire  heap_io_accel_0_req_valid; // @[Fringe.scala 107:20:@137096.4]
  wire  heap_io_accel_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@137096.4]
  wire [63:0] heap_io_accel_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@137096.4]
  wire  heap_io_accel_0_resp_valid; // @[Fringe.scala 107:20:@137096.4]
  wire  heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@137096.4]
  wire [63:0] heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@137096.4]
  wire  heap_io_host_0_req_valid; // @[Fringe.scala 107:20:@137096.4]
  wire  heap_io_host_0_req_bits_allocDealloc; // @[Fringe.scala 107:20:@137096.4]
  wire [63:0] heap_io_host_0_req_bits_sizeAddr; // @[Fringe.scala 107:20:@137096.4]
  wire  heap_io_host_0_resp_valid; // @[Fringe.scala 107:20:@137096.4]
  wire  heap_io_host_0_resp_bits_allocDealloc; // @[Fringe.scala 107:20:@137096.4]
  wire [63:0] heap_io_host_0_resp_bits_sizeAddr; // @[Fringe.scala 107:20:@137096.4]
  wire  regs_clock; // @[Fringe.scala 116:20:@137105.4]
  wire  regs_reset; // @[Fringe.scala 116:20:@137105.4]
  wire [31:0] regs_io_raddr; // @[Fringe.scala 116:20:@137105.4]
  wire  regs_io_wen; // @[Fringe.scala 116:20:@137105.4]
  wire [31:0] regs_io_waddr; // @[Fringe.scala 116:20:@137105.4]
  wire [63:0] regs_io_wdata; // @[Fringe.scala 116:20:@137105.4]
  wire [63:0] regs_io_rdata; // @[Fringe.scala 116:20:@137105.4]
  wire  regs_io_reset; // @[Fringe.scala 116:20:@137105.4]
  wire [63:0] regs_io_argIns_0; // @[Fringe.scala 116:20:@137105.4]
  wire [63:0] regs_io_argIns_1; // @[Fringe.scala 116:20:@137105.4]
  wire [63:0] regs_io_argIns_2; // @[Fringe.scala 116:20:@137105.4]
  wire [63:0] regs_io_argIns_3; // @[Fringe.scala 116:20:@137105.4]
  wire  regs_io_argOuts_0_valid; // @[Fringe.scala 116:20:@137105.4]
  wire [63:0] regs_io_argOuts_0_bits; // @[Fringe.scala 116:20:@137105.4]
  wire  regs_io_argOuts_1_valid; // @[Fringe.scala 116:20:@137105.4]
  wire [63:0] regs_io_argOuts_1_bits; // @[Fringe.scala 116:20:@137105.4]
  wire  timeoutCtr_clock; // @[Fringe.scala 143:26:@139155.4]
  wire  timeoutCtr_reset; // @[Fringe.scala 143:26:@139155.4]
  wire  timeoutCtr_io_enable; // @[Fringe.scala 143:26:@139155.4]
  wire  timeoutCtr_io_done; // @[Fringe.scala 143:26:@139155.4]
  wire  depulser_clock; // @[Fringe.scala 153:24:@139174.4]
  wire  depulser_reset; // @[Fringe.scala 153:24:@139174.4]
  wire  depulser_io_in; // @[Fringe.scala 153:24:@139174.4]
  wire  depulser_io_rst; // @[Fringe.scala 153:24:@139174.4]
  wire  depulser_io_out; // @[Fringe.scala 153:24:@139174.4]
  wire [63:0] _T_1020; // @[:@139132.4 :@139133.4]
  wire  curStatus_done; // @[Fringe.scala 133:45:@139134.4]
  wire  curStatus_timeout; // @[Fringe.scala 133:45:@139136.4]
  wire [2:0] curStatus_allocDealloc; // @[Fringe.scala 133:45:@139138.4]
  wire [58:0] curStatus_sizeAddr; // @[Fringe.scala 133:45:@139140.4]
  wire  _T_1025; // @[Fringe.scala 134:28:@139142.4]
  wire  _T_1029; // @[Fringe.scala 134:42:@139144.4]
  wire  _T_1030; // @[Fringe.scala 135:27:@139146.4]
  wire [63:0] _T_1040; // @[Fringe.scala 156:22:@139182.4]
  reg  _T_1047; // @[package.scala 152:20:@139185.4]
  reg [31:0] _RAND_0;
  wire  _T_1048; // @[package.scala 153:13:@139187.4]
  wire  _T_1049; // @[package.scala 153:8:@139188.4]
  wire  _T_1052; // @[Fringe.scala 160:55:@139192.4]
  wire  status_bits_done; // @[Fringe.scala 160:26:@139193.4]
  wire  _T_1055; // @[Fringe.scala 161:58:@139196.4]
  wire  status_bits_timeout; // @[Fringe.scala 161:29:@139197.4]
  wire [1:0] _T_1059; // @[Fringe.scala 162:57:@139199.4]
  wire [1:0] _T_1061; // @[Fringe.scala 162:34:@139200.4]
  wire [63:0] _T_1063; // @[Fringe.scala 163:30:@139202.4]
  wire [1:0] _T_1064; // @[Fringe.scala 171:37:@139205.4]
  wire [58:0] status_bits_sizeAddr; // @[Fringe.scala 158:20:@139184.4 Fringe.scala 163:24:@139203.4]
  wire [2:0] status_bits_allocDealloc; // @[Fringe.scala 158:20:@139184.4 Fringe.scala 162:28:@139201.4]
  wire [61:0] _T_1065; // @[Fringe.scala 171:37:@139206.4]
  wire  alloc; // @[Fringe.scala 202:38:@140836.4]
  wire  dealloc; // @[Fringe.scala 203:40:@140837.4]
  wire  _T_1569; // @[Fringe.scala 204:37:@140838.4]
  reg  _T_1572; // @[package.scala 152:20:@140839.4]
  reg [31:0] _RAND_1;
  wire  _T_1573; // @[package.scala 153:13:@140841.4]
  DRAMArbiter dramArbs_0 ( // @[Fringe.scala 91:25:@133223.4]
    .clock(dramArbs_0_clock),
    .reset(dramArbs_0_reset),
    .io_enable(dramArbs_0_io_enable),
    .io_app_stores_0_cmd_ready(dramArbs_0_io_app_stores_0_cmd_ready),
    .io_app_stores_0_cmd_valid(dramArbs_0_io_app_stores_0_cmd_valid),
    .io_app_stores_0_cmd_bits_addr(dramArbs_0_io_app_stores_0_cmd_bits_addr),
    .io_app_stores_0_cmd_bits_size(dramArbs_0_io_app_stores_0_cmd_bits_size),
    .io_app_stores_0_data_ready(dramArbs_0_io_app_stores_0_data_ready),
    .io_app_stores_0_data_valid(dramArbs_0_io_app_stores_0_data_valid),
    .io_app_stores_0_data_bits_wdata_0(dramArbs_0_io_app_stores_0_data_bits_wdata_0),
    .io_app_stores_0_data_bits_wstrb(dramArbs_0_io_app_stores_0_data_bits_wstrb),
    .io_app_stores_0_wresp_ready(dramArbs_0_io_app_stores_0_wresp_ready),
    .io_app_stores_0_wresp_valid(dramArbs_0_io_app_stores_0_wresp_valid),
    .io_app_stores_0_wresp_bits(dramArbs_0_io_app_stores_0_wresp_bits),
    .io_dram_cmd_ready(dramArbs_0_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_0_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_0_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_0_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_0_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_0_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_0_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_0_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_0_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_0_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_0_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_0_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_0_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_0_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_0_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_0_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_0_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_0_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_0_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_0_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_0_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_0_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_0_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_0_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_0_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_0_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_0_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_0_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_0_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_0_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_0_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_0_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_0_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_0_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_0_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_0_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_0_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_0_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_0_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_0_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_0_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_0_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_0_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_0_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_0_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_0_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_0_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_0_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_0_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_0_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_0_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_0_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_0_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_0_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_0_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_0_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_0_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_0_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_0_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_0_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_0_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_0_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_0_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_0_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_0_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_0_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_0_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_0_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_0_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_0_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_0_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_0_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_0_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_0_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_0_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_0_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_0_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_0_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_0_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_0_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_0_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_0_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_0_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_0_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_0_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_0_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_0_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_0_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_0_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_0_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_0_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_0_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_0_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_1 ( // @[Fringe.scala 91:25:@134216.4]
    .clock(dramArbs_1_clock),
    .reset(dramArbs_1_reset),
    .io_enable(dramArbs_1_io_enable),
    .io_dram_cmd_ready(dramArbs_1_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_1_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_1_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_1_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_1_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_1_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_1_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_1_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_1_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_1_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_1_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_1_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_1_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_1_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_1_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_1_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_1_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_1_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_1_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_1_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_1_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_1_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_1_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_1_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_1_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_1_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_1_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_1_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_1_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_1_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_1_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_1_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_1_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_1_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_1_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_1_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_1_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_1_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_1_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_1_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_1_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_1_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_1_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_1_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_1_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_1_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_1_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_1_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_1_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_1_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_1_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_1_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_1_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_1_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_1_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_1_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_1_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_1_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_1_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_1_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_1_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_1_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_1_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_1_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_1_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_1_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_1_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_1_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_1_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_1_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_1_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_1_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_1_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_1_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_1_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_1_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_1_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_1_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_1_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_1_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_1_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_1_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_1_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_1_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_1_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_1_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_1_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_1_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_1_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_1_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_1_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_1_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_1_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_2 ( // @[Fringe.scala 91:25:@135176.4]
    .clock(dramArbs_2_clock),
    .reset(dramArbs_2_reset),
    .io_enable(dramArbs_2_io_enable),
    .io_dram_cmd_ready(dramArbs_2_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_2_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_2_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_2_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_2_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_2_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_2_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_2_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_2_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_2_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_2_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_2_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_2_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_2_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_2_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_2_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_2_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_2_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_2_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_2_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_2_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_2_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_2_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_2_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_2_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_2_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_2_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_2_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_2_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_2_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_2_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_2_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_2_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_2_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_2_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_2_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_2_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_2_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_2_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_2_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_2_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_2_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_2_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_2_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_2_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_2_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_2_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_2_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_2_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_2_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_2_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_2_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_2_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_2_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_2_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_2_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_2_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_2_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_2_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_2_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_2_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_2_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_2_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_2_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_2_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_2_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_2_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_2_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_2_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_2_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_2_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_2_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_2_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_2_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_2_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_2_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_2_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_2_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_2_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_2_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_2_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_2_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_2_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_2_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_2_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_2_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_2_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_2_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_2_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_2_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_2_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_2_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_2_io_dram_wresp_bits_tag)
  );
  DRAMArbiter_1 dramArbs_3 ( // @[Fringe.scala 91:25:@136136.4]
    .clock(dramArbs_3_clock),
    .reset(dramArbs_3_reset),
    .io_enable(dramArbs_3_io_enable),
    .io_dram_cmd_ready(dramArbs_3_io_dram_cmd_ready),
    .io_dram_cmd_valid(dramArbs_3_io_dram_cmd_valid),
    .io_dram_cmd_bits_addr(dramArbs_3_io_dram_cmd_bits_addr),
    .io_dram_cmd_bits_size(dramArbs_3_io_dram_cmd_bits_size),
    .io_dram_cmd_bits_isWr(dramArbs_3_io_dram_cmd_bits_isWr),
    .io_dram_cmd_bits_tag(dramArbs_3_io_dram_cmd_bits_tag),
    .io_dram_wdata_ready(dramArbs_3_io_dram_wdata_ready),
    .io_dram_wdata_valid(dramArbs_3_io_dram_wdata_valid),
    .io_dram_wdata_bits_wdata_0(dramArbs_3_io_dram_wdata_bits_wdata_0),
    .io_dram_wdata_bits_wdata_1(dramArbs_3_io_dram_wdata_bits_wdata_1),
    .io_dram_wdata_bits_wdata_2(dramArbs_3_io_dram_wdata_bits_wdata_2),
    .io_dram_wdata_bits_wdata_3(dramArbs_3_io_dram_wdata_bits_wdata_3),
    .io_dram_wdata_bits_wdata_4(dramArbs_3_io_dram_wdata_bits_wdata_4),
    .io_dram_wdata_bits_wdata_5(dramArbs_3_io_dram_wdata_bits_wdata_5),
    .io_dram_wdata_bits_wdata_6(dramArbs_3_io_dram_wdata_bits_wdata_6),
    .io_dram_wdata_bits_wdata_7(dramArbs_3_io_dram_wdata_bits_wdata_7),
    .io_dram_wdata_bits_wdata_8(dramArbs_3_io_dram_wdata_bits_wdata_8),
    .io_dram_wdata_bits_wdata_9(dramArbs_3_io_dram_wdata_bits_wdata_9),
    .io_dram_wdata_bits_wdata_10(dramArbs_3_io_dram_wdata_bits_wdata_10),
    .io_dram_wdata_bits_wdata_11(dramArbs_3_io_dram_wdata_bits_wdata_11),
    .io_dram_wdata_bits_wdata_12(dramArbs_3_io_dram_wdata_bits_wdata_12),
    .io_dram_wdata_bits_wdata_13(dramArbs_3_io_dram_wdata_bits_wdata_13),
    .io_dram_wdata_bits_wdata_14(dramArbs_3_io_dram_wdata_bits_wdata_14),
    .io_dram_wdata_bits_wdata_15(dramArbs_3_io_dram_wdata_bits_wdata_15),
    .io_dram_wdata_bits_wstrb_0(dramArbs_3_io_dram_wdata_bits_wstrb_0),
    .io_dram_wdata_bits_wstrb_1(dramArbs_3_io_dram_wdata_bits_wstrb_1),
    .io_dram_wdata_bits_wstrb_2(dramArbs_3_io_dram_wdata_bits_wstrb_2),
    .io_dram_wdata_bits_wstrb_3(dramArbs_3_io_dram_wdata_bits_wstrb_3),
    .io_dram_wdata_bits_wstrb_4(dramArbs_3_io_dram_wdata_bits_wstrb_4),
    .io_dram_wdata_bits_wstrb_5(dramArbs_3_io_dram_wdata_bits_wstrb_5),
    .io_dram_wdata_bits_wstrb_6(dramArbs_3_io_dram_wdata_bits_wstrb_6),
    .io_dram_wdata_bits_wstrb_7(dramArbs_3_io_dram_wdata_bits_wstrb_7),
    .io_dram_wdata_bits_wstrb_8(dramArbs_3_io_dram_wdata_bits_wstrb_8),
    .io_dram_wdata_bits_wstrb_9(dramArbs_3_io_dram_wdata_bits_wstrb_9),
    .io_dram_wdata_bits_wstrb_10(dramArbs_3_io_dram_wdata_bits_wstrb_10),
    .io_dram_wdata_bits_wstrb_11(dramArbs_3_io_dram_wdata_bits_wstrb_11),
    .io_dram_wdata_bits_wstrb_12(dramArbs_3_io_dram_wdata_bits_wstrb_12),
    .io_dram_wdata_bits_wstrb_13(dramArbs_3_io_dram_wdata_bits_wstrb_13),
    .io_dram_wdata_bits_wstrb_14(dramArbs_3_io_dram_wdata_bits_wstrb_14),
    .io_dram_wdata_bits_wstrb_15(dramArbs_3_io_dram_wdata_bits_wstrb_15),
    .io_dram_wdata_bits_wstrb_16(dramArbs_3_io_dram_wdata_bits_wstrb_16),
    .io_dram_wdata_bits_wstrb_17(dramArbs_3_io_dram_wdata_bits_wstrb_17),
    .io_dram_wdata_bits_wstrb_18(dramArbs_3_io_dram_wdata_bits_wstrb_18),
    .io_dram_wdata_bits_wstrb_19(dramArbs_3_io_dram_wdata_bits_wstrb_19),
    .io_dram_wdata_bits_wstrb_20(dramArbs_3_io_dram_wdata_bits_wstrb_20),
    .io_dram_wdata_bits_wstrb_21(dramArbs_3_io_dram_wdata_bits_wstrb_21),
    .io_dram_wdata_bits_wstrb_22(dramArbs_3_io_dram_wdata_bits_wstrb_22),
    .io_dram_wdata_bits_wstrb_23(dramArbs_3_io_dram_wdata_bits_wstrb_23),
    .io_dram_wdata_bits_wstrb_24(dramArbs_3_io_dram_wdata_bits_wstrb_24),
    .io_dram_wdata_bits_wstrb_25(dramArbs_3_io_dram_wdata_bits_wstrb_25),
    .io_dram_wdata_bits_wstrb_26(dramArbs_3_io_dram_wdata_bits_wstrb_26),
    .io_dram_wdata_bits_wstrb_27(dramArbs_3_io_dram_wdata_bits_wstrb_27),
    .io_dram_wdata_bits_wstrb_28(dramArbs_3_io_dram_wdata_bits_wstrb_28),
    .io_dram_wdata_bits_wstrb_29(dramArbs_3_io_dram_wdata_bits_wstrb_29),
    .io_dram_wdata_bits_wstrb_30(dramArbs_3_io_dram_wdata_bits_wstrb_30),
    .io_dram_wdata_bits_wstrb_31(dramArbs_3_io_dram_wdata_bits_wstrb_31),
    .io_dram_wdata_bits_wstrb_32(dramArbs_3_io_dram_wdata_bits_wstrb_32),
    .io_dram_wdata_bits_wstrb_33(dramArbs_3_io_dram_wdata_bits_wstrb_33),
    .io_dram_wdata_bits_wstrb_34(dramArbs_3_io_dram_wdata_bits_wstrb_34),
    .io_dram_wdata_bits_wstrb_35(dramArbs_3_io_dram_wdata_bits_wstrb_35),
    .io_dram_wdata_bits_wstrb_36(dramArbs_3_io_dram_wdata_bits_wstrb_36),
    .io_dram_wdata_bits_wstrb_37(dramArbs_3_io_dram_wdata_bits_wstrb_37),
    .io_dram_wdata_bits_wstrb_38(dramArbs_3_io_dram_wdata_bits_wstrb_38),
    .io_dram_wdata_bits_wstrb_39(dramArbs_3_io_dram_wdata_bits_wstrb_39),
    .io_dram_wdata_bits_wstrb_40(dramArbs_3_io_dram_wdata_bits_wstrb_40),
    .io_dram_wdata_bits_wstrb_41(dramArbs_3_io_dram_wdata_bits_wstrb_41),
    .io_dram_wdata_bits_wstrb_42(dramArbs_3_io_dram_wdata_bits_wstrb_42),
    .io_dram_wdata_bits_wstrb_43(dramArbs_3_io_dram_wdata_bits_wstrb_43),
    .io_dram_wdata_bits_wstrb_44(dramArbs_3_io_dram_wdata_bits_wstrb_44),
    .io_dram_wdata_bits_wstrb_45(dramArbs_3_io_dram_wdata_bits_wstrb_45),
    .io_dram_wdata_bits_wstrb_46(dramArbs_3_io_dram_wdata_bits_wstrb_46),
    .io_dram_wdata_bits_wstrb_47(dramArbs_3_io_dram_wdata_bits_wstrb_47),
    .io_dram_wdata_bits_wstrb_48(dramArbs_3_io_dram_wdata_bits_wstrb_48),
    .io_dram_wdata_bits_wstrb_49(dramArbs_3_io_dram_wdata_bits_wstrb_49),
    .io_dram_wdata_bits_wstrb_50(dramArbs_3_io_dram_wdata_bits_wstrb_50),
    .io_dram_wdata_bits_wstrb_51(dramArbs_3_io_dram_wdata_bits_wstrb_51),
    .io_dram_wdata_bits_wstrb_52(dramArbs_3_io_dram_wdata_bits_wstrb_52),
    .io_dram_wdata_bits_wstrb_53(dramArbs_3_io_dram_wdata_bits_wstrb_53),
    .io_dram_wdata_bits_wstrb_54(dramArbs_3_io_dram_wdata_bits_wstrb_54),
    .io_dram_wdata_bits_wstrb_55(dramArbs_3_io_dram_wdata_bits_wstrb_55),
    .io_dram_wdata_bits_wstrb_56(dramArbs_3_io_dram_wdata_bits_wstrb_56),
    .io_dram_wdata_bits_wstrb_57(dramArbs_3_io_dram_wdata_bits_wstrb_57),
    .io_dram_wdata_bits_wstrb_58(dramArbs_3_io_dram_wdata_bits_wstrb_58),
    .io_dram_wdata_bits_wstrb_59(dramArbs_3_io_dram_wdata_bits_wstrb_59),
    .io_dram_wdata_bits_wstrb_60(dramArbs_3_io_dram_wdata_bits_wstrb_60),
    .io_dram_wdata_bits_wstrb_61(dramArbs_3_io_dram_wdata_bits_wstrb_61),
    .io_dram_wdata_bits_wstrb_62(dramArbs_3_io_dram_wdata_bits_wstrb_62),
    .io_dram_wdata_bits_wstrb_63(dramArbs_3_io_dram_wdata_bits_wstrb_63),
    .io_dram_wdata_bits_wlast(dramArbs_3_io_dram_wdata_bits_wlast),
    .io_dram_rresp_ready(dramArbs_3_io_dram_rresp_ready),
    .io_dram_wresp_ready(dramArbs_3_io_dram_wresp_ready),
    .io_dram_wresp_valid(dramArbs_3_io_dram_wresp_valid),
    .io_dram_wresp_bits_tag(dramArbs_3_io_dram_wresp_bits_tag)
  );
  DRAMHeap heap ( // @[Fringe.scala 107:20:@137096.4]
    .io_accel_0_req_valid(heap_io_accel_0_req_valid),
    .io_accel_0_req_bits_allocDealloc(heap_io_accel_0_req_bits_allocDealloc),
    .io_accel_0_req_bits_sizeAddr(heap_io_accel_0_req_bits_sizeAddr),
    .io_accel_0_resp_valid(heap_io_accel_0_resp_valid),
    .io_accel_0_resp_bits_allocDealloc(heap_io_accel_0_resp_bits_allocDealloc),
    .io_accel_0_resp_bits_sizeAddr(heap_io_accel_0_resp_bits_sizeAddr),
    .io_host_0_req_valid(heap_io_host_0_req_valid),
    .io_host_0_req_bits_allocDealloc(heap_io_host_0_req_bits_allocDealloc),
    .io_host_0_req_bits_sizeAddr(heap_io_host_0_req_bits_sizeAddr),
    .io_host_0_resp_valid(heap_io_host_0_resp_valid),
    .io_host_0_resp_bits_allocDealloc(heap_io_host_0_resp_bits_allocDealloc),
    .io_host_0_resp_bits_sizeAddr(heap_io_host_0_resp_bits_sizeAddr)
  );
  RegFile regs ( // @[Fringe.scala 116:20:@137105.4]
    .clock(regs_clock),
    .reset(regs_reset),
    .io_raddr(regs_io_raddr),
    .io_wen(regs_io_wen),
    .io_waddr(regs_io_waddr),
    .io_wdata(regs_io_wdata),
    .io_rdata(regs_io_rdata),
    .io_reset(regs_io_reset),
    .io_argIns_0(regs_io_argIns_0),
    .io_argIns_1(regs_io_argIns_1),
    .io_argIns_2(regs_io_argIns_2),
    .io_argIns_3(regs_io_argIns_3),
    .io_argOuts_0_valid(regs_io_argOuts_0_valid),
    .io_argOuts_0_bits(regs_io_argOuts_0_bits),
    .io_argOuts_1_valid(regs_io_argOuts_1_valid),
    .io_argOuts_1_bits(regs_io_argOuts_1_bits)
  );
  FringeCounter timeoutCtr ( // @[Fringe.scala 143:26:@139155.4]
    .clock(timeoutCtr_clock),
    .reset(timeoutCtr_reset),
    .io_enable(timeoutCtr_io_enable),
    .io_done(timeoutCtr_io_done)
  );
  Depulser depulser ( // @[Fringe.scala 153:24:@139174.4]
    .clock(depulser_clock),
    .reset(depulser_reset),
    .io_in(depulser_io_in),
    .io_rst(depulser_io_rst),
    .io_out(depulser_io_out)
  );
  assign _T_1020 = regs_io_argIns_1; // @[:@139132.4 :@139133.4]
  assign curStatus_done = _T_1020[0]; // @[Fringe.scala 133:45:@139134.4]
  assign curStatus_timeout = _T_1020[1]; // @[Fringe.scala 133:45:@139136.4]
  assign curStatus_allocDealloc = _T_1020[4:2]; // @[Fringe.scala 133:45:@139138.4]
  assign curStatus_sizeAddr = _T_1020[63:5]; // @[Fringe.scala 133:45:@139140.4]
  assign _T_1025 = regs_io_argIns_0[0]; // @[Fringe.scala 134:28:@139142.4]
  assign _T_1029 = curStatus_done == 1'h0; // @[Fringe.scala 134:42:@139144.4]
  assign _T_1030 = regs_io_argIns_0[1]; // @[Fringe.scala 135:27:@139146.4]
  assign _T_1040 = ~ regs_io_argIns_0; // @[Fringe.scala 156:22:@139182.4]
  assign _T_1048 = _T_1047 ^ heap_io_host_0_req_valid; // @[package.scala 153:13:@139187.4]
  assign _T_1049 = heap_io_host_0_req_valid & _T_1048; // @[package.scala 153:8:@139188.4]
  assign _T_1052 = _T_1025 & depulser_io_out; // @[Fringe.scala 160:55:@139192.4]
  assign status_bits_done = depulser_io_out ? _T_1052 : curStatus_done; // @[Fringe.scala 160:26:@139193.4]
  assign _T_1055 = _T_1025 & timeoutCtr_io_done; // @[Fringe.scala 161:58:@139196.4]
  assign status_bits_timeout = depulser_io_out ? _T_1055 : curStatus_timeout; // @[Fringe.scala 161:29:@139197.4]
  assign _T_1059 = heap_io_host_0_req_bits_allocDealloc ? 2'h1 : 2'h2; // @[Fringe.scala 162:57:@139199.4]
  assign _T_1061 = heap_io_host_0_req_valid ? _T_1059 : 2'h0; // @[Fringe.scala 162:34:@139200.4]
  assign _T_1063 = heap_io_host_0_req_valid ? heap_io_host_0_req_bits_sizeAddr : 64'h0; // @[Fringe.scala 163:30:@139202.4]
  assign _T_1064 = {status_bits_timeout,status_bits_done}; // @[Fringe.scala 171:37:@139205.4]
  assign status_bits_sizeAddr = _T_1063[58:0]; // @[Fringe.scala 158:20:@139184.4 Fringe.scala 163:24:@139203.4]
  assign status_bits_allocDealloc = {{1'd0}, _T_1061}; // @[Fringe.scala 158:20:@139184.4 Fringe.scala 162:28:@139201.4]
  assign _T_1065 = {status_bits_sizeAddr,status_bits_allocDealloc}; // @[Fringe.scala 171:37:@139206.4]
  assign alloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 202:38:@140836.4]
  assign dealloc = curStatus_allocDealloc == 3'h4; // @[Fringe.scala 203:40:@140837.4]
  assign _T_1569 = alloc | dealloc; // @[Fringe.scala 204:37:@140838.4]
  assign _T_1573 = _T_1572 ^ _T_1569; // @[package.scala 153:13:@140841.4]
  assign io_rdata = regs_io_rdata; // @[Fringe.scala 125:14:@139130.4]
  assign io_enable = _T_1025 & _T_1029; // @[Fringe.scala 136:13:@139150.4]
  assign io_reset = _T_1030 | reset; // @[Fringe.scala 137:12:@139151.4]
  assign io_argIns_0 = regs_io_argIns_2; // @[Fringe.scala 151:51:@139172.4]
  assign io_argIns_1 = regs_io_argIns_3; // @[Fringe.scala 151:51:@139173.4]
  assign io_memStreams_stores_0_cmd_ready = dramArbs_0_io_app_stores_0_cmd_ready; // @[Fringe.scala 101:72:@134142.4]
  assign io_memStreams_stores_0_data_ready = dramArbs_0_io_app_stores_0_data_ready; // @[Fringe.scala 101:72:@134138.4]
  assign io_memStreams_stores_0_wresp_valid = dramArbs_0_io_app_stores_0_wresp_valid; // @[Fringe.scala 101:72:@134133.4]
  assign io_memStreams_stores_0_wresp_bits = dramArbs_0_io_app_stores_0_wresp_bits; // @[Fringe.scala 101:72:@134132.4]
  assign io_dram_0_cmd_valid = dramArbs_0_io_dram_cmd_valid; // @[Fringe.scala 195:72:@140334.4]
  assign io_dram_0_cmd_bits_addr = dramArbs_0_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@140333.4]
  assign io_dram_0_cmd_bits_size = dramArbs_0_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@140332.4]
  assign io_dram_0_cmd_bits_isWr = dramArbs_0_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@140330.4]
  assign io_dram_0_cmd_bits_tag = dramArbs_0_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@140329.4]
  assign io_dram_0_wdata_valid = dramArbs_0_io_dram_wdata_valid; // @[Fringe.scala 195:72:@140327.4]
  assign io_dram_0_wdata_bits_wdata_0 = dramArbs_0_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@140311.4]
  assign io_dram_0_wdata_bits_wdata_1 = dramArbs_0_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@140312.4]
  assign io_dram_0_wdata_bits_wdata_2 = dramArbs_0_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@140313.4]
  assign io_dram_0_wdata_bits_wdata_3 = dramArbs_0_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@140314.4]
  assign io_dram_0_wdata_bits_wdata_4 = dramArbs_0_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@140315.4]
  assign io_dram_0_wdata_bits_wdata_5 = dramArbs_0_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@140316.4]
  assign io_dram_0_wdata_bits_wdata_6 = dramArbs_0_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@140317.4]
  assign io_dram_0_wdata_bits_wdata_7 = dramArbs_0_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@140318.4]
  assign io_dram_0_wdata_bits_wdata_8 = dramArbs_0_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@140319.4]
  assign io_dram_0_wdata_bits_wdata_9 = dramArbs_0_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@140320.4]
  assign io_dram_0_wdata_bits_wdata_10 = dramArbs_0_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@140321.4]
  assign io_dram_0_wdata_bits_wdata_11 = dramArbs_0_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@140322.4]
  assign io_dram_0_wdata_bits_wdata_12 = dramArbs_0_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@140323.4]
  assign io_dram_0_wdata_bits_wdata_13 = dramArbs_0_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@140324.4]
  assign io_dram_0_wdata_bits_wdata_14 = dramArbs_0_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@140325.4]
  assign io_dram_0_wdata_bits_wdata_15 = dramArbs_0_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@140326.4]
  assign io_dram_0_wdata_bits_wstrb_0 = dramArbs_0_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@140247.4]
  assign io_dram_0_wdata_bits_wstrb_1 = dramArbs_0_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@140248.4]
  assign io_dram_0_wdata_bits_wstrb_2 = dramArbs_0_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@140249.4]
  assign io_dram_0_wdata_bits_wstrb_3 = dramArbs_0_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@140250.4]
  assign io_dram_0_wdata_bits_wstrb_4 = dramArbs_0_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@140251.4]
  assign io_dram_0_wdata_bits_wstrb_5 = dramArbs_0_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@140252.4]
  assign io_dram_0_wdata_bits_wstrb_6 = dramArbs_0_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@140253.4]
  assign io_dram_0_wdata_bits_wstrb_7 = dramArbs_0_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@140254.4]
  assign io_dram_0_wdata_bits_wstrb_8 = dramArbs_0_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@140255.4]
  assign io_dram_0_wdata_bits_wstrb_9 = dramArbs_0_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@140256.4]
  assign io_dram_0_wdata_bits_wstrb_10 = dramArbs_0_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@140257.4]
  assign io_dram_0_wdata_bits_wstrb_11 = dramArbs_0_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@140258.4]
  assign io_dram_0_wdata_bits_wstrb_12 = dramArbs_0_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@140259.4]
  assign io_dram_0_wdata_bits_wstrb_13 = dramArbs_0_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@140260.4]
  assign io_dram_0_wdata_bits_wstrb_14 = dramArbs_0_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@140261.4]
  assign io_dram_0_wdata_bits_wstrb_15 = dramArbs_0_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@140262.4]
  assign io_dram_0_wdata_bits_wstrb_16 = dramArbs_0_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@140263.4]
  assign io_dram_0_wdata_bits_wstrb_17 = dramArbs_0_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@140264.4]
  assign io_dram_0_wdata_bits_wstrb_18 = dramArbs_0_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@140265.4]
  assign io_dram_0_wdata_bits_wstrb_19 = dramArbs_0_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@140266.4]
  assign io_dram_0_wdata_bits_wstrb_20 = dramArbs_0_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@140267.4]
  assign io_dram_0_wdata_bits_wstrb_21 = dramArbs_0_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@140268.4]
  assign io_dram_0_wdata_bits_wstrb_22 = dramArbs_0_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@140269.4]
  assign io_dram_0_wdata_bits_wstrb_23 = dramArbs_0_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@140270.4]
  assign io_dram_0_wdata_bits_wstrb_24 = dramArbs_0_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@140271.4]
  assign io_dram_0_wdata_bits_wstrb_25 = dramArbs_0_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@140272.4]
  assign io_dram_0_wdata_bits_wstrb_26 = dramArbs_0_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@140273.4]
  assign io_dram_0_wdata_bits_wstrb_27 = dramArbs_0_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@140274.4]
  assign io_dram_0_wdata_bits_wstrb_28 = dramArbs_0_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@140275.4]
  assign io_dram_0_wdata_bits_wstrb_29 = dramArbs_0_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@140276.4]
  assign io_dram_0_wdata_bits_wstrb_30 = dramArbs_0_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@140277.4]
  assign io_dram_0_wdata_bits_wstrb_31 = dramArbs_0_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@140278.4]
  assign io_dram_0_wdata_bits_wstrb_32 = dramArbs_0_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@140279.4]
  assign io_dram_0_wdata_bits_wstrb_33 = dramArbs_0_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@140280.4]
  assign io_dram_0_wdata_bits_wstrb_34 = dramArbs_0_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@140281.4]
  assign io_dram_0_wdata_bits_wstrb_35 = dramArbs_0_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@140282.4]
  assign io_dram_0_wdata_bits_wstrb_36 = dramArbs_0_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@140283.4]
  assign io_dram_0_wdata_bits_wstrb_37 = dramArbs_0_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@140284.4]
  assign io_dram_0_wdata_bits_wstrb_38 = dramArbs_0_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@140285.4]
  assign io_dram_0_wdata_bits_wstrb_39 = dramArbs_0_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@140286.4]
  assign io_dram_0_wdata_bits_wstrb_40 = dramArbs_0_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@140287.4]
  assign io_dram_0_wdata_bits_wstrb_41 = dramArbs_0_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@140288.4]
  assign io_dram_0_wdata_bits_wstrb_42 = dramArbs_0_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@140289.4]
  assign io_dram_0_wdata_bits_wstrb_43 = dramArbs_0_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@140290.4]
  assign io_dram_0_wdata_bits_wstrb_44 = dramArbs_0_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@140291.4]
  assign io_dram_0_wdata_bits_wstrb_45 = dramArbs_0_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@140292.4]
  assign io_dram_0_wdata_bits_wstrb_46 = dramArbs_0_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@140293.4]
  assign io_dram_0_wdata_bits_wstrb_47 = dramArbs_0_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@140294.4]
  assign io_dram_0_wdata_bits_wstrb_48 = dramArbs_0_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@140295.4]
  assign io_dram_0_wdata_bits_wstrb_49 = dramArbs_0_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@140296.4]
  assign io_dram_0_wdata_bits_wstrb_50 = dramArbs_0_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@140297.4]
  assign io_dram_0_wdata_bits_wstrb_51 = dramArbs_0_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@140298.4]
  assign io_dram_0_wdata_bits_wstrb_52 = dramArbs_0_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@140299.4]
  assign io_dram_0_wdata_bits_wstrb_53 = dramArbs_0_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@140300.4]
  assign io_dram_0_wdata_bits_wstrb_54 = dramArbs_0_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@140301.4]
  assign io_dram_0_wdata_bits_wstrb_55 = dramArbs_0_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@140302.4]
  assign io_dram_0_wdata_bits_wstrb_56 = dramArbs_0_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@140303.4]
  assign io_dram_0_wdata_bits_wstrb_57 = dramArbs_0_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@140304.4]
  assign io_dram_0_wdata_bits_wstrb_58 = dramArbs_0_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@140305.4]
  assign io_dram_0_wdata_bits_wstrb_59 = dramArbs_0_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@140306.4]
  assign io_dram_0_wdata_bits_wstrb_60 = dramArbs_0_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@140307.4]
  assign io_dram_0_wdata_bits_wstrb_61 = dramArbs_0_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@140308.4]
  assign io_dram_0_wdata_bits_wstrb_62 = dramArbs_0_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@140309.4]
  assign io_dram_0_wdata_bits_wstrb_63 = dramArbs_0_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@140310.4]
  assign io_dram_0_wdata_bits_wlast = dramArbs_0_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@140246.4]
  assign io_dram_0_rresp_ready = dramArbs_0_io_dram_rresp_ready; // @[Fringe.scala 195:72:@140245.4]
  assign io_dram_0_wresp_ready = dramArbs_0_io_dram_wresp_ready; // @[Fringe.scala 195:72:@140226.4]
  assign io_dram_1_cmd_valid = dramArbs_1_io_dram_cmd_valid; // @[Fringe.scala 195:72:@140446.4]
  assign io_dram_1_cmd_bits_addr = dramArbs_1_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@140445.4]
  assign io_dram_1_cmd_bits_size = dramArbs_1_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@140444.4]
  assign io_dram_1_cmd_bits_isWr = dramArbs_1_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@140442.4]
  assign io_dram_1_cmd_bits_tag = dramArbs_1_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@140441.4]
  assign io_dram_1_wdata_valid = dramArbs_1_io_dram_wdata_valid; // @[Fringe.scala 195:72:@140439.4]
  assign io_dram_1_wdata_bits_wdata_0 = dramArbs_1_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@140423.4]
  assign io_dram_1_wdata_bits_wdata_1 = dramArbs_1_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@140424.4]
  assign io_dram_1_wdata_bits_wdata_2 = dramArbs_1_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@140425.4]
  assign io_dram_1_wdata_bits_wdata_3 = dramArbs_1_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@140426.4]
  assign io_dram_1_wdata_bits_wdata_4 = dramArbs_1_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@140427.4]
  assign io_dram_1_wdata_bits_wdata_5 = dramArbs_1_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@140428.4]
  assign io_dram_1_wdata_bits_wdata_6 = dramArbs_1_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@140429.4]
  assign io_dram_1_wdata_bits_wdata_7 = dramArbs_1_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@140430.4]
  assign io_dram_1_wdata_bits_wdata_8 = dramArbs_1_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@140431.4]
  assign io_dram_1_wdata_bits_wdata_9 = dramArbs_1_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@140432.4]
  assign io_dram_1_wdata_bits_wdata_10 = dramArbs_1_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@140433.4]
  assign io_dram_1_wdata_bits_wdata_11 = dramArbs_1_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@140434.4]
  assign io_dram_1_wdata_bits_wdata_12 = dramArbs_1_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@140435.4]
  assign io_dram_1_wdata_bits_wdata_13 = dramArbs_1_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@140436.4]
  assign io_dram_1_wdata_bits_wdata_14 = dramArbs_1_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@140437.4]
  assign io_dram_1_wdata_bits_wdata_15 = dramArbs_1_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@140438.4]
  assign io_dram_1_wdata_bits_wstrb_0 = dramArbs_1_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@140359.4]
  assign io_dram_1_wdata_bits_wstrb_1 = dramArbs_1_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@140360.4]
  assign io_dram_1_wdata_bits_wstrb_2 = dramArbs_1_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@140361.4]
  assign io_dram_1_wdata_bits_wstrb_3 = dramArbs_1_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@140362.4]
  assign io_dram_1_wdata_bits_wstrb_4 = dramArbs_1_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@140363.4]
  assign io_dram_1_wdata_bits_wstrb_5 = dramArbs_1_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@140364.4]
  assign io_dram_1_wdata_bits_wstrb_6 = dramArbs_1_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@140365.4]
  assign io_dram_1_wdata_bits_wstrb_7 = dramArbs_1_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@140366.4]
  assign io_dram_1_wdata_bits_wstrb_8 = dramArbs_1_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@140367.4]
  assign io_dram_1_wdata_bits_wstrb_9 = dramArbs_1_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@140368.4]
  assign io_dram_1_wdata_bits_wstrb_10 = dramArbs_1_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@140369.4]
  assign io_dram_1_wdata_bits_wstrb_11 = dramArbs_1_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@140370.4]
  assign io_dram_1_wdata_bits_wstrb_12 = dramArbs_1_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@140371.4]
  assign io_dram_1_wdata_bits_wstrb_13 = dramArbs_1_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@140372.4]
  assign io_dram_1_wdata_bits_wstrb_14 = dramArbs_1_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@140373.4]
  assign io_dram_1_wdata_bits_wstrb_15 = dramArbs_1_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@140374.4]
  assign io_dram_1_wdata_bits_wstrb_16 = dramArbs_1_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@140375.4]
  assign io_dram_1_wdata_bits_wstrb_17 = dramArbs_1_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@140376.4]
  assign io_dram_1_wdata_bits_wstrb_18 = dramArbs_1_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@140377.4]
  assign io_dram_1_wdata_bits_wstrb_19 = dramArbs_1_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@140378.4]
  assign io_dram_1_wdata_bits_wstrb_20 = dramArbs_1_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@140379.4]
  assign io_dram_1_wdata_bits_wstrb_21 = dramArbs_1_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@140380.4]
  assign io_dram_1_wdata_bits_wstrb_22 = dramArbs_1_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@140381.4]
  assign io_dram_1_wdata_bits_wstrb_23 = dramArbs_1_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@140382.4]
  assign io_dram_1_wdata_bits_wstrb_24 = dramArbs_1_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@140383.4]
  assign io_dram_1_wdata_bits_wstrb_25 = dramArbs_1_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@140384.4]
  assign io_dram_1_wdata_bits_wstrb_26 = dramArbs_1_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@140385.4]
  assign io_dram_1_wdata_bits_wstrb_27 = dramArbs_1_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@140386.4]
  assign io_dram_1_wdata_bits_wstrb_28 = dramArbs_1_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@140387.4]
  assign io_dram_1_wdata_bits_wstrb_29 = dramArbs_1_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@140388.4]
  assign io_dram_1_wdata_bits_wstrb_30 = dramArbs_1_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@140389.4]
  assign io_dram_1_wdata_bits_wstrb_31 = dramArbs_1_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@140390.4]
  assign io_dram_1_wdata_bits_wstrb_32 = dramArbs_1_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@140391.4]
  assign io_dram_1_wdata_bits_wstrb_33 = dramArbs_1_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@140392.4]
  assign io_dram_1_wdata_bits_wstrb_34 = dramArbs_1_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@140393.4]
  assign io_dram_1_wdata_bits_wstrb_35 = dramArbs_1_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@140394.4]
  assign io_dram_1_wdata_bits_wstrb_36 = dramArbs_1_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@140395.4]
  assign io_dram_1_wdata_bits_wstrb_37 = dramArbs_1_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@140396.4]
  assign io_dram_1_wdata_bits_wstrb_38 = dramArbs_1_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@140397.4]
  assign io_dram_1_wdata_bits_wstrb_39 = dramArbs_1_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@140398.4]
  assign io_dram_1_wdata_bits_wstrb_40 = dramArbs_1_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@140399.4]
  assign io_dram_1_wdata_bits_wstrb_41 = dramArbs_1_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@140400.4]
  assign io_dram_1_wdata_bits_wstrb_42 = dramArbs_1_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@140401.4]
  assign io_dram_1_wdata_bits_wstrb_43 = dramArbs_1_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@140402.4]
  assign io_dram_1_wdata_bits_wstrb_44 = dramArbs_1_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@140403.4]
  assign io_dram_1_wdata_bits_wstrb_45 = dramArbs_1_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@140404.4]
  assign io_dram_1_wdata_bits_wstrb_46 = dramArbs_1_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@140405.4]
  assign io_dram_1_wdata_bits_wstrb_47 = dramArbs_1_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@140406.4]
  assign io_dram_1_wdata_bits_wstrb_48 = dramArbs_1_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@140407.4]
  assign io_dram_1_wdata_bits_wstrb_49 = dramArbs_1_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@140408.4]
  assign io_dram_1_wdata_bits_wstrb_50 = dramArbs_1_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@140409.4]
  assign io_dram_1_wdata_bits_wstrb_51 = dramArbs_1_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@140410.4]
  assign io_dram_1_wdata_bits_wstrb_52 = dramArbs_1_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@140411.4]
  assign io_dram_1_wdata_bits_wstrb_53 = dramArbs_1_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@140412.4]
  assign io_dram_1_wdata_bits_wstrb_54 = dramArbs_1_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@140413.4]
  assign io_dram_1_wdata_bits_wstrb_55 = dramArbs_1_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@140414.4]
  assign io_dram_1_wdata_bits_wstrb_56 = dramArbs_1_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@140415.4]
  assign io_dram_1_wdata_bits_wstrb_57 = dramArbs_1_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@140416.4]
  assign io_dram_1_wdata_bits_wstrb_58 = dramArbs_1_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@140417.4]
  assign io_dram_1_wdata_bits_wstrb_59 = dramArbs_1_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@140418.4]
  assign io_dram_1_wdata_bits_wstrb_60 = dramArbs_1_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@140419.4]
  assign io_dram_1_wdata_bits_wstrb_61 = dramArbs_1_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@140420.4]
  assign io_dram_1_wdata_bits_wstrb_62 = dramArbs_1_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@140421.4]
  assign io_dram_1_wdata_bits_wstrb_63 = dramArbs_1_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@140422.4]
  assign io_dram_1_wdata_bits_wlast = dramArbs_1_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@140358.4]
  assign io_dram_1_rresp_ready = dramArbs_1_io_dram_rresp_ready; // @[Fringe.scala 195:72:@140357.4]
  assign io_dram_1_wresp_ready = dramArbs_1_io_dram_wresp_ready; // @[Fringe.scala 195:72:@140338.4]
  assign io_dram_2_cmd_valid = dramArbs_2_io_dram_cmd_valid; // @[Fringe.scala 195:72:@140558.4]
  assign io_dram_2_cmd_bits_addr = dramArbs_2_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@140557.4]
  assign io_dram_2_cmd_bits_size = dramArbs_2_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@140556.4]
  assign io_dram_2_cmd_bits_isWr = dramArbs_2_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@140554.4]
  assign io_dram_2_cmd_bits_tag = dramArbs_2_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@140553.4]
  assign io_dram_2_wdata_valid = dramArbs_2_io_dram_wdata_valid; // @[Fringe.scala 195:72:@140551.4]
  assign io_dram_2_wdata_bits_wdata_0 = dramArbs_2_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@140535.4]
  assign io_dram_2_wdata_bits_wdata_1 = dramArbs_2_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@140536.4]
  assign io_dram_2_wdata_bits_wdata_2 = dramArbs_2_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@140537.4]
  assign io_dram_2_wdata_bits_wdata_3 = dramArbs_2_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@140538.4]
  assign io_dram_2_wdata_bits_wdata_4 = dramArbs_2_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@140539.4]
  assign io_dram_2_wdata_bits_wdata_5 = dramArbs_2_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@140540.4]
  assign io_dram_2_wdata_bits_wdata_6 = dramArbs_2_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@140541.4]
  assign io_dram_2_wdata_bits_wdata_7 = dramArbs_2_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@140542.4]
  assign io_dram_2_wdata_bits_wdata_8 = dramArbs_2_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@140543.4]
  assign io_dram_2_wdata_bits_wdata_9 = dramArbs_2_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@140544.4]
  assign io_dram_2_wdata_bits_wdata_10 = dramArbs_2_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@140545.4]
  assign io_dram_2_wdata_bits_wdata_11 = dramArbs_2_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@140546.4]
  assign io_dram_2_wdata_bits_wdata_12 = dramArbs_2_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@140547.4]
  assign io_dram_2_wdata_bits_wdata_13 = dramArbs_2_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@140548.4]
  assign io_dram_2_wdata_bits_wdata_14 = dramArbs_2_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@140549.4]
  assign io_dram_2_wdata_bits_wdata_15 = dramArbs_2_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@140550.4]
  assign io_dram_2_wdata_bits_wstrb_0 = dramArbs_2_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@140471.4]
  assign io_dram_2_wdata_bits_wstrb_1 = dramArbs_2_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@140472.4]
  assign io_dram_2_wdata_bits_wstrb_2 = dramArbs_2_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@140473.4]
  assign io_dram_2_wdata_bits_wstrb_3 = dramArbs_2_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@140474.4]
  assign io_dram_2_wdata_bits_wstrb_4 = dramArbs_2_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@140475.4]
  assign io_dram_2_wdata_bits_wstrb_5 = dramArbs_2_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@140476.4]
  assign io_dram_2_wdata_bits_wstrb_6 = dramArbs_2_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@140477.4]
  assign io_dram_2_wdata_bits_wstrb_7 = dramArbs_2_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@140478.4]
  assign io_dram_2_wdata_bits_wstrb_8 = dramArbs_2_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@140479.4]
  assign io_dram_2_wdata_bits_wstrb_9 = dramArbs_2_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@140480.4]
  assign io_dram_2_wdata_bits_wstrb_10 = dramArbs_2_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@140481.4]
  assign io_dram_2_wdata_bits_wstrb_11 = dramArbs_2_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@140482.4]
  assign io_dram_2_wdata_bits_wstrb_12 = dramArbs_2_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@140483.4]
  assign io_dram_2_wdata_bits_wstrb_13 = dramArbs_2_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@140484.4]
  assign io_dram_2_wdata_bits_wstrb_14 = dramArbs_2_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@140485.4]
  assign io_dram_2_wdata_bits_wstrb_15 = dramArbs_2_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@140486.4]
  assign io_dram_2_wdata_bits_wstrb_16 = dramArbs_2_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@140487.4]
  assign io_dram_2_wdata_bits_wstrb_17 = dramArbs_2_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@140488.4]
  assign io_dram_2_wdata_bits_wstrb_18 = dramArbs_2_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@140489.4]
  assign io_dram_2_wdata_bits_wstrb_19 = dramArbs_2_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@140490.4]
  assign io_dram_2_wdata_bits_wstrb_20 = dramArbs_2_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@140491.4]
  assign io_dram_2_wdata_bits_wstrb_21 = dramArbs_2_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@140492.4]
  assign io_dram_2_wdata_bits_wstrb_22 = dramArbs_2_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@140493.4]
  assign io_dram_2_wdata_bits_wstrb_23 = dramArbs_2_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@140494.4]
  assign io_dram_2_wdata_bits_wstrb_24 = dramArbs_2_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@140495.4]
  assign io_dram_2_wdata_bits_wstrb_25 = dramArbs_2_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@140496.4]
  assign io_dram_2_wdata_bits_wstrb_26 = dramArbs_2_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@140497.4]
  assign io_dram_2_wdata_bits_wstrb_27 = dramArbs_2_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@140498.4]
  assign io_dram_2_wdata_bits_wstrb_28 = dramArbs_2_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@140499.4]
  assign io_dram_2_wdata_bits_wstrb_29 = dramArbs_2_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@140500.4]
  assign io_dram_2_wdata_bits_wstrb_30 = dramArbs_2_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@140501.4]
  assign io_dram_2_wdata_bits_wstrb_31 = dramArbs_2_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@140502.4]
  assign io_dram_2_wdata_bits_wstrb_32 = dramArbs_2_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@140503.4]
  assign io_dram_2_wdata_bits_wstrb_33 = dramArbs_2_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@140504.4]
  assign io_dram_2_wdata_bits_wstrb_34 = dramArbs_2_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@140505.4]
  assign io_dram_2_wdata_bits_wstrb_35 = dramArbs_2_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@140506.4]
  assign io_dram_2_wdata_bits_wstrb_36 = dramArbs_2_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@140507.4]
  assign io_dram_2_wdata_bits_wstrb_37 = dramArbs_2_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@140508.4]
  assign io_dram_2_wdata_bits_wstrb_38 = dramArbs_2_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@140509.4]
  assign io_dram_2_wdata_bits_wstrb_39 = dramArbs_2_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@140510.4]
  assign io_dram_2_wdata_bits_wstrb_40 = dramArbs_2_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@140511.4]
  assign io_dram_2_wdata_bits_wstrb_41 = dramArbs_2_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@140512.4]
  assign io_dram_2_wdata_bits_wstrb_42 = dramArbs_2_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@140513.4]
  assign io_dram_2_wdata_bits_wstrb_43 = dramArbs_2_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@140514.4]
  assign io_dram_2_wdata_bits_wstrb_44 = dramArbs_2_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@140515.4]
  assign io_dram_2_wdata_bits_wstrb_45 = dramArbs_2_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@140516.4]
  assign io_dram_2_wdata_bits_wstrb_46 = dramArbs_2_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@140517.4]
  assign io_dram_2_wdata_bits_wstrb_47 = dramArbs_2_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@140518.4]
  assign io_dram_2_wdata_bits_wstrb_48 = dramArbs_2_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@140519.4]
  assign io_dram_2_wdata_bits_wstrb_49 = dramArbs_2_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@140520.4]
  assign io_dram_2_wdata_bits_wstrb_50 = dramArbs_2_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@140521.4]
  assign io_dram_2_wdata_bits_wstrb_51 = dramArbs_2_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@140522.4]
  assign io_dram_2_wdata_bits_wstrb_52 = dramArbs_2_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@140523.4]
  assign io_dram_2_wdata_bits_wstrb_53 = dramArbs_2_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@140524.4]
  assign io_dram_2_wdata_bits_wstrb_54 = dramArbs_2_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@140525.4]
  assign io_dram_2_wdata_bits_wstrb_55 = dramArbs_2_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@140526.4]
  assign io_dram_2_wdata_bits_wstrb_56 = dramArbs_2_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@140527.4]
  assign io_dram_2_wdata_bits_wstrb_57 = dramArbs_2_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@140528.4]
  assign io_dram_2_wdata_bits_wstrb_58 = dramArbs_2_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@140529.4]
  assign io_dram_2_wdata_bits_wstrb_59 = dramArbs_2_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@140530.4]
  assign io_dram_2_wdata_bits_wstrb_60 = dramArbs_2_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@140531.4]
  assign io_dram_2_wdata_bits_wstrb_61 = dramArbs_2_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@140532.4]
  assign io_dram_2_wdata_bits_wstrb_62 = dramArbs_2_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@140533.4]
  assign io_dram_2_wdata_bits_wstrb_63 = dramArbs_2_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@140534.4]
  assign io_dram_2_wdata_bits_wlast = dramArbs_2_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@140470.4]
  assign io_dram_2_rresp_ready = dramArbs_2_io_dram_rresp_ready; // @[Fringe.scala 195:72:@140469.4]
  assign io_dram_2_wresp_ready = dramArbs_2_io_dram_wresp_ready; // @[Fringe.scala 195:72:@140450.4]
  assign io_dram_3_cmd_valid = dramArbs_3_io_dram_cmd_valid; // @[Fringe.scala 195:72:@140670.4]
  assign io_dram_3_cmd_bits_addr = dramArbs_3_io_dram_cmd_bits_addr; // @[Fringe.scala 195:72:@140669.4]
  assign io_dram_3_cmd_bits_size = dramArbs_3_io_dram_cmd_bits_size; // @[Fringe.scala 195:72:@140668.4]
  assign io_dram_3_cmd_bits_isWr = dramArbs_3_io_dram_cmd_bits_isWr; // @[Fringe.scala 195:72:@140666.4]
  assign io_dram_3_cmd_bits_tag = dramArbs_3_io_dram_cmd_bits_tag; // @[Fringe.scala 195:72:@140665.4]
  assign io_dram_3_wdata_valid = dramArbs_3_io_dram_wdata_valid; // @[Fringe.scala 195:72:@140663.4]
  assign io_dram_3_wdata_bits_wdata_0 = dramArbs_3_io_dram_wdata_bits_wdata_0; // @[Fringe.scala 195:72:@140647.4]
  assign io_dram_3_wdata_bits_wdata_1 = dramArbs_3_io_dram_wdata_bits_wdata_1; // @[Fringe.scala 195:72:@140648.4]
  assign io_dram_3_wdata_bits_wdata_2 = dramArbs_3_io_dram_wdata_bits_wdata_2; // @[Fringe.scala 195:72:@140649.4]
  assign io_dram_3_wdata_bits_wdata_3 = dramArbs_3_io_dram_wdata_bits_wdata_3; // @[Fringe.scala 195:72:@140650.4]
  assign io_dram_3_wdata_bits_wdata_4 = dramArbs_3_io_dram_wdata_bits_wdata_4; // @[Fringe.scala 195:72:@140651.4]
  assign io_dram_3_wdata_bits_wdata_5 = dramArbs_3_io_dram_wdata_bits_wdata_5; // @[Fringe.scala 195:72:@140652.4]
  assign io_dram_3_wdata_bits_wdata_6 = dramArbs_3_io_dram_wdata_bits_wdata_6; // @[Fringe.scala 195:72:@140653.4]
  assign io_dram_3_wdata_bits_wdata_7 = dramArbs_3_io_dram_wdata_bits_wdata_7; // @[Fringe.scala 195:72:@140654.4]
  assign io_dram_3_wdata_bits_wdata_8 = dramArbs_3_io_dram_wdata_bits_wdata_8; // @[Fringe.scala 195:72:@140655.4]
  assign io_dram_3_wdata_bits_wdata_9 = dramArbs_3_io_dram_wdata_bits_wdata_9; // @[Fringe.scala 195:72:@140656.4]
  assign io_dram_3_wdata_bits_wdata_10 = dramArbs_3_io_dram_wdata_bits_wdata_10; // @[Fringe.scala 195:72:@140657.4]
  assign io_dram_3_wdata_bits_wdata_11 = dramArbs_3_io_dram_wdata_bits_wdata_11; // @[Fringe.scala 195:72:@140658.4]
  assign io_dram_3_wdata_bits_wdata_12 = dramArbs_3_io_dram_wdata_bits_wdata_12; // @[Fringe.scala 195:72:@140659.4]
  assign io_dram_3_wdata_bits_wdata_13 = dramArbs_3_io_dram_wdata_bits_wdata_13; // @[Fringe.scala 195:72:@140660.4]
  assign io_dram_3_wdata_bits_wdata_14 = dramArbs_3_io_dram_wdata_bits_wdata_14; // @[Fringe.scala 195:72:@140661.4]
  assign io_dram_3_wdata_bits_wdata_15 = dramArbs_3_io_dram_wdata_bits_wdata_15; // @[Fringe.scala 195:72:@140662.4]
  assign io_dram_3_wdata_bits_wstrb_0 = dramArbs_3_io_dram_wdata_bits_wstrb_0; // @[Fringe.scala 195:72:@140583.4]
  assign io_dram_3_wdata_bits_wstrb_1 = dramArbs_3_io_dram_wdata_bits_wstrb_1; // @[Fringe.scala 195:72:@140584.4]
  assign io_dram_3_wdata_bits_wstrb_2 = dramArbs_3_io_dram_wdata_bits_wstrb_2; // @[Fringe.scala 195:72:@140585.4]
  assign io_dram_3_wdata_bits_wstrb_3 = dramArbs_3_io_dram_wdata_bits_wstrb_3; // @[Fringe.scala 195:72:@140586.4]
  assign io_dram_3_wdata_bits_wstrb_4 = dramArbs_3_io_dram_wdata_bits_wstrb_4; // @[Fringe.scala 195:72:@140587.4]
  assign io_dram_3_wdata_bits_wstrb_5 = dramArbs_3_io_dram_wdata_bits_wstrb_5; // @[Fringe.scala 195:72:@140588.4]
  assign io_dram_3_wdata_bits_wstrb_6 = dramArbs_3_io_dram_wdata_bits_wstrb_6; // @[Fringe.scala 195:72:@140589.4]
  assign io_dram_3_wdata_bits_wstrb_7 = dramArbs_3_io_dram_wdata_bits_wstrb_7; // @[Fringe.scala 195:72:@140590.4]
  assign io_dram_3_wdata_bits_wstrb_8 = dramArbs_3_io_dram_wdata_bits_wstrb_8; // @[Fringe.scala 195:72:@140591.4]
  assign io_dram_3_wdata_bits_wstrb_9 = dramArbs_3_io_dram_wdata_bits_wstrb_9; // @[Fringe.scala 195:72:@140592.4]
  assign io_dram_3_wdata_bits_wstrb_10 = dramArbs_3_io_dram_wdata_bits_wstrb_10; // @[Fringe.scala 195:72:@140593.4]
  assign io_dram_3_wdata_bits_wstrb_11 = dramArbs_3_io_dram_wdata_bits_wstrb_11; // @[Fringe.scala 195:72:@140594.4]
  assign io_dram_3_wdata_bits_wstrb_12 = dramArbs_3_io_dram_wdata_bits_wstrb_12; // @[Fringe.scala 195:72:@140595.4]
  assign io_dram_3_wdata_bits_wstrb_13 = dramArbs_3_io_dram_wdata_bits_wstrb_13; // @[Fringe.scala 195:72:@140596.4]
  assign io_dram_3_wdata_bits_wstrb_14 = dramArbs_3_io_dram_wdata_bits_wstrb_14; // @[Fringe.scala 195:72:@140597.4]
  assign io_dram_3_wdata_bits_wstrb_15 = dramArbs_3_io_dram_wdata_bits_wstrb_15; // @[Fringe.scala 195:72:@140598.4]
  assign io_dram_3_wdata_bits_wstrb_16 = dramArbs_3_io_dram_wdata_bits_wstrb_16; // @[Fringe.scala 195:72:@140599.4]
  assign io_dram_3_wdata_bits_wstrb_17 = dramArbs_3_io_dram_wdata_bits_wstrb_17; // @[Fringe.scala 195:72:@140600.4]
  assign io_dram_3_wdata_bits_wstrb_18 = dramArbs_3_io_dram_wdata_bits_wstrb_18; // @[Fringe.scala 195:72:@140601.4]
  assign io_dram_3_wdata_bits_wstrb_19 = dramArbs_3_io_dram_wdata_bits_wstrb_19; // @[Fringe.scala 195:72:@140602.4]
  assign io_dram_3_wdata_bits_wstrb_20 = dramArbs_3_io_dram_wdata_bits_wstrb_20; // @[Fringe.scala 195:72:@140603.4]
  assign io_dram_3_wdata_bits_wstrb_21 = dramArbs_3_io_dram_wdata_bits_wstrb_21; // @[Fringe.scala 195:72:@140604.4]
  assign io_dram_3_wdata_bits_wstrb_22 = dramArbs_3_io_dram_wdata_bits_wstrb_22; // @[Fringe.scala 195:72:@140605.4]
  assign io_dram_3_wdata_bits_wstrb_23 = dramArbs_3_io_dram_wdata_bits_wstrb_23; // @[Fringe.scala 195:72:@140606.4]
  assign io_dram_3_wdata_bits_wstrb_24 = dramArbs_3_io_dram_wdata_bits_wstrb_24; // @[Fringe.scala 195:72:@140607.4]
  assign io_dram_3_wdata_bits_wstrb_25 = dramArbs_3_io_dram_wdata_bits_wstrb_25; // @[Fringe.scala 195:72:@140608.4]
  assign io_dram_3_wdata_bits_wstrb_26 = dramArbs_3_io_dram_wdata_bits_wstrb_26; // @[Fringe.scala 195:72:@140609.4]
  assign io_dram_3_wdata_bits_wstrb_27 = dramArbs_3_io_dram_wdata_bits_wstrb_27; // @[Fringe.scala 195:72:@140610.4]
  assign io_dram_3_wdata_bits_wstrb_28 = dramArbs_3_io_dram_wdata_bits_wstrb_28; // @[Fringe.scala 195:72:@140611.4]
  assign io_dram_3_wdata_bits_wstrb_29 = dramArbs_3_io_dram_wdata_bits_wstrb_29; // @[Fringe.scala 195:72:@140612.4]
  assign io_dram_3_wdata_bits_wstrb_30 = dramArbs_3_io_dram_wdata_bits_wstrb_30; // @[Fringe.scala 195:72:@140613.4]
  assign io_dram_3_wdata_bits_wstrb_31 = dramArbs_3_io_dram_wdata_bits_wstrb_31; // @[Fringe.scala 195:72:@140614.4]
  assign io_dram_3_wdata_bits_wstrb_32 = dramArbs_3_io_dram_wdata_bits_wstrb_32; // @[Fringe.scala 195:72:@140615.4]
  assign io_dram_3_wdata_bits_wstrb_33 = dramArbs_3_io_dram_wdata_bits_wstrb_33; // @[Fringe.scala 195:72:@140616.4]
  assign io_dram_3_wdata_bits_wstrb_34 = dramArbs_3_io_dram_wdata_bits_wstrb_34; // @[Fringe.scala 195:72:@140617.4]
  assign io_dram_3_wdata_bits_wstrb_35 = dramArbs_3_io_dram_wdata_bits_wstrb_35; // @[Fringe.scala 195:72:@140618.4]
  assign io_dram_3_wdata_bits_wstrb_36 = dramArbs_3_io_dram_wdata_bits_wstrb_36; // @[Fringe.scala 195:72:@140619.4]
  assign io_dram_3_wdata_bits_wstrb_37 = dramArbs_3_io_dram_wdata_bits_wstrb_37; // @[Fringe.scala 195:72:@140620.4]
  assign io_dram_3_wdata_bits_wstrb_38 = dramArbs_3_io_dram_wdata_bits_wstrb_38; // @[Fringe.scala 195:72:@140621.4]
  assign io_dram_3_wdata_bits_wstrb_39 = dramArbs_3_io_dram_wdata_bits_wstrb_39; // @[Fringe.scala 195:72:@140622.4]
  assign io_dram_3_wdata_bits_wstrb_40 = dramArbs_3_io_dram_wdata_bits_wstrb_40; // @[Fringe.scala 195:72:@140623.4]
  assign io_dram_3_wdata_bits_wstrb_41 = dramArbs_3_io_dram_wdata_bits_wstrb_41; // @[Fringe.scala 195:72:@140624.4]
  assign io_dram_3_wdata_bits_wstrb_42 = dramArbs_3_io_dram_wdata_bits_wstrb_42; // @[Fringe.scala 195:72:@140625.4]
  assign io_dram_3_wdata_bits_wstrb_43 = dramArbs_3_io_dram_wdata_bits_wstrb_43; // @[Fringe.scala 195:72:@140626.4]
  assign io_dram_3_wdata_bits_wstrb_44 = dramArbs_3_io_dram_wdata_bits_wstrb_44; // @[Fringe.scala 195:72:@140627.4]
  assign io_dram_3_wdata_bits_wstrb_45 = dramArbs_3_io_dram_wdata_bits_wstrb_45; // @[Fringe.scala 195:72:@140628.4]
  assign io_dram_3_wdata_bits_wstrb_46 = dramArbs_3_io_dram_wdata_bits_wstrb_46; // @[Fringe.scala 195:72:@140629.4]
  assign io_dram_3_wdata_bits_wstrb_47 = dramArbs_3_io_dram_wdata_bits_wstrb_47; // @[Fringe.scala 195:72:@140630.4]
  assign io_dram_3_wdata_bits_wstrb_48 = dramArbs_3_io_dram_wdata_bits_wstrb_48; // @[Fringe.scala 195:72:@140631.4]
  assign io_dram_3_wdata_bits_wstrb_49 = dramArbs_3_io_dram_wdata_bits_wstrb_49; // @[Fringe.scala 195:72:@140632.4]
  assign io_dram_3_wdata_bits_wstrb_50 = dramArbs_3_io_dram_wdata_bits_wstrb_50; // @[Fringe.scala 195:72:@140633.4]
  assign io_dram_3_wdata_bits_wstrb_51 = dramArbs_3_io_dram_wdata_bits_wstrb_51; // @[Fringe.scala 195:72:@140634.4]
  assign io_dram_3_wdata_bits_wstrb_52 = dramArbs_3_io_dram_wdata_bits_wstrb_52; // @[Fringe.scala 195:72:@140635.4]
  assign io_dram_3_wdata_bits_wstrb_53 = dramArbs_3_io_dram_wdata_bits_wstrb_53; // @[Fringe.scala 195:72:@140636.4]
  assign io_dram_3_wdata_bits_wstrb_54 = dramArbs_3_io_dram_wdata_bits_wstrb_54; // @[Fringe.scala 195:72:@140637.4]
  assign io_dram_3_wdata_bits_wstrb_55 = dramArbs_3_io_dram_wdata_bits_wstrb_55; // @[Fringe.scala 195:72:@140638.4]
  assign io_dram_3_wdata_bits_wstrb_56 = dramArbs_3_io_dram_wdata_bits_wstrb_56; // @[Fringe.scala 195:72:@140639.4]
  assign io_dram_3_wdata_bits_wstrb_57 = dramArbs_3_io_dram_wdata_bits_wstrb_57; // @[Fringe.scala 195:72:@140640.4]
  assign io_dram_3_wdata_bits_wstrb_58 = dramArbs_3_io_dram_wdata_bits_wstrb_58; // @[Fringe.scala 195:72:@140641.4]
  assign io_dram_3_wdata_bits_wstrb_59 = dramArbs_3_io_dram_wdata_bits_wstrb_59; // @[Fringe.scala 195:72:@140642.4]
  assign io_dram_3_wdata_bits_wstrb_60 = dramArbs_3_io_dram_wdata_bits_wstrb_60; // @[Fringe.scala 195:72:@140643.4]
  assign io_dram_3_wdata_bits_wstrb_61 = dramArbs_3_io_dram_wdata_bits_wstrb_61; // @[Fringe.scala 195:72:@140644.4]
  assign io_dram_3_wdata_bits_wstrb_62 = dramArbs_3_io_dram_wdata_bits_wstrb_62; // @[Fringe.scala 195:72:@140645.4]
  assign io_dram_3_wdata_bits_wstrb_63 = dramArbs_3_io_dram_wdata_bits_wstrb_63; // @[Fringe.scala 195:72:@140646.4]
  assign io_dram_3_wdata_bits_wlast = dramArbs_3_io_dram_wdata_bits_wlast; // @[Fringe.scala 195:72:@140582.4]
  assign io_dram_3_rresp_ready = dramArbs_3_io_dram_rresp_ready; // @[Fringe.scala 195:72:@140581.4]
  assign io_dram_3_wresp_ready = dramArbs_3_io_dram_wresp_ready; // @[Fringe.scala 195:72:@140562.4]
  assign io_heap_0_resp_valid = heap_io_accel_0_resp_valid; // @[Fringe.scala 108:17:@137101.4]
  assign io_heap_0_resp_bits_allocDealloc = heap_io_accel_0_resp_bits_allocDealloc; // @[Fringe.scala 108:17:@137100.4]
  assign io_heap_0_resp_bits_sizeAddr = heap_io_accel_0_resp_bits_sizeAddr; // @[Fringe.scala 108:17:@137099.4]
  assign dramArbs_0_clock = clock; // @[:@133224.4]
  assign dramArbs_0_reset = _T_1030 | reset; // @[:@133225.4 Fringe.scala 187:30:@140216.4]
  assign dramArbs_0_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@140220.4]
  assign dramArbs_0_io_app_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[Fringe.scala 101:72:@134141.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[Fringe.scala 101:72:@134140.4]
  assign dramArbs_0_io_app_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[Fringe.scala 101:72:@134139.4]
  assign dramArbs_0_io_app_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[Fringe.scala 101:72:@134137.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[Fringe.scala 101:72:@134136.4]
  assign dramArbs_0_io_app_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[Fringe.scala 101:72:@134135.4]
  assign dramArbs_0_io_app_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[Fringe.scala 101:72:@134134.4]
  assign dramArbs_0_io_dram_cmd_ready = io_dram_0_cmd_ready; // @[Fringe.scala 195:72:@140335.4]
  assign dramArbs_0_io_dram_wdata_ready = io_dram_0_wdata_ready; // @[Fringe.scala 195:72:@140328.4]
  assign dramArbs_0_io_dram_wresp_valid = io_dram_0_wresp_valid; // @[Fringe.scala 195:72:@140225.4]
  assign dramArbs_0_io_dram_wresp_bits_tag = io_dram_0_wresp_bits_tag; // @[Fringe.scala 195:72:@140224.4]
  assign dramArbs_1_clock = clock; // @[:@134217.4]
  assign dramArbs_1_reset = _T_1030 | reset; // @[:@134218.4 Fringe.scala 187:30:@140217.4]
  assign dramArbs_1_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@140221.4]
  assign dramArbs_1_io_dram_cmd_ready = io_dram_1_cmd_ready; // @[Fringe.scala 195:72:@140447.4]
  assign dramArbs_1_io_dram_wdata_ready = io_dram_1_wdata_ready; // @[Fringe.scala 195:72:@140440.4]
  assign dramArbs_1_io_dram_wresp_valid = io_dram_1_wresp_valid; // @[Fringe.scala 195:72:@140337.4]
  assign dramArbs_1_io_dram_wresp_bits_tag = io_dram_1_wresp_bits_tag; // @[Fringe.scala 195:72:@140336.4]
  assign dramArbs_2_clock = clock; // @[:@135177.4]
  assign dramArbs_2_reset = _T_1030 | reset; // @[:@135178.4 Fringe.scala 187:30:@140218.4]
  assign dramArbs_2_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@140222.4]
  assign dramArbs_2_io_dram_cmd_ready = io_dram_2_cmd_ready; // @[Fringe.scala 195:72:@140559.4]
  assign dramArbs_2_io_dram_wdata_ready = io_dram_2_wdata_ready; // @[Fringe.scala 195:72:@140552.4]
  assign dramArbs_2_io_dram_wresp_valid = io_dram_2_wresp_valid; // @[Fringe.scala 195:72:@140449.4]
  assign dramArbs_2_io_dram_wresp_bits_tag = io_dram_2_wresp_bits_tag; // @[Fringe.scala 195:72:@140448.4]
  assign dramArbs_3_clock = clock; // @[:@136137.4]
  assign dramArbs_3_reset = _T_1030 | reset; // @[:@136138.4 Fringe.scala 187:30:@140219.4]
  assign dramArbs_3_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 192:36:@140223.4]
  assign dramArbs_3_io_dram_cmd_ready = io_dram_3_cmd_ready; // @[Fringe.scala 195:72:@140671.4]
  assign dramArbs_3_io_dram_wdata_ready = io_dram_3_wdata_ready; // @[Fringe.scala 195:72:@140664.4]
  assign dramArbs_3_io_dram_wresp_valid = io_dram_3_wresp_valid; // @[Fringe.scala 195:72:@140561.4]
  assign dramArbs_3_io_dram_wresp_bits_tag = io_dram_3_wresp_bits_tag; // @[Fringe.scala 195:72:@140560.4]
  assign heap_io_accel_0_req_valid = io_heap_0_req_valid; // @[Fringe.scala 108:17:@137104.4]
  assign heap_io_accel_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[Fringe.scala 108:17:@137103.4]
  assign heap_io_accel_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[Fringe.scala 108:17:@137102.4]
  assign heap_io_host_0_resp_valid = _T_1569 & _T_1573; // @[Fringe.scala 204:22:@140843.4]
  assign heap_io_host_0_resp_bits_allocDealloc = curStatus_allocDealloc == 3'h3; // @[Fringe.scala 205:34:@140844.4]
  assign heap_io_host_0_resp_bits_sizeAddr = {{5'd0}, curStatus_sizeAddr}; // @[Fringe.scala 206:30:@140845.4]
  assign regs_clock = clock; // @[:@137106.4]
  assign regs_reset = reset; // @[:@137107.4 Fringe.scala 139:14:@139154.4]
  assign regs_io_raddr = io_raddr; // @[Fringe.scala 118:17:@139126.4]
  assign regs_io_wen = io_wen; // @[Fringe.scala 120:15:@139128.4]
  assign regs_io_waddr = io_waddr; // @[Fringe.scala 119:17:@139127.4]
  assign regs_io_wdata = io_wdata; // @[Fringe.scala 121:17:@139129.4]
  assign regs_io_reset = _T_1030 | reset; // @[Fringe.scala 138:17:@139152.4]
  assign regs_io_argOuts_0_valid = depulser_io_out | _T_1049; // @[Fringe.scala 170:23:@139204.4]
  assign regs_io_argOuts_0_bits = {_T_1065,_T_1064}; // @[Fringe.scala 171:22:@139208.4]
  assign regs_io_argOuts_1_valid = io_argOuts_0_valid; // @[Fringe.scala 176:23:@139211.4]
  assign regs_io_argOuts_1_bits = io_argOuts_0_bits; // @[Fringe.scala 175:22:@139210.4]
  assign timeoutCtr_clock = clock; // @[:@139156.4]
  assign timeoutCtr_reset = reset; // @[:@139157.4]
  assign timeoutCtr_io_enable = _T_1025 & _T_1029; // @[Fringe.scala 149:24:@139171.4]
  assign depulser_clock = clock; // @[:@139175.4]
  assign depulser_reset = reset; // @[:@139176.4]
  assign depulser_io_in = io_done | timeoutCtr_io_done; // @[Fringe.scala 155:18:@139181.4]
  assign depulser_io_rst = _T_1040[0]; // @[Fringe.scala 156:19:@139183.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1047 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_1572 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_1047 <= 1'h0;
    end else begin
      _T_1047 <= heap_io_host_0_req_valid;
    end
    if (reset) begin
      _T_1572 <= 1'h0;
    end else begin
      _T_1572 <= _T_1569;
    end
  end
endmodule
module AXI4LiteToRFBridge( // @[:@140860.2]
  input         clock, // @[:@140861.4]
  input         reset, // @[:@140862.4]
  input  [31:0] io_S_AXI_AWADDR, // @[:@140863.4]
  input  [2:0]  io_S_AXI_AWPROT, // @[:@140863.4]
  input         io_S_AXI_AWVALID, // @[:@140863.4]
  output        io_S_AXI_AWREADY, // @[:@140863.4]
  input  [31:0] io_S_AXI_ARADDR, // @[:@140863.4]
  input  [2:0]  io_S_AXI_ARPROT, // @[:@140863.4]
  input         io_S_AXI_ARVALID, // @[:@140863.4]
  output        io_S_AXI_ARREADY, // @[:@140863.4]
  input  [31:0] io_S_AXI_WDATA, // @[:@140863.4]
  input  [3:0]  io_S_AXI_WSTRB, // @[:@140863.4]
  input         io_S_AXI_WVALID, // @[:@140863.4]
  output        io_S_AXI_WREADY, // @[:@140863.4]
  output [31:0] io_S_AXI_RDATA, // @[:@140863.4]
  output [1:0]  io_S_AXI_RRESP, // @[:@140863.4]
  output        io_S_AXI_RVALID, // @[:@140863.4]
  input         io_S_AXI_RREADY, // @[:@140863.4]
  output [1:0]  io_S_AXI_BRESP, // @[:@140863.4]
  output        io_S_AXI_BVALID, // @[:@140863.4]
  input         io_S_AXI_BREADY, // @[:@140863.4]
  output [31:0] io_raddr, // @[:@140863.4]
  output        io_wen, // @[:@140863.4]
  output [31:0] io_waddr, // @[:@140863.4]
  output [31:0] io_wdata, // @[:@140863.4]
  input  [31:0] io_rdata // @[:@140863.4]
);
  wire [31:0] d_rf_rdata; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [31:0] d_rf_wdata; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [31:0] d_rf_waddr; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_rf_wen; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [31:0] d_rf_raddr; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_ARESETN; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_ACLK; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [31:0] d_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [2:0] d_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [31:0] d_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [2:0] d_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [31:0] d_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [3:0] d_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [31:0] d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [1:0] d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire [1:0] d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  wire  d_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
  AXI4LiteToRFBridgeVerilog d ( // @[AXI4LiteToRFBridge.scala 36:17:@140865.4]
    .rf_rdata(d_rf_rdata),
    .rf_wdata(d_rf_wdata),
    .rf_waddr(d_rf_waddr),
    .rf_wen(d_rf_wen),
    .rf_raddr(d_rf_raddr),
    .S_AXI_ARESETN(d_S_AXI_ARESETN),
    .S_AXI_ACLK(d_S_AXI_ACLK),
    .S_AXI_AWADDR(d_S_AXI_AWADDR),
    .S_AXI_AWPROT(d_S_AXI_AWPROT),
    .S_AXI_AWVALID(d_S_AXI_AWVALID),
    .S_AXI_AWREADY(d_S_AXI_AWREADY),
    .S_AXI_ARADDR(d_S_AXI_ARADDR),
    .S_AXI_ARPROT(d_S_AXI_ARPROT),
    .S_AXI_ARVALID(d_S_AXI_ARVALID),
    .S_AXI_ARREADY(d_S_AXI_ARREADY),
    .S_AXI_WDATA(d_S_AXI_WDATA),
    .S_AXI_WSTRB(d_S_AXI_WSTRB),
    .S_AXI_WVALID(d_S_AXI_WVALID),
    .S_AXI_WREADY(d_S_AXI_WREADY),
    .S_AXI_RDATA(d_S_AXI_RDATA),
    .S_AXI_RRESP(d_S_AXI_RRESP),
    .S_AXI_RVALID(d_S_AXI_RVALID),
    .S_AXI_RREADY(d_S_AXI_RREADY),
    .S_AXI_BRESP(d_S_AXI_BRESP),
    .S_AXI_BVALID(d_S_AXI_BVALID),
    .S_AXI_BREADY(d_S_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = d_S_AXI_AWREADY; // @[AXI4LiteToRFBridge.scala 38:14:@140889.4]
  assign io_S_AXI_ARREADY = d_S_AXI_ARREADY; // @[AXI4LiteToRFBridge.scala 38:14:@140885.4]
  assign io_S_AXI_WREADY = d_S_AXI_WREADY; // @[AXI4LiteToRFBridge.scala 38:14:@140881.4]
  assign io_S_AXI_RDATA = d_S_AXI_RDATA; // @[AXI4LiteToRFBridge.scala 38:14:@140880.4]
  assign io_S_AXI_RRESP = d_S_AXI_RRESP; // @[AXI4LiteToRFBridge.scala 38:14:@140879.4]
  assign io_S_AXI_RVALID = d_S_AXI_RVALID; // @[AXI4LiteToRFBridge.scala 38:14:@140878.4]
  assign io_S_AXI_BRESP = d_S_AXI_BRESP; // @[AXI4LiteToRFBridge.scala 38:14:@140876.4]
  assign io_S_AXI_BVALID = d_S_AXI_BVALID; // @[AXI4LiteToRFBridge.scala 38:14:@140875.4]
  assign io_raddr = d_rf_raddr; // @[AXI4LiteToRFBridge.scala 42:12:@140897.4]
  assign io_wen = d_rf_wen; // @[AXI4LiteToRFBridge.scala 45:12:@140900.4]
  assign io_waddr = d_rf_waddr; // @[AXI4LiteToRFBridge.scala 43:12:@140898.4]
  assign io_wdata = d_rf_wdata; // @[AXI4LiteToRFBridge.scala 44:12:@140899.4]
  assign d_rf_rdata = io_rdata; // @[AXI4LiteToRFBridge.scala 46:17:@140901.4]
  assign d_S_AXI_ARESETN = ~ reset; // @[AXI4LiteToRFBridge.scala 40:22:@140896.4]
  assign d_S_AXI_ACLK = clock; // @[AXI4LiteToRFBridge.scala 39:19:@140893.4]
  assign d_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[AXI4LiteToRFBridge.scala 38:14:@140892.4]
  assign d_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[AXI4LiteToRFBridge.scala 38:14:@140891.4]
  assign d_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[AXI4LiteToRFBridge.scala 38:14:@140890.4]
  assign d_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[AXI4LiteToRFBridge.scala 38:14:@140888.4]
  assign d_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[AXI4LiteToRFBridge.scala 38:14:@140887.4]
  assign d_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[AXI4LiteToRFBridge.scala 38:14:@140886.4]
  assign d_S_AXI_WDATA = io_S_AXI_WDATA; // @[AXI4LiteToRFBridge.scala 38:14:@140884.4]
  assign d_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[AXI4LiteToRFBridge.scala 38:14:@140883.4]
  assign d_S_AXI_WVALID = io_S_AXI_WVALID; // @[AXI4LiteToRFBridge.scala 38:14:@140882.4]
  assign d_S_AXI_RREADY = io_S_AXI_RREADY; // @[AXI4LiteToRFBridge.scala 38:14:@140877.4]
  assign d_S_AXI_BREADY = io_S_AXI_BREADY; // @[AXI4LiteToRFBridge.scala 38:14:@140874.4]
endmodule
module MAGToAXI4Bridge( // @[:@140903.2]
  output         io_in_cmd_ready, // @[:@140906.4]
  input          io_in_cmd_valid, // @[:@140906.4]
  input  [63:0]  io_in_cmd_bits_addr, // @[:@140906.4]
  input  [31:0]  io_in_cmd_bits_size, // @[:@140906.4]
  input          io_in_cmd_bits_isWr, // @[:@140906.4]
  input  [31:0]  io_in_cmd_bits_tag, // @[:@140906.4]
  output         io_in_wdata_ready, // @[:@140906.4]
  input          io_in_wdata_valid, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_0, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_1, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_2, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_3, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_4, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_5, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_6, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_7, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_8, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_9, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_10, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_11, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_12, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_13, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_14, // @[:@140906.4]
  input  [31:0]  io_in_wdata_bits_wdata_15, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_0, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_1, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_2, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_3, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_4, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_5, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_6, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_7, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_8, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_9, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_10, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_11, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_12, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_13, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_14, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_15, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_16, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_17, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_18, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_19, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_20, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_21, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_22, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_23, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_24, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_25, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_26, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_27, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_28, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_29, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_30, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_31, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_32, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_33, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_34, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_35, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_36, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_37, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_38, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_39, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_40, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_41, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_42, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_43, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_44, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_45, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_46, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_47, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_48, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_49, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_50, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_51, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_52, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_53, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_54, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_55, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_56, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_57, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_58, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_59, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_60, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_61, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_62, // @[:@140906.4]
  input          io_in_wdata_bits_wstrb_63, // @[:@140906.4]
  input          io_in_wdata_bits_wlast, // @[:@140906.4]
  input          io_in_rresp_ready, // @[:@140906.4]
  input          io_in_wresp_ready, // @[:@140906.4]
  output         io_in_wresp_valid, // @[:@140906.4]
  output [31:0]  io_in_wresp_bits_tag, // @[:@140906.4]
  output [31:0]  io_M_AXI_AWID, // @[:@140906.4]
  output [31:0]  io_M_AXI_AWADDR, // @[:@140906.4]
  output [7:0]   io_M_AXI_AWLEN, // @[:@140906.4]
  output         io_M_AXI_AWVALID, // @[:@140906.4]
  input          io_M_AXI_AWREADY, // @[:@140906.4]
  output [31:0]  io_M_AXI_ARID, // @[:@140906.4]
  output [31:0]  io_M_AXI_ARADDR, // @[:@140906.4]
  output [7:0]   io_M_AXI_ARLEN, // @[:@140906.4]
  output         io_M_AXI_ARVALID, // @[:@140906.4]
  input          io_M_AXI_ARREADY, // @[:@140906.4]
  output [511:0] io_M_AXI_WDATA, // @[:@140906.4]
  output [63:0]  io_M_AXI_WSTRB, // @[:@140906.4]
  output         io_M_AXI_WLAST, // @[:@140906.4]
  output         io_M_AXI_WVALID, // @[:@140906.4]
  input          io_M_AXI_WREADY, // @[:@140906.4]
  output         io_M_AXI_RREADY, // @[:@140906.4]
  input  [31:0]  io_M_AXI_BID, // @[:@140906.4]
  input          io_M_AXI_BVALID, // @[:@140906.4]
  output         io_M_AXI_BREADY // @[:@140906.4]
);
  wire [32:0] _T_218; // @[MAGToAXI4Bridge.scala 27:29:@141063.4]
  wire [32:0] _T_219; // @[MAGToAXI4Bridge.scala 27:29:@141064.4]
  wire [31:0] _T_220; // @[MAGToAXI4Bridge.scala 27:29:@141065.4]
  wire  _T_228; // @[MAGToAXI4Bridge.scala 35:42:@141073.4]
  wire [319:0] _T_250; // @[Cat.scala 30:58:@141100.4]
  wire [479:0] _T_255; // @[Cat.scala 30:58:@141105.4]
  wire [9:0] _T_265; // @[Cat.scala 30:58:@141116.4]
  wire [18:0] _T_274; // @[Cat.scala 30:58:@141125.4]
  wire [27:0] _T_283; // @[Cat.scala 30:58:@141134.4]
  wire [36:0] _T_292; // @[Cat.scala 30:58:@141143.4]
  wire [45:0] _T_301; // @[Cat.scala 30:58:@141152.4]
  wire [54:0] _T_310; // @[Cat.scala 30:58:@141161.4]
  wire [62:0] _T_318; // @[Cat.scala 30:58:@141169.4]
  assign _T_218 = io_in_cmd_bits_size - 32'h1; // @[MAGToAXI4Bridge.scala 27:29:@141063.4]
  assign _T_219 = $unsigned(_T_218); // @[MAGToAXI4Bridge.scala 27:29:@141064.4]
  assign _T_220 = _T_219[31:0]; // @[MAGToAXI4Bridge.scala 27:29:@141065.4]
  assign _T_228 = io_in_cmd_bits_isWr == 1'h0; // @[MAGToAXI4Bridge.scala 35:42:@141073.4]
  assign _T_250 = {io_in_wdata_bits_wdata_15,io_in_wdata_bits_wdata_14,io_in_wdata_bits_wdata_13,io_in_wdata_bits_wdata_12,io_in_wdata_bits_wdata_11,io_in_wdata_bits_wdata_10,io_in_wdata_bits_wdata_9,io_in_wdata_bits_wdata_8,io_in_wdata_bits_wdata_7,io_in_wdata_bits_wdata_6}; // @[Cat.scala 30:58:@141100.4]
  assign _T_255 = {_T_250,io_in_wdata_bits_wdata_5,io_in_wdata_bits_wdata_4,io_in_wdata_bits_wdata_3,io_in_wdata_bits_wdata_2,io_in_wdata_bits_wdata_1}; // @[Cat.scala 30:58:@141105.4]
  assign _T_265 = {io_in_wdata_bits_wstrb_63,io_in_wdata_bits_wstrb_62,io_in_wdata_bits_wstrb_61,io_in_wdata_bits_wstrb_60,io_in_wdata_bits_wstrb_59,io_in_wdata_bits_wstrb_58,io_in_wdata_bits_wstrb_57,io_in_wdata_bits_wstrb_56,io_in_wdata_bits_wstrb_55,io_in_wdata_bits_wstrb_54}; // @[Cat.scala 30:58:@141116.4]
  assign _T_274 = {_T_265,io_in_wdata_bits_wstrb_53,io_in_wdata_bits_wstrb_52,io_in_wdata_bits_wstrb_51,io_in_wdata_bits_wstrb_50,io_in_wdata_bits_wstrb_49,io_in_wdata_bits_wstrb_48,io_in_wdata_bits_wstrb_47,io_in_wdata_bits_wstrb_46,io_in_wdata_bits_wstrb_45}; // @[Cat.scala 30:58:@141125.4]
  assign _T_283 = {_T_274,io_in_wdata_bits_wstrb_44,io_in_wdata_bits_wstrb_43,io_in_wdata_bits_wstrb_42,io_in_wdata_bits_wstrb_41,io_in_wdata_bits_wstrb_40,io_in_wdata_bits_wstrb_39,io_in_wdata_bits_wstrb_38,io_in_wdata_bits_wstrb_37,io_in_wdata_bits_wstrb_36}; // @[Cat.scala 30:58:@141134.4]
  assign _T_292 = {_T_283,io_in_wdata_bits_wstrb_35,io_in_wdata_bits_wstrb_34,io_in_wdata_bits_wstrb_33,io_in_wdata_bits_wstrb_32,io_in_wdata_bits_wstrb_31,io_in_wdata_bits_wstrb_30,io_in_wdata_bits_wstrb_29,io_in_wdata_bits_wstrb_28,io_in_wdata_bits_wstrb_27}; // @[Cat.scala 30:58:@141143.4]
  assign _T_301 = {_T_292,io_in_wdata_bits_wstrb_26,io_in_wdata_bits_wstrb_25,io_in_wdata_bits_wstrb_24,io_in_wdata_bits_wstrb_23,io_in_wdata_bits_wstrb_22,io_in_wdata_bits_wstrb_21,io_in_wdata_bits_wstrb_20,io_in_wdata_bits_wstrb_19,io_in_wdata_bits_wstrb_18}; // @[Cat.scala 30:58:@141152.4]
  assign _T_310 = {_T_301,io_in_wdata_bits_wstrb_17,io_in_wdata_bits_wstrb_16,io_in_wdata_bits_wstrb_15,io_in_wdata_bits_wstrb_14,io_in_wdata_bits_wstrb_13,io_in_wdata_bits_wstrb_12,io_in_wdata_bits_wstrb_11,io_in_wdata_bits_wstrb_10,io_in_wdata_bits_wstrb_9}; // @[Cat.scala 30:58:@141161.4]
  assign _T_318 = {_T_310,io_in_wdata_bits_wstrb_8,io_in_wdata_bits_wstrb_7,io_in_wdata_bits_wstrb_6,io_in_wdata_bits_wstrb_5,io_in_wdata_bits_wstrb_4,io_in_wdata_bits_wstrb_3,io_in_wdata_bits_wstrb_2,io_in_wdata_bits_wstrb_1}; // @[Cat.scala 30:58:@141169.4]
  assign io_in_cmd_ready = io_in_cmd_bits_isWr ? io_M_AXI_AWREADY : io_M_AXI_ARREADY; // @[MAGToAXI4Bridge.scala 36:21:@141077.4]
  assign io_in_wdata_ready = io_M_AXI_WREADY; // @[MAGToAXI4Bridge.scala 56:21:@141174.4]
  assign io_in_wresp_valid = io_M_AXI_BVALID; // @[MAGToAXI4Bridge.scala 71:21:@141227.4]
  assign io_in_wresp_bits_tag = io_M_AXI_BID; // @[MAGToAXI4Bridge.scala 74:24:@141229.4]
  assign io_M_AXI_AWID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 39:21:@141078.4]
  assign io_M_AXI_AWADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 40:21:@141079.4]
  assign io_M_AXI_AWLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 41:21:@141083.4]
  assign io_M_AXI_AWVALID = io_in_cmd_valid & io_in_cmd_bits_isWr; // @[MAGToAXI4Bridge.scala 49:21:@141091.4]
  assign io_M_AXI_ARID = io_in_cmd_bits_tag; // @[MAGToAXI4Bridge.scala 25:21:@141061.4]
  assign io_M_AXI_ARADDR = io_in_cmd_bits_addr[31:0]; // @[MAGToAXI4Bridge.scala 26:21:@141062.4]
  assign io_M_AXI_ARLEN = _T_220[7:0]; // @[MAGToAXI4Bridge.scala 27:21:@141066.4]
  assign io_M_AXI_ARVALID = io_in_cmd_valid & _T_228; // @[MAGToAXI4Bridge.scala 35:21:@141075.4]
  assign io_M_AXI_WDATA = {_T_255,io_in_wdata_bits_wdata_0}; // @[MAGToAXI4Bridge.scala 52:21:@141107.4]
  assign io_M_AXI_WSTRB = {_T_318,io_in_wdata_bits_wstrb_0}; // @[MAGToAXI4Bridge.scala 53:21:@141171.4]
  assign io_M_AXI_WLAST = io_in_wdata_bits_wlast; // @[MAGToAXI4Bridge.scala 54:21:@141172.4]
  assign io_M_AXI_WVALID = io_in_wdata_valid; // @[MAGToAXI4Bridge.scala 55:21:@141173.4]
  assign io_M_AXI_RREADY = io_in_rresp_ready; // @[MAGToAXI4Bridge.scala 64:19:@141224.4]
  assign io_M_AXI_BREADY = io_in_wresp_ready; // @[MAGToAXI4Bridge.scala 67:19:@141225.4]
endmodule
module FringeZynq( // @[:@142215.2]
  input          clock, // @[:@142216.4]
  input          reset, // @[:@142217.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@142218.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@142218.4]
  input          io_S_AXI_AWVALID, // @[:@142218.4]
  output         io_S_AXI_AWREADY, // @[:@142218.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@142218.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@142218.4]
  input          io_S_AXI_ARVALID, // @[:@142218.4]
  output         io_S_AXI_ARREADY, // @[:@142218.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@142218.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@142218.4]
  input          io_S_AXI_WVALID, // @[:@142218.4]
  output         io_S_AXI_WREADY, // @[:@142218.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@142218.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@142218.4]
  output         io_S_AXI_RVALID, // @[:@142218.4]
  input          io_S_AXI_RREADY, // @[:@142218.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@142218.4]
  output         io_S_AXI_BVALID, // @[:@142218.4]
  input          io_S_AXI_BREADY, // @[:@142218.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@142218.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@142218.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@142218.4]
  output         io_M_AXI_0_AWVALID, // @[:@142218.4]
  input          io_M_AXI_0_AWREADY, // @[:@142218.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@142218.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@142218.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@142218.4]
  output         io_M_AXI_0_ARVALID, // @[:@142218.4]
  input          io_M_AXI_0_ARREADY, // @[:@142218.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@142218.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@142218.4]
  output         io_M_AXI_0_WLAST, // @[:@142218.4]
  output         io_M_AXI_0_WVALID, // @[:@142218.4]
  input          io_M_AXI_0_WREADY, // @[:@142218.4]
  output         io_M_AXI_0_RREADY, // @[:@142218.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@142218.4]
  input          io_M_AXI_0_BVALID, // @[:@142218.4]
  output         io_M_AXI_0_BREADY, // @[:@142218.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@142218.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@142218.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@142218.4]
  output         io_M_AXI_1_AWVALID, // @[:@142218.4]
  input          io_M_AXI_1_AWREADY, // @[:@142218.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@142218.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@142218.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@142218.4]
  output         io_M_AXI_1_ARVALID, // @[:@142218.4]
  input          io_M_AXI_1_ARREADY, // @[:@142218.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@142218.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@142218.4]
  output         io_M_AXI_1_WLAST, // @[:@142218.4]
  output         io_M_AXI_1_WVALID, // @[:@142218.4]
  input          io_M_AXI_1_WREADY, // @[:@142218.4]
  output         io_M_AXI_1_RREADY, // @[:@142218.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@142218.4]
  input          io_M_AXI_1_BVALID, // @[:@142218.4]
  output         io_M_AXI_1_BREADY, // @[:@142218.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@142218.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@142218.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@142218.4]
  output         io_M_AXI_2_AWVALID, // @[:@142218.4]
  input          io_M_AXI_2_AWREADY, // @[:@142218.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@142218.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@142218.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@142218.4]
  output         io_M_AXI_2_ARVALID, // @[:@142218.4]
  input          io_M_AXI_2_ARREADY, // @[:@142218.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@142218.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@142218.4]
  output         io_M_AXI_2_WLAST, // @[:@142218.4]
  output         io_M_AXI_2_WVALID, // @[:@142218.4]
  input          io_M_AXI_2_WREADY, // @[:@142218.4]
  output         io_M_AXI_2_RREADY, // @[:@142218.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@142218.4]
  input          io_M_AXI_2_BVALID, // @[:@142218.4]
  output         io_M_AXI_2_BREADY, // @[:@142218.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@142218.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@142218.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@142218.4]
  output         io_M_AXI_3_AWVALID, // @[:@142218.4]
  input          io_M_AXI_3_AWREADY, // @[:@142218.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@142218.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@142218.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@142218.4]
  output         io_M_AXI_3_ARVALID, // @[:@142218.4]
  input          io_M_AXI_3_ARREADY, // @[:@142218.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@142218.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@142218.4]
  output         io_M_AXI_3_WLAST, // @[:@142218.4]
  output         io_M_AXI_3_WVALID, // @[:@142218.4]
  input          io_M_AXI_3_WREADY, // @[:@142218.4]
  output         io_M_AXI_3_RREADY, // @[:@142218.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@142218.4]
  input          io_M_AXI_3_BVALID, // @[:@142218.4]
  output         io_M_AXI_3_BREADY, // @[:@142218.4]
  output         io_enable, // @[:@142218.4]
  input          io_done, // @[:@142218.4]
  output         io_reset, // @[:@142218.4]
  output [63:0]  io_argIns_0, // @[:@142218.4]
  output [63:0]  io_argIns_1, // @[:@142218.4]
  input          io_argOuts_0_valid, // @[:@142218.4]
  input  [63:0]  io_argOuts_0_bits, // @[:@142218.4]
  output         io_memStreams_stores_0_cmd_ready, // @[:@142218.4]
  input          io_memStreams_stores_0_cmd_valid, // @[:@142218.4]
  input  [63:0]  io_memStreams_stores_0_cmd_bits_addr, // @[:@142218.4]
  input  [31:0]  io_memStreams_stores_0_cmd_bits_size, // @[:@142218.4]
  output         io_memStreams_stores_0_data_ready, // @[:@142218.4]
  input          io_memStreams_stores_0_data_valid, // @[:@142218.4]
  input  [31:0]  io_memStreams_stores_0_data_bits_wdata_0, // @[:@142218.4]
  input          io_memStreams_stores_0_data_bits_wstrb, // @[:@142218.4]
  input          io_memStreams_stores_0_wresp_ready, // @[:@142218.4]
  output         io_memStreams_stores_0_wresp_valid, // @[:@142218.4]
  output         io_memStreams_stores_0_wresp_bits, // @[:@142218.4]
  input          io_heap_0_req_valid, // @[:@142218.4]
  input          io_heap_0_req_bits_allocDealloc, // @[:@142218.4]
  input  [63:0]  io_heap_0_req_bits_sizeAddr, // @[:@142218.4]
  output         io_heap_0_resp_valid, // @[:@142218.4]
  output         io_heap_0_resp_bits_allocDealloc, // @[:@142218.4]
  output [63:0]  io_heap_0_resp_bits_sizeAddr // @[:@142218.4]
);
  wire  fringeCommon_clock; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_reset; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_raddr; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_wen; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_waddr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_wdata; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_rdata; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_enable; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_done; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_reset; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_argIns_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_argIns_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_argOuts_0_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_argOuts_0_bits; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_cmd_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_0_wresp_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_0_wresp_bits_tag; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_cmd_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_1_wresp_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_1_wresp_bits_tag; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_cmd_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_2_wresp_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_2_wresp_bits_tag; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_cmd_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_dram_3_wresp_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire [31:0] fringeCommon_io_dram_3_wresp_bits_tag; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_heap_0_req_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 69:28:@142689.4]
  wire  fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 69:28:@142689.4]
  wire [63:0] fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 69:28:@142689.4]
  wire  AXI4LiteToRFBridge_clock; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_reset; // @[FringeZynq.scala 90:31:@143595.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_AWADDR; // @[FringeZynq.scala 90:31:@143595.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_AWPROT; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWVALID; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 90:31:@143595.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_ARADDR; // @[FringeZynq.scala 90:31:@143595.4]
  wire [2:0] AXI4LiteToRFBridge_io_S_AXI_ARPROT; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARVALID; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 90:31:@143595.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_WDATA; // @[FringeZynq.scala 90:31:@143595.4]
  wire [3:0] AXI4LiteToRFBridge_io_S_AXI_WSTRB; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WVALID; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 90:31:@143595.4]
  wire [31:0] AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 90:31:@143595.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_RREADY; // @[FringeZynq.scala 90:31:@143595.4]
  wire [1:0] AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_S_AXI_BREADY; // @[FringeZynq.scala 90:31:@143595.4]
  wire [31:0] AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 90:31:@143595.4]
  wire  AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 90:31:@143595.4]
  wire [31:0] AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 90:31:@143595.4]
  wire [31:0] AXI4LiteToRFBridge_io_wdata; // @[FringeZynq.scala 90:31:@143595.4]
  wire [31:0] AXI4LiteToRFBridge_io_rdata; // @[FringeZynq.scala 90:31:@143595.4]
  wire  MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@143745.4]
  wire [63:0] MAGToAXI4Bridge_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@143745.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@143745.4]
  wire [7:0] MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@143745.4]
  wire [511:0] MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@143745.4]
  wire [63:0] MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@143745.4]
  wire [31:0] MAGToAXI4Bridge_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@143745.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@143901.4]
  wire [63:0] MAGToAXI4Bridge_1_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@143901.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@143901.4]
  wire [7:0] MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@143901.4]
  wire [511:0] MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@143901.4]
  wire [63:0] MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@143901.4]
  wire [31:0] MAGToAXI4Bridge_1_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@143901.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@144057.4]
  wire [63:0] MAGToAXI4Bridge_2_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@144057.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@144057.4]
  wire [7:0] MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@144057.4]
  wire [511:0] MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@144057.4]
  wire [63:0] MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@144057.4]
  wire [31:0] MAGToAXI4Bridge_2_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@144057.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_valid; // @[FringeZynq.scala 131:27:@144213.4]
  wire [63:0] MAGToAXI4Bridge_3_io_in_cmd_bits_addr; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_size; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_cmd_bits_isWr; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_cmd_bits_tag; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_valid; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wdata_bits_wlast; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_rresp_ready; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_ready; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 131:27:@144213.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_AWREADY; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 131:27:@144213.4]
  wire [7:0] MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_ARREADY; // @[FringeZynq.scala 131:27:@144213.4]
  wire [511:0] MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 131:27:@144213.4]
  wire [63:0] MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_WREADY; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 131:27:@144213.4]
  wire [31:0] MAGToAXI4Bridge_3_io_M_AXI_BID; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BVALID; // @[FringeZynq.scala 131:27:@144213.4]
  wire  MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 131:27:@144213.4]
  Fringe fringeCommon ( // @[FringeZynq.scala 69:28:@142689.4]
    .clock(fringeCommon_clock),
    .reset(fringeCommon_reset),
    .io_raddr(fringeCommon_io_raddr),
    .io_wen(fringeCommon_io_wen),
    .io_waddr(fringeCommon_io_waddr),
    .io_wdata(fringeCommon_io_wdata),
    .io_rdata(fringeCommon_io_rdata),
    .io_enable(fringeCommon_io_enable),
    .io_done(fringeCommon_io_done),
    .io_reset(fringeCommon_io_reset),
    .io_argIns_0(fringeCommon_io_argIns_0),
    .io_argIns_1(fringeCommon_io_argIns_1),
    .io_argOuts_0_valid(fringeCommon_io_argOuts_0_valid),
    .io_argOuts_0_bits(fringeCommon_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(fringeCommon_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(fringeCommon_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(fringeCommon_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(fringeCommon_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(fringeCommon_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(fringeCommon_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(fringeCommon_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(fringeCommon_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(fringeCommon_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(fringeCommon_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(fringeCommon_io_memStreams_stores_0_wresp_bits),
    .io_dram_0_cmd_ready(fringeCommon_io_dram_0_cmd_ready),
    .io_dram_0_cmd_valid(fringeCommon_io_dram_0_cmd_valid),
    .io_dram_0_cmd_bits_addr(fringeCommon_io_dram_0_cmd_bits_addr),
    .io_dram_0_cmd_bits_size(fringeCommon_io_dram_0_cmd_bits_size),
    .io_dram_0_cmd_bits_isWr(fringeCommon_io_dram_0_cmd_bits_isWr),
    .io_dram_0_cmd_bits_tag(fringeCommon_io_dram_0_cmd_bits_tag),
    .io_dram_0_wdata_ready(fringeCommon_io_dram_0_wdata_ready),
    .io_dram_0_wdata_valid(fringeCommon_io_dram_0_wdata_valid),
    .io_dram_0_wdata_bits_wdata_0(fringeCommon_io_dram_0_wdata_bits_wdata_0),
    .io_dram_0_wdata_bits_wdata_1(fringeCommon_io_dram_0_wdata_bits_wdata_1),
    .io_dram_0_wdata_bits_wdata_2(fringeCommon_io_dram_0_wdata_bits_wdata_2),
    .io_dram_0_wdata_bits_wdata_3(fringeCommon_io_dram_0_wdata_bits_wdata_3),
    .io_dram_0_wdata_bits_wdata_4(fringeCommon_io_dram_0_wdata_bits_wdata_4),
    .io_dram_0_wdata_bits_wdata_5(fringeCommon_io_dram_0_wdata_bits_wdata_5),
    .io_dram_0_wdata_bits_wdata_6(fringeCommon_io_dram_0_wdata_bits_wdata_6),
    .io_dram_0_wdata_bits_wdata_7(fringeCommon_io_dram_0_wdata_bits_wdata_7),
    .io_dram_0_wdata_bits_wdata_8(fringeCommon_io_dram_0_wdata_bits_wdata_8),
    .io_dram_0_wdata_bits_wdata_9(fringeCommon_io_dram_0_wdata_bits_wdata_9),
    .io_dram_0_wdata_bits_wdata_10(fringeCommon_io_dram_0_wdata_bits_wdata_10),
    .io_dram_0_wdata_bits_wdata_11(fringeCommon_io_dram_0_wdata_bits_wdata_11),
    .io_dram_0_wdata_bits_wdata_12(fringeCommon_io_dram_0_wdata_bits_wdata_12),
    .io_dram_0_wdata_bits_wdata_13(fringeCommon_io_dram_0_wdata_bits_wdata_13),
    .io_dram_0_wdata_bits_wdata_14(fringeCommon_io_dram_0_wdata_bits_wdata_14),
    .io_dram_0_wdata_bits_wdata_15(fringeCommon_io_dram_0_wdata_bits_wdata_15),
    .io_dram_0_wdata_bits_wstrb_0(fringeCommon_io_dram_0_wdata_bits_wstrb_0),
    .io_dram_0_wdata_bits_wstrb_1(fringeCommon_io_dram_0_wdata_bits_wstrb_1),
    .io_dram_0_wdata_bits_wstrb_2(fringeCommon_io_dram_0_wdata_bits_wstrb_2),
    .io_dram_0_wdata_bits_wstrb_3(fringeCommon_io_dram_0_wdata_bits_wstrb_3),
    .io_dram_0_wdata_bits_wstrb_4(fringeCommon_io_dram_0_wdata_bits_wstrb_4),
    .io_dram_0_wdata_bits_wstrb_5(fringeCommon_io_dram_0_wdata_bits_wstrb_5),
    .io_dram_0_wdata_bits_wstrb_6(fringeCommon_io_dram_0_wdata_bits_wstrb_6),
    .io_dram_0_wdata_bits_wstrb_7(fringeCommon_io_dram_0_wdata_bits_wstrb_7),
    .io_dram_0_wdata_bits_wstrb_8(fringeCommon_io_dram_0_wdata_bits_wstrb_8),
    .io_dram_0_wdata_bits_wstrb_9(fringeCommon_io_dram_0_wdata_bits_wstrb_9),
    .io_dram_0_wdata_bits_wstrb_10(fringeCommon_io_dram_0_wdata_bits_wstrb_10),
    .io_dram_0_wdata_bits_wstrb_11(fringeCommon_io_dram_0_wdata_bits_wstrb_11),
    .io_dram_0_wdata_bits_wstrb_12(fringeCommon_io_dram_0_wdata_bits_wstrb_12),
    .io_dram_0_wdata_bits_wstrb_13(fringeCommon_io_dram_0_wdata_bits_wstrb_13),
    .io_dram_0_wdata_bits_wstrb_14(fringeCommon_io_dram_0_wdata_bits_wstrb_14),
    .io_dram_0_wdata_bits_wstrb_15(fringeCommon_io_dram_0_wdata_bits_wstrb_15),
    .io_dram_0_wdata_bits_wstrb_16(fringeCommon_io_dram_0_wdata_bits_wstrb_16),
    .io_dram_0_wdata_bits_wstrb_17(fringeCommon_io_dram_0_wdata_bits_wstrb_17),
    .io_dram_0_wdata_bits_wstrb_18(fringeCommon_io_dram_0_wdata_bits_wstrb_18),
    .io_dram_0_wdata_bits_wstrb_19(fringeCommon_io_dram_0_wdata_bits_wstrb_19),
    .io_dram_0_wdata_bits_wstrb_20(fringeCommon_io_dram_0_wdata_bits_wstrb_20),
    .io_dram_0_wdata_bits_wstrb_21(fringeCommon_io_dram_0_wdata_bits_wstrb_21),
    .io_dram_0_wdata_bits_wstrb_22(fringeCommon_io_dram_0_wdata_bits_wstrb_22),
    .io_dram_0_wdata_bits_wstrb_23(fringeCommon_io_dram_0_wdata_bits_wstrb_23),
    .io_dram_0_wdata_bits_wstrb_24(fringeCommon_io_dram_0_wdata_bits_wstrb_24),
    .io_dram_0_wdata_bits_wstrb_25(fringeCommon_io_dram_0_wdata_bits_wstrb_25),
    .io_dram_0_wdata_bits_wstrb_26(fringeCommon_io_dram_0_wdata_bits_wstrb_26),
    .io_dram_0_wdata_bits_wstrb_27(fringeCommon_io_dram_0_wdata_bits_wstrb_27),
    .io_dram_0_wdata_bits_wstrb_28(fringeCommon_io_dram_0_wdata_bits_wstrb_28),
    .io_dram_0_wdata_bits_wstrb_29(fringeCommon_io_dram_0_wdata_bits_wstrb_29),
    .io_dram_0_wdata_bits_wstrb_30(fringeCommon_io_dram_0_wdata_bits_wstrb_30),
    .io_dram_0_wdata_bits_wstrb_31(fringeCommon_io_dram_0_wdata_bits_wstrb_31),
    .io_dram_0_wdata_bits_wstrb_32(fringeCommon_io_dram_0_wdata_bits_wstrb_32),
    .io_dram_0_wdata_bits_wstrb_33(fringeCommon_io_dram_0_wdata_bits_wstrb_33),
    .io_dram_0_wdata_bits_wstrb_34(fringeCommon_io_dram_0_wdata_bits_wstrb_34),
    .io_dram_0_wdata_bits_wstrb_35(fringeCommon_io_dram_0_wdata_bits_wstrb_35),
    .io_dram_0_wdata_bits_wstrb_36(fringeCommon_io_dram_0_wdata_bits_wstrb_36),
    .io_dram_0_wdata_bits_wstrb_37(fringeCommon_io_dram_0_wdata_bits_wstrb_37),
    .io_dram_0_wdata_bits_wstrb_38(fringeCommon_io_dram_0_wdata_bits_wstrb_38),
    .io_dram_0_wdata_bits_wstrb_39(fringeCommon_io_dram_0_wdata_bits_wstrb_39),
    .io_dram_0_wdata_bits_wstrb_40(fringeCommon_io_dram_0_wdata_bits_wstrb_40),
    .io_dram_0_wdata_bits_wstrb_41(fringeCommon_io_dram_0_wdata_bits_wstrb_41),
    .io_dram_0_wdata_bits_wstrb_42(fringeCommon_io_dram_0_wdata_bits_wstrb_42),
    .io_dram_0_wdata_bits_wstrb_43(fringeCommon_io_dram_0_wdata_bits_wstrb_43),
    .io_dram_0_wdata_bits_wstrb_44(fringeCommon_io_dram_0_wdata_bits_wstrb_44),
    .io_dram_0_wdata_bits_wstrb_45(fringeCommon_io_dram_0_wdata_bits_wstrb_45),
    .io_dram_0_wdata_bits_wstrb_46(fringeCommon_io_dram_0_wdata_bits_wstrb_46),
    .io_dram_0_wdata_bits_wstrb_47(fringeCommon_io_dram_0_wdata_bits_wstrb_47),
    .io_dram_0_wdata_bits_wstrb_48(fringeCommon_io_dram_0_wdata_bits_wstrb_48),
    .io_dram_0_wdata_bits_wstrb_49(fringeCommon_io_dram_0_wdata_bits_wstrb_49),
    .io_dram_0_wdata_bits_wstrb_50(fringeCommon_io_dram_0_wdata_bits_wstrb_50),
    .io_dram_0_wdata_bits_wstrb_51(fringeCommon_io_dram_0_wdata_bits_wstrb_51),
    .io_dram_0_wdata_bits_wstrb_52(fringeCommon_io_dram_0_wdata_bits_wstrb_52),
    .io_dram_0_wdata_bits_wstrb_53(fringeCommon_io_dram_0_wdata_bits_wstrb_53),
    .io_dram_0_wdata_bits_wstrb_54(fringeCommon_io_dram_0_wdata_bits_wstrb_54),
    .io_dram_0_wdata_bits_wstrb_55(fringeCommon_io_dram_0_wdata_bits_wstrb_55),
    .io_dram_0_wdata_bits_wstrb_56(fringeCommon_io_dram_0_wdata_bits_wstrb_56),
    .io_dram_0_wdata_bits_wstrb_57(fringeCommon_io_dram_0_wdata_bits_wstrb_57),
    .io_dram_0_wdata_bits_wstrb_58(fringeCommon_io_dram_0_wdata_bits_wstrb_58),
    .io_dram_0_wdata_bits_wstrb_59(fringeCommon_io_dram_0_wdata_bits_wstrb_59),
    .io_dram_0_wdata_bits_wstrb_60(fringeCommon_io_dram_0_wdata_bits_wstrb_60),
    .io_dram_0_wdata_bits_wstrb_61(fringeCommon_io_dram_0_wdata_bits_wstrb_61),
    .io_dram_0_wdata_bits_wstrb_62(fringeCommon_io_dram_0_wdata_bits_wstrb_62),
    .io_dram_0_wdata_bits_wstrb_63(fringeCommon_io_dram_0_wdata_bits_wstrb_63),
    .io_dram_0_wdata_bits_wlast(fringeCommon_io_dram_0_wdata_bits_wlast),
    .io_dram_0_rresp_ready(fringeCommon_io_dram_0_rresp_ready),
    .io_dram_0_wresp_ready(fringeCommon_io_dram_0_wresp_ready),
    .io_dram_0_wresp_valid(fringeCommon_io_dram_0_wresp_valid),
    .io_dram_0_wresp_bits_tag(fringeCommon_io_dram_0_wresp_bits_tag),
    .io_dram_1_cmd_ready(fringeCommon_io_dram_1_cmd_ready),
    .io_dram_1_cmd_valid(fringeCommon_io_dram_1_cmd_valid),
    .io_dram_1_cmd_bits_addr(fringeCommon_io_dram_1_cmd_bits_addr),
    .io_dram_1_cmd_bits_size(fringeCommon_io_dram_1_cmd_bits_size),
    .io_dram_1_cmd_bits_isWr(fringeCommon_io_dram_1_cmd_bits_isWr),
    .io_dram_1_cmd_bits_tag(fringeCommon_io_dram_1_cmd_bits_tag),
    .io_dram_1_wdata_ready(fringeCommon_io_dram_1_wdata_ready),
    .io_dram_1_wdata_valid(fringeCommon_io_dram_1_wdata_valid),
    .io_dram_1_wdata_bits_wdata_0(fringeCommon_io_dram_1_wdata_bits_wdata_0),
    .io_dram_1_wdata_bits_wdata_1(fringeCommon_io_dram_1_wdata_bits_wdata_1),
    .io_dram_1_wdata_bits_wdata_2(fringeCommon_io_dram_1_wdata_bits_wdata_2),
    .io_dram_1_wdata_bits_wdata_3(fringeCommon_io_dram_1_wdata_bits_wdata_3),
    .io_dram_1_wdata_bits_wdata_4(fringeCommon_io_dram_1_wdata_bits_wdata_4),
    .io_dram_1_wdata_bits_wdata_5(fringeCommon_io_dram_1_wdata_bits_wdata_5),
    .io_dram_1_wdata_bits_wdata_6(fringeCommon_io_dram_1_wdata_bits_wdata_6),
    .io_dram_1_wdata_bits_wdata_7(fringeCommon_io_dram_1_wdata_bits_wdata_7),
    .io_dram_1_wdata_bits_wdata_8(fringeCommon_io_dram_1_wdata_bits_wdata_8),
    .io_dram_1_wdata_bits_wdata_9(fringeCommon_io_dram_1_wdata_bits_wdata_9),
    .io_dram_1_wdata_bits_wdata_10(fringeCommon_io_dram_1_wdata_bits_wdata_10),
    .io_dram_1_wdata_bits_wdata_11(fringeCommon_io_dram_1_wdata_bits_wdata_11),
    .io_dram_1_wdata_bits_wdata_12(fringeCommon_io_dram_1_wdata_bits_wdata_12),
    .io_dram_1_wdata_bits_wdata_13(fringeCommon_io_dram_1_wdata_bits_wdata_13),
    .io_dram_1_wdata_bits_wdata_14(fringeCommon_io_dram_1_wdata_bits_wdata_14),
    .io_dram_1_wdata_bits_wdata_15(fringeCommon_io_dram_1_wdata_bits_wdata_15),
    .io_dram_1_wdata_bits_wstrb_0(fringeCommon_io_dram_1_wdata_bits_wstrb_0),
    .io_dram_1_wdata_bits_wstrb_1(fringeCommon_io_dram_1_wdata_bits_wstrb_1),
    .io_dram_1_wdata_bits_wstrb_2(fringeCommon_io_dram_1_wdata_bits_wstrb_2),
    .io_dram_1_wdata_bits_wstrb_3(fringeCommon_io_dram_1_wdata_bits_wstrb_3),
    .io_dram_1_wdata_bits_wstrb_4(fringeCommon_io_dram_1_wdata_bits_wstrb_4),
    .io_dram_1_wdata_bits_wstrb_5(fringeCommon_io_dram_1_wdata_bits_wstrb_5),
    .io_dram_1_wdata_bits_wstrb_6(fringeCommon_io_dram_1_wdata_bits_wstrb_6),
    .io_dram_1_wdata_bits_wstrb_7(fringeCommon_io_dram_1_wdata_bits_wstrb_7),
    .io_dram_1_wdata_bits_wstrb_8(fringeCommon_io_dram_1_wdata_bits_wstrb_8),
    .io_dram_1_wdata_bits_wstrb_9(fringeCommon_io_dram_1_wdata_bits_wstrb_9),
    .io_dram_1_wdata_bits_wstrb_10(fringeCommon_io_dram_1_wdata_bits_wstrb_10),
    .io_dram_1_wdata_bits_wstrb_11(fringeCommon_io_dram_1_wdata_bits_wstrb_11),
    .io_dram_1_wdata_bits_wstrb_12(fringeCommon_io_dram_1_wdata_bits_wstrb_12),
    .io_dram_1_wdata_bits_wstrb_13(fringeCommon_io_dram_1_wdata_bits_wstrb_13),
    .io_dram_1_wdata_bits_wstrb_14(fringeCommon_io_dram_1_wdata_bits_wstrb_14),
    .io_dram_1_wdata_bits_wstrb_15(fringeCommon_io_dram_1_wdata_bits_wstrb_15),
    .io_dram_1_wdata_bits_wstrb_16(fringeCommon_io_dram_1_wdata_bits_wstrb_16),
    .io_dram_1_wdata_bits_wstrb_17(fringeCommon_io_dram_1_wdata_bits_wstrb_17),
    .io_dram_1_wdata_bits_wstrb_18(fringeCommon_io_dram_1_wdata_bits_wstrb_18),
    .io_dram_1_wdata_bits_wstrb_19(fringeCommon_io_dram_1_wdata_bits_wstrb_19),
    .io_dram_1_wdata_bits_wstrb_20(fringeCommon_io_dram_1_wdata_bits_wstrb_20),
    .io_dram_1_wdata_bits_wstrb_21(fringeCommon_io_dram_1_wdata_bits_wstrb_21),
    .io_dram_1_wdata_bits_wstrb_22(fringeCommon_io_dram_1_wdata_bits_wstrb_22),
    .io_dram_1_wdata_bits_wstrb_23(fringeCommon_io_dram_1_wdata_bits_wstrb_23),
    .io_dram_1_wdata_bits_wstrb_24(fringeCommon_io_dram_1_wdata_bits_wstrb_24),
    .io_dram_1_wdata_bits_wstrb_25(fringeCommon_io_dram_1_wdata_bits_wstrb_25),
    .io_dram_1_wdata_bits_wstrb_26(fringeCommon_io_dram_1_wdata_bits_wstrb_26),
    .io_dram_1_wdata_bits_wstrb_27(fringeCommon_io_dram_1_wdata_bits_wstrb_27),
    .io_dram_1_wdata_bits_wstrb_28(fringeCommon_io_dram_1_wdata_bits_wstrb_28),
    .io_dram_1_wdata_bits_wstrb_29(fringeCommon_io_dram_1_wdata_bits_wstrb_29),
    .io_dram_1_wdata_bits_wstrb_30(fringeCommon_io_dram_1_wdata_bits_wstrb_30),
    .io_dram_1_wdata_bits_wstrb_31(fringeCommon_io_dram_1_wdata_bits_wstrb_31),
    .io_dram_1_wdata_bits_wstrb_32(fringeCommon_io_dram_1_wdata_bits_wstrb_32),
    .io_dram_1_wdata_bits_wstrb_33(fringeCommon_io_dram_1_wdata_bits_wstrb_33),
    .io_dram_1_wdata_bits_wstrb_34(fringeCommon_io_dram_1_wdata_bits_wstrb_34),
    .io_dram_1_wdata_bits_wstrb_35(fringeCommon_io_dram_1_wdata_bits_wstrb_35),
    .io_dram_1_wdata_bits_wstrb_36(fringeCommon_io_dram_1_wdata_bits_wstrb_36),
    .io_dram_1_wdata_bits_wstrb_37(fringeCommon_io_dram_1_wdata_bits_wstrb_37),
    .io_dram_1_wdata_bits_wstrb_38(fringeCommon_io_dram_1_wdata_bits_wstrb_38),
    .io_dram_1_wdata_bits_wstrb_39(fringeCommon_io_dram_1_wdata_bits_wstrb_39),
    .io_dram_1_wdata_bits_wstrb_40(fringeCommon_io_dram_1_wdata_bits_wstrb_40),
    .io_dram_1_wdata_bits_wstrb_41(fringeCommon_io_dram_1_wdata_bits_wstrb_41),
    .io_dram_1_wdata_bits_wstrb_42(fringeCommon_io_dram_1_wdata_bits_wstrb_42),
    .io_dram_1_wdata_bits_wstrb_43(fringeCommon_io_dram_1_wdata_bits_wstrb_43),
    .io_dram_1_wdata_bits_wstrb_44(fringeCommon_io_dram_1_wdata_bits_wstrb_44),
    .io_dram_1_wdata_bits_wstrb_45(fringeCommon_io_dram_1_wdata_bits_wstrb_45),
    .io_dram_1_wdata_bits_wstrb_46(fringeCommon_io_dram_1_wdata_bits_wstrb_46),
    .io_dram_1_wdata_bits_wstrb_47(fringeCommon_io_dram_1_wdata_bits_wstrb_47),
    .io_dram_1_wdata_bits_wstrb_48(fringeCommon_io_dram_1_wdata_bits_wstrb_48),
    .io_dram_1_wdata_bits_wstrb_49(fringeCommon_io_dram_1_wdata_bits_wstrb_49),
    .io_dram_1_wdata_bits_wstrb_50(fringeCommon_io_dram_1_wdata_bits_wstrb_50),
    .io_dram_1_wdata_bits_wstrb_51(fringeCommon_io_dram_1_wdata_bits_wstrb_51),
    .io_dram_1_wdata_bits_wstrb_52(fringeCommon_io_dram_1_wdata_bits_wstrb_52),
    .io_dram_1_wdata_bits_wstrb_53(fringeCommon_io_dram_1_wdata_bits_wstrb_53),
    .io_dram_1_wdata_bits_wstrb_54(fringeCommon_io_dram_1_wdata_bits_wstrb_54),
    .io_dram_1_wdata_bits_wstrb_55(fringeCommon_io_dram_1_wdata_bits_wstrb_55),
    .io_dram_1_wdata_bits_wstrb_56(fringeCommon_io_dram_1_wdata_bits_wstrb_56),
    .io_dram_1_wdata_bits_wstrb_57(fringeCommon_io_dram_1_wdata_bits_wstrb_57),
    .io_dram_1_wdata_bits_wstrb_58(fringeCommon_io_dram_1_wdata_bits_wstrb_58),
    .io_dram_1_wdata_bits_wstrb_59(fringeCommon_io_dram_1_wdata_bits_wstrb_59),
    .io_dram_1_wdata_bits_wstrb_60(fringeCommon_io_dram_1_wdata_bits_wstrb_60),
    .io_dram_1_wdata_bits_wstrb_61(fringeCommon_io_dram_1_wdata_bits_wstrb_61),
    .io_dram_1_wdata_bits_wstrb_62(fringeCommon_io_dram_1_wdata_bits_wstrb_62),
    .io_dram_1_wdata_bits_wstrb_63(fringeCommon_io_dram_1_wdata_bits_wstrb_63),
    .io_dram_1_wdata_bits_wlast(fringeCommon_io_dram_1_wdata_bits_wlast),
    .io_dram_1_rresp_ready(fringeCommon_io_dram_1_rresp_ready),
    .io_dram_1_wresp_ready(fringeCommon_io_dram_1_wresp_ready),
    .io_dram_1_wresp_valid(fringeCommon_io_dram_1_wresp_valid),
    .io_dram_1_wresp_bits_tag(fringeCommon_io_dram_1_wresp_bits_tag),
    .io_dram_2_cmd_ready(fringeCommon_io_dram_2_cmd_ready),
    .io_dram_2_cmd_valid(fringeCommon_io_dram_2_cmd_valid),
    .io_dram_2_cmd_bits_addr(fringeCommon_io_dram_2_cmd_bits_addr),
    .io_dram_2_cmd_bits_size(fringeCommon_io_dram_2_cmd_bits_size),
    .io_dram_2_cmd_bits_isWr(fringeCommon_io_dram_2_cmd_bits_isWr),
    .io_dram_2_cmd_bits_tag(fringeCommon_io_dram_2_cmd_bits_tag),
    .io_dram_2_wdata_ready(fringeCommon_io_dram_2_wdata_ready),
    .io_dram_2_wdata_valid(fringeCommon_io_dram_2_wdata_valid),
    .io_dram_2_wdata_bits_wdata_0(fringeCommon_io_dram_2_wdata_bits_wdata_0),
    .io_dram_2_wdata_bits_wdata_1(fringeCommon_io_dram_2_wdata_bits_wdata_1),
    .io_dram_2_wdata_bits_wdata_2(fringeCommon_io_dram_2_wdata_bits_wdata_2),
    .io_dram_2_wdata_bits_wdata_3(fringeCommon_io_dram_2_wdata_bits_wdata_3),
    .io_dram_2_wdata_bits_wdata_4(fringeCommon_io_dram_2_wdata_bits_wdata_4),
    .io_dram_2_wdata_bits_wdata_5(fringeCommon_io_dram_2_wdata_bits_wdata_5),
    .io_dram_2_wdata_bits_wdata_6(fringeCommon_io_dram_2_wdata_bits_wdata_6),
    .io_dram_2_wdata_bits_wdata_7(fringeCommon_io_dram_2_wdata_bits_wdata_7),
    .io_dram_2_wdata_bits_wdata_8(fringeCommon_io_dram_2_wdata_bits_wdata_8),
    .io_dram_2_wdata_bits_wdata_9(fringeCommon_io_dram_2_wdata_bits_wdata_9),
    .io_dram_2_wdata_bits_wdata_10(fringeCommon_io_dram_2_wdata_bits_wdata_10),
    .io_dram_2_wdata_bits_wdata_11(fringeCommon_io_dram_2_wdata_bits_wdata_11),
    .io_dram_2_wdata_bits_wdata_12(fringeCommon_io_dram_2_wdata_bits_wdata_12),
    .io_dram_2_wdata_bits_wdata_13(fringeCommon_io_dram_2_wdata_bits_wdata_13),
    .io_dram_2_wdata_bits_wdata_14(fringeCommon_io_dram_2_wdata_bits_wdata_14),
    .io_dram_2_wdata_bits_wdata_15(fringeCommon_io_dram_2_wdata_bits_wdata_15),
    .io_dram_2_wdata_bits_wstrb_0(fringeCommon_io_dram_2_wdata_bits_wstrb_0),
    .io_dram_2_wdata_bits_wstrb_1(fringeCommon_io_dram_2_wdata_bits_wstrb_1),
    .io_dram_2_wdata_bits_wstrb_2(fringeCommon_io_dram_2_wdata_bits_wstrb_2),
    .io_dram_2_wdata_bits_wstrb_3(fringeCommon_io_dram_2_wdata_bits_wstrb_3),
    .io_dram_2_wdata_bits_wstrb_4(fringeCommon_io_dram_2_wdata_bits_wstrb_4),
    .io_dram_2_wdata_bits_wstrb_5(fringeCommon_io_dram_2_wdata_bits_wstrb_5),
    .io_dram_2_wdata_bits_wstrb_6(fringeCommon_io_dram_2_wdata_bits_wstrb_6),
    .io_dram_2_wdata_bits_wstrb_7(fringeCommon_io_dram_2_wdata_bits_wstrb_7),
    .io_dram_2_wdata_bits_wstrb_8(fringeCommon_io_dram_2_wdata_bits_wstrb_8),
    .io_dram_2_wdata_bits_wstrb_9(fringeCommon_io_dram_2_wdata_bits_wstrb_9),
    .io_dram_2_wdata_bits_wstrb_10(fringeCommon_io_dram_2_wdata_bits_wstrb_10),
    .io_dram_2_wdata_bits_wstrb_11(fringeCommon_io_dram_2_wdata_bits_wstrb_11),
    .io_dram_2_wdata_bits_wstrb_12(fringeCommon_io_dram_2_wdata_bits_wstrb_12),
    .io_dram_2_wdata_bits_wstrb_13(fringeCommon_io_dram_2_wdata_bits_wstrb_13),
    .io_dram_2_wdata_bits_wstrb_14(fringeCommon_io_dram_2_wdata_bits_wstrb_14),
    .io_dram_2_wdata_bits_wstrb_15(fringeCommon_io_dram_2_wdata_bits_wstrb_15),
    .io_dram_2_wdata_bits_wstrb_16(fringeCommon_io_dram_2_wdata_bits_wstrb_16),
    .io_dram_2_wdata_bits_wstrb_17(fringeCommon_io_dram_2_wdata_bits_wstrb_17),
    .io_dram_2_wdata_bits_wstrb_18(fringeCommon_io_dram_2_wdata_bits_wstrb_18),
    .io_dram_2_wdata_bits_wstrb_19(fringeCommon_io_dram_2_wdata_bits_wstrb_19),
    .io_dram_2_wdata_bits_wstrb_20(fringeCommon_io_dram_2_wdata_bits_wstrb_20),
    .io_dram_2_wdata_bits_wstrb_21(fringeCommon_io_dram_2_wdata_bits_wstrb_21),
    .io_dram_2_wdata_bits_wstrb_22(fringeCommon_io_dram_2_wdata_bits_wstrb_22),
    .io_dram_2_wdata_bits_wstrb_23(fringeCommon_io_dram_2_wdata_bits_wstrb_23),
    .io_dram_2_wdata_bits_wstrb_24(fringeCommon_io_dram_2_wdata_bits_wstrb_24),
    .io_dram_2_wdata_bits_wstrb_25(fringeCommon_io_dram_2_wdata_bits_wstrb_25),
    .io_dram_2_wdata_bits_wstrb_26(fringeCommon_io_dram_2_wdata_bits_wstrb_26),
    .io_dram_2_wdata_bits_wstrb_27(fringeCommon_io_dram_2_wdata_bits_wstrb_27),
    .io_dram_2_wdata_bits_wstrb_28(fringeCommon_io_dram_2_wdata_bits_wstrb_28),
    .io_dram_2_wdata_bits_wstrb_29(fringeCommon_io_dram_2_wdata_bits_wstrb_29),
    .io_dram_2_wdata_bits_wstrb_30(fringeCommon_io_dram_2_wdata_bits_wstrb_30),
    .io_dram_2_wdata_bits_wstrb_31(fringeCommon_io_dram_2_wdata_bits_wstrb_31),
    .io_dram_2_wdata_bits_wstrb_32(fringeCommon_io_dram_2_wdata_bits_wstrb_32),
    .io_dram_2_wdata_bits_wstrb_33(fringeCommon_io_dram_2_wdata_bits_wstrb_33),
    .io_dram_2_wdata_bits_wstrb_34(fringeCommon_io_dram_2_wdata_bits_wstrb_34),
    .io_dram_2_wdata_bits_wstrb_35(fringeCommon_io_dram_2_wdata_bits_wstrb_35),
    .io_dram_2_wdata_bits_wstrb_36(fringeCommon_io_dram_2_wdata_bits_wstrb_36),
    .io_dram_2_wdata_bits_wstrb_37(fringeCommon_io_dram_2_wdata_bits_wstrb_37),
    .io_dram_2_wdata_bits_wstrb_38(fringeCommon_io_dram_2_wdata_bits_wstrb_38),
    .io_dram_2_wdata_bits_wstrb_39(fringeCommon_io_dram_2_wdata_bits_wstrb_39),
    .io_dram_2_wdata_bits_wstrb_40(fringeCommon_io_dram_2_wdata_bits_wstrb_40),
    .io_dram_2_wdata_bits_wstrb_41(fringeCommon_io_dram_2_wdata_bits_wstrb_41),
    .io_dram_2_wdata_bits_wstrb_42(fringeCommon_io_dram_2_wdata_bits_wstrb_42),
    .io_dram_2_wdata_bits_wstrb_43(fringeCommon_io_dram_2_wdata_bits_wstrb_43),
    .io_dram_2_wdata_bits_wstrb_44(fringeCommon_io_dram_2_wdata_bits_wstrb_44),
    .io_dram_2_wdata_bits_wstrb_45(fringeCommon_io_dram_2_wdata_bits_wstrb_45),
    .io_dram_2_wdata_bits_wstrb_46(fringeCommon_io_dram_2_wdata_bits_wstrb_46),
    .io_dram_2_wdata_bits_wstrb_47(fringeCommon_io_dram_2_wdata_bits_wstrb_47),
    .io_dram_2_wdata_bits_wstrb_48(fringeCommon_io_dram_2_wdata_bits_wstrb_48),
    .io_dram_2_wdata_bits_wstrb_49(fringeCommon_io_dram_2_wdata_bits_wstrb_49),
    .io_dram_2_wdata_bits_wstrb_50(fringeCommon_io_dram_2_wdata_bits_wstrb_50),
    .io_dram_2_wdata_bits_wstrb_51(fringeCommon_io_dram_2_wdata_bits_wstrb_51),
    .io_dram_2_wdata_bits_wstrb_52(fringeCommon_io_dram_2_wdata_bits_wstrb_52),
    .io_dram_2_wdata_bits_wstrb_53(fringeCommon_io_dram_2_wdata_bits_wstrb_53),
    .io_dram_2_wdata_bits_wstrb_54(fringeCommon_io_dram_2_wdata_bits_wstrb_54),
    .io_dram_2_wdata_bits_wstrb_55(fringeCommon_io_dram_2_wdata_bits_wstrb_55),
    .io_dram_2_wdata_bits_wstrb_56(fringeCommon_io_dram_2_wdata_bits_wstrb_56),
    .io_dram_2_wdata_bits_wstrb_57(fringeCommon_io_dram_2_wdata_bits_wstrb_57),
    .io_dram_2_wdata_bits_wstrb_58(fringeCommon_io_dram_2_wdata_bits_wstrb_58),
    .io_dram_2_wdata_bits_wstrb_59(fringeCommon_io_dram_2_wdata_bits_wstrb_59),
    .io_dram_2_wdata_bits_wstrb_60(fringeCommon_io_dram_2_wdata_bits_wstrb_60),
    .io_dram_2_wdata_bits_wstrb_61(fringeCommon_io_dram_2_wdata_bits_wstrb_61),
    .io_dram_2_wdata_bits_wstrb_62(fringeCommon_io_dram_2_wdata_bits_wstrb_62),
    .io_dram_2_wdata_bits_wstrb_63(fringeCommon_io_dram_2_wdata_bits_wstrb_63),
    .io_dram_2_wdata_bits_wlast(fringeCommon_io_dram_2_wdata_bits_wlast),
    .io_dram_2_rresp_ready(fringeCommon_io_dram_2_rresp_ready),
    .io_dram_2_wresp_ready(fringeCommon_io_dram_2_wresp_ready),
    .io_dram_2_wresp_valid(fringeCommon_io_dram_2_wresp_valid),
    .io_dram_2_wresp_bits_tag(fringeCommon_io_dram_2_wresp_bits_tag),
    .io_dram_3_cmd_ready(fringeCommon_io_dram_3_cmd_ready),
    .io_dram_3_cmd_valid(fringeCommon_io_dram_3_cmd_valid),
    .io_dram_3_cmd_bits_addr(fringeCommon_io_dram_3_cmd_bits_addr),
    .io_dram_3_cmd_bits_size(fringeCommon_io_dram_3_cmd_bits_size),
    .io_dram_3_cmd_bits_isWr(fringeCommon_io_dram_3_cmd_bits_isWr),
    .io_dram_3_cmd_bits_tag(fringeCommon_io_dram_3_cmd_bits_tag),
    .io_dram_3_wdata_ready(fringeCommon_io_dram_3_wdata_ready),
    .io_dram_3_wdata_valid(fringeCommon_io_dram_3_wdata_valid),
    .io_dram_3_wdata_bits_wdata_0(fringeCommon_io_dram_3_wdata_bits_wdata_0),
    .io_dram_3_wdata_bits_wdata_1(fringeCommon_io_dram_3_wdata_bits_wdata_1),
    .io_dram_3_wdata_bits_wdata_2(fringeCommon_io_dram_3_wdata_bits_wdata_2),
    .io_dram_3_wdata_bits_wdata_3(fringeCommon_io_dram_3_wdata_bits_wdata_3),
    .io_dram_3_wdata_bits_wdata_4(fringeCommon_io_dram_3_wdata_bits_wdata_4),
    .io_dram_3_wdata_bits_wdata_5(fringeCommon_io_dram_3_wdata_bits_wdata_5),
    .io_dram_3_wdata_bits_wdata_6(fringeCommon_io_dram_3_wdata_bits_wdata_6),
    .io_dram_3_wdata_bits_wdata_7(fringeCommon_io_dram_3_wdata_bits_wdata_7),
    .io_dram_3_wdata_bits_wdata_8(fringeCommon_io_dram_3_wdata_bits_wdata_8),
    .io_dram_3_wdata_bits_wdata_9(fringeCommon_io_dram_3_wdata_bits_wdata_9),
    .io_dram_3_wdata_bits_wdata_10(fringeCommon_io_dram_3_wdata_bits_wdata_10),
    .io_dram_3_wdata_bits_wdata_11(fringeCommon_io_dram_3_wdata_bits_wdata_11),
    .io_dram_3_wdata_bits_wdata_12(fringeCommon_io_dram_3_wdata_bits_wdata_12),
    .io_dram_3_wdata_bits_wdata_13(fringeCommon_io_dram_3_wdata_bits_wdata_13),
    .io_dram_3_wdata_bits_wdata_14(fringeCommon_io_dram_3_wdata_bits_wdata_14),
    .io_dram_3_wdata_bits_wdata_15(fringeCommon_io_dram_3_wdata_bits_wdata_15),
    .io_dram_3_wdata_bits_wstrb_0(fringeCommon_io_dram_3_wdata_bits_wstrb_0),
    .io_dram_3_wdata_bits_wstrb_1(fringeCommon_io_dram_3_wdata_bits_wstrb_1),
    .io_dram_3_wdata_bits_wstrb_2(fringeCommon_io_dram_3_wdata_bits_wstrb_2),
    .io_dram_3_wdata_bits_wstrb_3(fringeCommon_io_dram_3_wdata_bits_wstrb_3),
    .io_dram_3_wdata_bits_wstrb_4(fringeCommon_io_dram_3_wdata_bits_wstrb_4),
    .io_dram_3_wdata_bits_wstrb_5(fringeCommon_io_dram_3_wdata_bits_wstrb_5),
    .io_dram_3_wdata_bits_wstrb_6(fringeCommon_io_dram_3_wdata_bits_wstrb_6),
    .io_dram_3_wdata_bits_wstrb_7(fringeCommon_io_dram_3_wdata_bits_wstrb_7),
    .io_dram_3_wdata_bits_wstrb_8(fringeCommon_io_dram_3_wdata_bits_wstrb_8),
    .io_dram_3_wdata_bits_wstrb_9(fringeCommon_io_dram_3_wdata_bits_wstrb_9),
    .io_dram_3_wdata_bits_wstrb_10(fringeCommon_io_dram_3_wdata_bits_wstrb_10),
    .io_dram_3_wdata_bits_wstrb_11(fringeCommon_io_dram_3_wdata_bits_wstrb_11),
    .io_dram_3_wdata_bits_wstrb_12(fringeCommon_io_dram_3_wdata_bits_wstrb_12),
    .io_dram_3_wdata_bits_wstrb_13(fringeCommon_io_dram_3_wdata_bits_wstrb_13),
    .io_dram_3_wdata_bits_wstrb_14(fringeCommon_io_dram_3_wdata_bits_wstrb_14),
    .io_dram_3_wdata_bits_wstrb_15(fringeCommon_io_dram_3_wdata_bits_wstrb_15),
    .io_dram_3_wdata_bits_wstrb_16(fringeCommon_io_dram_3_wdata_bits_wstrb_16),
    .io_dram_3_wdata_bits_wstrb_17(fringeCommon_io_dram_3_wdata_bits_wstrb_17),
    .io_dram_3_wdata_bits_wstrb_18(fringeCommon_io_dram_3_wdata_bits_wstrb_18),
    .io_dram_3_wdata_bits_wstrb_19(fringeCommon_io_dram_3_wdata_bits_wstrb_19),
    .io_dram_3_wdata_bits_wstrb_20(fringeCommon_io_dram_3_wdata_bits_wstrb_20),
    .io_dram_3_wdata_bits_wstrb_21(fringeCommon_io_dram_3_wdata_bits_wstrb_21),
    .io_dram_3_wdata_bits_wstrb_22(fringeCommon_io_dram_3_wdata_bits_wstrb_22),
    .io_dram_3_wdata_bits_wstrb_23(fringeCommon_io_dram_3_wdata_bits_wstrb_23),
    .io_dram_3_wdata_bits_wstrb_24(fringeCommon_io_dram_3_wdata_bits_wstrb_24),
    .io_dram_3_wdata_bits_wstrb_25(fringeCommon_io_dram_3_wdata_bits_wstrb_25),
    .io_dram_3_wdata_bits_wstrb_26(fringeCommon_io_dram_3_wdata_bits_wstrb_26),
    .io_dram_3_wdata_bits_wstrb_27(fringeCommon_io_dram_3_wdata_bits_wstrb_27),
    .io_dram_3_wdata_bits_wstrb_28(fringeCommon_io_dram_3_wdata_bits_wstrb_28),
    .io_dram_3_wdata_bits_wstrb_29(fringeCommon_io_dram_3_wdata_bits_wstrb_29),
    .io_dram_3_wdata_bits_wstrb_30(fringeCommon_io_dram_3_wdata_bits_wstrb_30),
    .io_dram_3_wdata_bits_wstrb_31(fringeCommon_io_dram_3_wdata_bits_wstrb_31),
    .io_dram_3_wdata_bits_wstrb_32(fringeCommon_io_dram_3_wdata_bits_wstrb_32),
    .io_dram_3_wdata_bits_wstrb_33(fringeCommon_io_dram_3_wdata_bits_wstrb_33),
    .io_dram_3_wdata_bits_wstrb_34(fringeCommon_io_dram_3_wdata_bits_wstrb_34),
    .io_dram_3_wdata_bits_wstrb_35(fringeCommon_io_dram_3_wdata_bits_wstrb_35),
    .io_dram_3_wdata_bits_wstrb_36(fringeCommon_io_dram_3_wdata_bits_wstrb_36),
    .io_dram_3_wdata_bits_wstrb_37(fringeCommon_io_dram_3_wdata_bits_wstrb_37),
    .io_dram_3_wdata_bits_wstrb_38(fringeCommon_io_dram_3_wdata_bits_wstrb_38),
    .io_dram_3_wdata_bits_wstrb_39(fringeCommon_io_dram_3_wdata_bits_wstrb_39),
    .io_dram_3_wdata_bits_wstrb_40(fringeCommon_io_dram_3_wdata_bits_wstrb_40),
    .io_dram_3_wdata_bits_wstrb_41(fringeCommon_io_dram_3_wdata_bits_wstrb_41),
    .io_dram_3_wdata_bits_wstrb_42(fringeCommon_io_dram_3_wdata_bits_wstrb_42),
    .io_dram_3_wdata_bits_wstrb_43(fringeCommon_io_dram_3_wdata_bits_wstrb_43),
    .io_dram_3_wdata_bits_wstrb_44(fringeCommon_io_dram_3_wdata_bits_wstrb_44),
    .io_dram_3_wdata_bits_wstrb_45(fringeCommon_io_dram_3_wdata_bits_wstrb_45),
    .io_dram_3_wdata_bits_wstrb_46(fringeCommon_io_dram_3_wdata_bits_wstrb_46),
    .io_dram_3_wdata_bits_wstrb_47(fringeCommon_io_dram_3_wdata_bits_wstrb_47),
    .io_dram_3_wdata_bits_wstrb_48(fringeCommon_io_dram_3_wdata_bits_wstrb_48),
    .io_dram_3_wdata_bits_wstrb_49(fringeCommon_io_dram_3_wdata_bits_wstrb_49),
    .io_dram_3_wdata_bits_wstrb_50(fringeCommon_io_dram_3_wdata_bits_wstrb_50),
    .io_dram_3_wdata_bits_wstrb_51(fringeCommon_io_dram_3_wdata_bits_wstrb_51),
    .io_dram_3_wdata_bits_wstrb_52(fringeCommon_io_dram_3_wdata_bits_wstrb_52),
    .io_dram_3_wdata_bits_wstrb_53(fringeCommon_io_dram_3_wdata_bits_wstrb_53),
    .io_dram_3_wdata_bits_wstrb_54(fringeCommon_io_dram_3_wdata_bits_wstrb_54),
    .io_dram_3_wdata_bits_wstrb_55(fringeCommon_io_dram_3_wdata_bits_wstrb_55),
    .io_dram_3_wdata_bits_wstrb_56(fringeCommon_io_dram_3_wdata_bits_wstrb_56),
    .io_dram_3_wdata_bits_wstrb_57(fringeCommon_io_dram_3_wdata_bits_wstrb_57),
    .io_dram_3_wdata_bits_wstrb_58(fringeCommon_io_dram_3_wdata_bits_wstrb_58),
    .io_dram_3_wdata_bits_wstrb_59(fringeCommon_io_dram_3_wdata_bits_wstrb_59),
    .io_dram_3_wdata_bits_wstrb_60(fringeCommon_io_dram_3_wdata_bits_wstrb_60),
    .io_dram_3_wdata_bits_wstrb_61(fringeCommon_io_dram_3_wdata_bits_wstrb_61),
    .io_dram_3_wdata_bits_wstrb_62(fringeCommon_io_dram_3_wdata_bits_wstrb_62),
    .io_dram_3_wdata_bits_wstrb_63(fringeCommon_io_dram_3_wdata_bits_wstrb_63),
    .io_dram_3_wdata_bits_wlast(fringeCommon_io_dram_3_wdata_bits_wlast),
    .io_dram_3_rresp_ready(fringeCommon_io_dram_3_rresp_ready),
    .io_dram_3_wresp_ready(fringeCommon_io_dram_3_wresp_ready),
    .io_dram_3_wresp_valid(fringeCommon_io_dram_3_wresp_valid),
    .io_dram_3_wresp_bits_tag(fringeCommon_io_dram_3_wresp_bits_tag),
    .io_heap_0_req_valid(fringeCommon_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(fringeCommon_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(fringeCommon_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(fringeCommon_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(fringeCommon_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(fringeCommon_io_heap_0_resp_bits_sizeAddr)
  );
  AXI4LiteToRFBridge AXI4LiteToRFBridge ( // @[FringeZynq.scala 90:31:@143595.4]
    .clock(AXI4LiteToRFBridge_clock),
    .reset(AXI4LiteToRFBridge_reset),
    .io_S_AXI_AWADDR(AXI4LiteToRFBridge_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(AXI4LiteToRFBridge_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(AXI4LiteToRFBridge_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(AXI4LiteToRFBridge_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(AXI4LiteToRFBridge_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(AXI4LiteToRFBridge_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(AXI4LiteToRFBridge_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(AXI4LiteToRFBridge_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(AXI4LiteToRFBridge_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(AXI4LiteToRFBridge_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(AXI4LiteToRFBridge_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(AXI4LiteToRFBridge_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(AXI4LiteToRFBridge_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(AXI4LiteToRFBridge_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(AXI4LiteToRFBridge_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(AXI4LiteToRFBridge_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(AXI4LiteToRFBridge_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(AXI4LiteToRFBridge_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(AXI4LiteToRFBridge_io_S_AXI_BREADY),
    .io_raddr(AXI4LiteToRFBridge_io_raddr),
    .io_wen(AXI4LiteToRFBridge_io_wen),
    .io_waddr(AXI4LiteToRFBridge_io_waddr),
    .io_wdata(AXI4LiteToRFBridge_io_wdata),
    .io_rdata(AXI4LiteToRFBridge_io_rdata)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge ( // @[FringeZynq.scala 131:27:@143745.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_1 ( // @[FringeZynq.scala 131:27:@143901.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_1_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_1_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_1_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_1_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_1_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_1_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_1_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_1_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_1_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_1_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_1_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_1_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_1_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_1_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_1_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_1_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_1_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_1_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_1_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_1_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_1_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_1_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_1_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_1_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_1_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_1_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_1_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_1_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_1_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_1_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_1_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_1_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_2 ( // @[FringeZynq.scala 131:27:@144057.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_2_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_2_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_2_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_2_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_2_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_2_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_2_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_2_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_2_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_2_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_2_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_2_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_2_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_2_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_2_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_2_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_2_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_2_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_2_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_2_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_2_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_2_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_2_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_2_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_2_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_2_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_2_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_2_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_2_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_2_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_2_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_2_io_M_AXI_BREADY)
  );
  MAGToAXI4Bridge MAGToAXI4Bridge_3 ( // @[FringeZynq.scala 131:27:@144213.4]
    .io_in_cmd_ready(MAGToAXI4Bridge_3_io_in_cmd_ready),
    .io_in_cmd_valid(MAGToAXI4Bridge_3_io_in_cmd_valid),
    .io_in_cmd_bits_addr(MAGToAXI4Bridge_3_io_in_cmd_bits_addr),
    .io_in_cmd_bits_size(MAGToAXI4Bridge_3_io_in_cmd_bits_size),
    .io_in_cmd_bits_isWr(MAGToAXI4Bridge_3_io_in_cmd_bits_isWr),
    .io_in_cmd_bits_tag(MAGToAXI4Bridge_3_io_in_cmd_bits_tag),
    .io_in_wdata_ready(MAGToAXI4Bridge_3_io_in_wdata_ready),
    .io_in_wdata_valid(MAGToAXI4Bridge_3_io_in_wdata_valid),
    .io_in_wdata_bits_wdata_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0),
    .io_in_wdata_bits_wdata_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1),
    .io_in_wdata_bits_wdata_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2),
    .io_in_wdata_bits_wdata_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3),
    .io_in_wdata_bits_wdata_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4),
    .io_in_wdata_bits_wdata_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5),
    .io_in_wdata_bits_wdata_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6),
    .io_in_wdata_bits_wdata_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7),
    .io_in_wdata_bits_wdata_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8),
    .io_in_wdata_bits_wdata_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9),
    .io_in_wdata_bits_wdata_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10),
    .io_in_wdata_bits_wdata_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11),
    .io_in_wdata_bits_wdata_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12),
    .io_in_wdata_bits_wdata_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13),
    .io_in_wdata_bits_wdata_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14),
    .io_in_wdata_bits_wdata_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15),
    .io_in_wdata_bits_wstrb_0(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0),
    .io_in_wdata_bits_wstrb_1(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1),
    .io_in_wdata_bits_wstrb_2(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2),
    .io_in_wdata_bits_wstrb_3(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3),
    .io_in_wdata_bits_wstrb_4(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4),
    .io_in_wdata_bits_wstrb_5(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5),
    .io_in_wdata_bits_wstrb_6(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6),
    .io_in_wdata_bits_wstrb_7(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7),
    .io_in_wdata_bits_wstrb_8(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8),
    .io_in_wdata_bits_wstrb_9(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9),
    .io_in_wdata_bits_wstrb_10(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10),
    .io_in_wdata_bits_wstrb_11(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11),
    .io_in_wdata_bits_wstrb_12(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12),
    .io_in_wdata_bits_wstrb_13(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13),
    .io_in_wdata_bits_wstrb_14(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14),
    .io_in_wdata_bits_wstrb_15(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15),
    .io_in_wdata_bits_wstrb_16(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16),
    .io_in_wdata_bits_wstrb_17(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17),
    .io_in_wdata_bits_wstrb_18(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18),
    .io_in_wdata_bits_wstrb_19(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19),
    .io_in_wdata_bits_wstrb_20(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20),
    .io_in_wdata_bits_wstrb_21(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21),
    .io_in_wdata_bits_wstrb_22(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22),
    .io_in_wdata_bits_wstrb_23(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23),
    .io_in_wdata_bits_wstrb_24(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24),
    .io_in_wdata_bits_wstrb_25(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25),
    .io_in_wdata_bits_wstrb_26(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26),
    .io_in_wdata_bits_wstrb_27(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27),
    .io_in_wdata_bits_wstrb_28(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28),
    .io_in_wdata_bits_wstrb_29(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29),
    .io_in_wdata_bits_wstrb_30(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30),
    .io_in_wdata_bits_wstrb_31(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31),
    .io_in_wdata_bits_wstrb_32(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32),
    .io_in_wdata_bits_wstrb_33(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33),
    .io_in_wdata_bits_wstrb_34(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34),
    .io_in_wdata_bits_wstrb_35(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35),
    .io_in_wdata_bits_wstrb_36(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36),
    .io_in_wdata_bits_wstrb_37(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37),
    .io_in_wdata_bits_wstrb_38(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38),
    .io_in_wdata_bits_wstrb_39(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39),
    .io_in_wdata_bits_wstrb_40(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40),
    .io_in_wdata_bits_wstrb_41(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41),
    .io_in_wdata_bits_wstrb_42(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42),
    .io_in_wdata_bits_wstrb_43(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43),
    .io_in_wdata_bits_wstrb_44(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44),
    .io_in_wdata_bits_wstrb_45(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45),
    .io_in_wdata_bits_wstrb_46(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46),
    .io_in_wdata_bits_wstrb_47(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47),
    .io_in_wdata_bits_wstrb_48(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48),
    .io_in_wdata_bits_wstrb_49(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49),
    .io_in_wdata_bits_wstrb_50(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50),
    .io_in_wdata_bits_wstrb_51(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51),
    .io_in_wdata_bits_wstrb_52(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52),
    .io_in_wdata_bits_wstrb_53(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53),
    .io_in_wdata_bits_wstrb_54(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54),
    .io_in_wdata_bits_wstrb_55(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55),
    .io_in_wdata_bits_wstrb_56(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56),
    .io_in_wdata_bits_wstrb_57(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57),
    .io_in_wdata_bits_wstrb_58(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58),
    .io_in_wdata_bits_wstrb_59(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59),
    .io_in_wdata_bits_wstrb_60(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60),
    .io_in_wdata_bits_wstrb_61(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61),
    .io_in_wdata_bits_wstrb_62(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62),
    .io_in_wdata_bits_wstrb_63(MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63),
    .io_in_wdata_bits_wlast(MAGToAXI4Bridge_3_io_in_wdata_bits_wlast),
    .io_in_rresp_ready(MAGToAXI4Bridge_3_io_in_rresp_ready),
    .io_in_wresp_ready(MAGToAXI4Bridge_3_io_in_wresp_ready),
    .io_in_wresp_valid(MAGToAXI4Bridge_3_io_in_wresp_valid),
    .io_in_wresp_bits_tag(MAGToAXI4Bridge_3_io_in_wresp_bits_tag),
    .io_M_AXI_AWID(MAGToAXI4Bridge_3_io_M_AXI_AWID),
    .io_M_AXI_AWADDR(MAGToAXI4Bridge_3_io_M_AXI_AWADDR),
    .io_M_AXI_AWLEN(MAGToAXI4Bridge_3_io_M_AXI_AWLEN),
    .io_M_AXI_AWVALID(MAGToAXI4Bridge_3_io_M_AXI_AWVALID),
    .io_M_AXI_AWREADY(MAGToAXI4Bridge_3_io_M_AXI_AWREADY),
    .io_M_AXI_ARID(MAGToAXI4Bridge_3_io_M_AXI_ARID),
    .io_M_AXI_ARADDR(MAGToAXI4Bridge_3_io_M_AXI_ARADDR),
    .io_M_AXI_ARLEN(MAGToAXI4Bridge_3_io_M_AXI_ARLEN),
    .io_M_AXI_ARVALID(MAGToAXI4Bridge_3_io_M_AXI_ARVALID),
    .io_M_AXI_ARREADY(MAGToAXI4Bridge_3_io_M_AXI_ARREADY),
    .io_M_AXI_WDATA(MAGToAXI4Bridge_3_io_M_AXI_WDATA),
    .io_M_AXI_WSTRB(MAGToAXI4Bridge_3_io_M_AXI_WSTRB),
    .io_M_AXI_WLAST(MAGToAXI4Bridge_3_io_M_AXI_WLAST),
    .io_M_AXI_WVALID(MAGToAXI4Bridge_3_io_M_AXI_WVALID),
    .io_M_AXI_WREADY(MAGToAXI4Bridge_3_io_M_AXI_WREADY),
    .io_M_AXI_RREADY(MAGToAXI4Bridge_3_io_M_AXI_RREADY),
    .io_M_AXI_BID(MAGToAXI4Bridge_3_io_M_AXI_BID),
    .io_M_AXI_BVALID(MAGToAXI4Bridge_3_io_M_AXI_BVALID),
    .io_M_AXI_BREADY(MAGToAXI4Bridge_3_io_M_AXI_BREADY)
  );
  assign io_S_AXI_AWREADY = AXI4LiteToRFBridge_io_S_AXI_AWREADY; // @[FringeZynq.scala 91:28:@143613.4]
  assign io_S_AXI_ARREADY = AXI4LiteToRFBridge_io_S_AXI_ARREADY; // @[FringeZynq.scala 91:28:@143609.4]
  assign io_S_AXI_WREADY = AXI4LiteToRFBridge_io_S_AXI_WREADY; // @[FringeZynq.scala 91:28:@143605.4]
  assign io_S_AXI_RDATA = AXI4LiteToRFBridge_io_S_AXI_RDATA; // @[FringeZynq.scala 91:28:@143604.4]
  assign io_S_AXI_RRESP = AXI4LiteToRFBridge_io_S_AXI_RRESP; // @[FringeZynq.scala 91:28:@143603.4]
  assign io_S_AXI_RVALID = AXI4LiteToRFBridge_io_S_AXI_RVALID; // @[FringeZynq.scala 91:28:@143602.4]
  assign io_S_AXI_BRESP = AXI4LiteToRFBridge_io_S_AXI_BRESP; // @[FringeZynq.scala 91:28:@143600.4]
  assign io_S_AXI_BVALID = AXI4LiteToRFBridge_io_S_AXI_BVALID; // @[FringeZynq.scala 91:28:@143599.4]
  assign io_M_AXI_0_AWID = MAGToAXI4Bridge_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@143900.4]
  assign io_M_AXI_0_AWADDR = MAGToAXI4Bridge_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@143898.4]
  assign io_M_AXI_0_AWLEN = MAGToAXI4Bridge_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@143897.4]
  assign io_M_AXI_0_AWVALID = MAGToAXI4Bridge_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@143890.4]
  assign io_M_AXI_0_ARID = MAGToAXI4Bridge_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@143888.4]
  assign io_M_AXI_0_ARADDR = MAGToAXI4Bridge_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@143886.4]
  assign io_M_AXI_0_ARLEN = MAGToAXI4Bridge_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@143885.4]
  assign io_M_AXI_0_ARVALID = MAGToAXI4Bridge_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@143878.4]
  assign io_M_AXI_0_WDATA = MAGToAXI4Bridge_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@143876.4]
  assign io_M_AXI_0_WSTRB = MAGToAXI4Bridge_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@143875.4]
  assign io_M_AXI_0_WLAST = MAGToAXI4Bridge_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@143874.4]
  assign io_M_AXI_0_WVALID = MAGToAXI4Bridge_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@143873.4]
  assign io_M_AXI_0_RREADY = MAGToAXI4Bridge_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@143865.4]
  assign io_M_AXI_0_BREADY = MAGToAXI4Bridge_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@143860.4]
  assign io_M_AXI_1_AWID = MAGToAXI4Bridge_1_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@144056.4]
  assign io_M_AXI_1_AWADDR = MAGToAXI4Bridge_1_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@144054.4]
  assign io_M_AXI_1_AWLEN = MAGToAXI4Bridge_1_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@144053.4]
  assign io_M_AXI_1_AWVALID = MAGToAXI4Bridge_1_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@144046.4]
  assign io_M_AXI_1_ARID = MAGToAXI4Bridge_1_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@144044.4]
  assign io_M_AXI_1_ARADDR = MAGToAXI4Bridge_1_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@144042.4]
  assign io_M_AXI_1_ARLEN = MAGToAXI4Bridge_1_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@144041.4]
  assign io_M_AXI_1_ARVALID = MAGToAXI4Bridge_1_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@144034.4]
  assign io_M_AXI_1_WDATA = MAGToAXI4Bridge_1_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@144032.4]
  assign io_M_AXI_1_WSTRB = MAGToAXI4Bridge_1_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@144031.4]
  assign io_M_AXI_1_WLAST = MAGToAXI4Bridge_1_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@144030.4]
  assign io_M_AXI_1_WVALID = MAGToAXI4Bridge_1_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@144029.4]
  assign io_M_AXI_1_RREADY = MAGToAXI4Bridge_1_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@144021.4]
  assign io_M_AXI_1_BREADY = MAGToAXI4Bridge_1_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@144016.4]
  assign io_M_AXI_2_AWID = MAGToAXI4Bridge_2_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@144212.4]
  assign io_M_AXI_2_AWADDR = MAGToAXI4Bridge_2_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@144210.4]
  assign io_M_AXI_2_AWLEN = MAGToAXI4Bridge_2_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@144209.4]
  assign io_M_AXI_2_AWVALID = MAGToAXI4Bridge_2_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@144202.4]
  assign io_M_AXI_2_ARID = MAGToAXI4Bridge_2_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@144200.4]
  assign io_M_AXI_2_ARADDR = MAGToAXI4Bridge_2_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@144198.4]
  assign io_M_AXI_2_ARLEN = MAGToAXI4Bridge_2_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@144197.4]
  assign io_M_AXI_2_ARVALID = MAGToAXI4Bridge_2_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@144190.4]
  assign io_M_AXI_2_WDATA = MAGToAXI4Bridge_2_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@144188.4]
  assign io_M_AXI_2_WSTRB = MAGToAXI4Bridge_2_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@144187.4]
  assign io_M_AXI_2_WLAST = MAGToAXI4Bridge_2_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@144186.4]
  assign io_M_AXI_2_WVALID = MAGToAXI4Bridge_2_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@144185.4]
  assign io_M_AXI_2_RREADY = MAGToAXI4Bridge_2_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@144177.4]
  assign io_M_AXI_2_BREADY = MAGToAXI4Bridge_2_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@144172.4]
  assign io_M_AXI_3_AWID = MAGToAXI4Bridge_3_io_M_AXI_AWID; // @[FringeZynq.scala 133:10:@144368.4]
  assign io_M_AXI_3_AWADDR = MAGToAXI4Bridge_3_io_M_AXI_AWADDR; // @[FringeZynq.scala 133:10:@144366.4]
  assign io_M_AXI_3_AWLEN = MAGToAXI4Bridge_3_io_M_AXI_AWLEN; // @[FringeZynq.scala 133:10:@144365.4]
  assign io_M_AXI_3_AWVALID = MAGToAXI4Bridge_3_io_M_AXI_AWVALID; // @[FringeZynq.scala 133:10:@144358.4]
  assign io_M_AXI_3_ARID = MAGToAXI4Bridge_3_io_M_AXI_ARID; // @[FringeZynq.scala 133:10:@144356.4]
  assign io_M_AXI_3_ARADDR = MAGToAXI4Bridge_3_io_M_AXI_ARADDR; // @[FringeZynq.scala 133:10:@144354.4]
  assign io_M_AXI_3_ARLEN = MAGToAXI4Bridge_3_io_M_AXI_ARLEN; // @[FringeZynq.scala 133:10:@144353.4]
  assign io_M_AXI_3_ARVALID = MAGToAXI4Bridge_3_io_M_AXI_ARVALID; // @[FringeZynq.scala 133:10:@144346.4]
  assign io_M_AXI_3_WDATA = MAGToAXI4Bridge_3_io_M_AXI_WDATA; // @[FringeZynq.scala 133:10:@144344.4]
  assign io_M_AXI_3_WSTRB = MAGToAXI4Bridge_3_io_M_AXI_WSTRB; // @[FringeZynq.scala 133:10:@144343.4]
  assign io_M_AXI_3_WLAST = MAGToAXI4Bridge_3_io_M_AXI_WLAST; // @[FringeZynq.scala 133:10:@144342.4]
  assign io_M_AXI_3_WVALID = MAGToAXI4Bridge_3_io_M_AXI_WVALID; // @[FringeZynq.scala 133:10:@144341.4]
  assign io_M_AXI_3_RREADY = MAGToAXI4Bridge_3_io_M_AXI_RREADY; // @[FringeZynq.scala 133:10:@144333.4]
  assign io_M_AXI_3_BREADY = MAGToAXI4Bridge_3_io_M_AXI_BREADY; // @[FringeZynq.scala 133:10:@144328.4]
  assign io_enable = fringeCommon_io_enable; // @[FringeZynq.scala 115:13:@143623.4]
  assign io_reset = fringeCommon_io_reset; // @[FringeZynq.scala 119:12:@143627.4]
  assign io_argIns_0 = fringeCommon_io_argIns_0; // @[FringeZynq.scala 121:13:@143628.4]
  assign io_argIns_1 = fringeCommon_io_argIns_1; // @[FringeZynq.scala 121:13:@143629.4]
  assign io_memStreams_stores_0_cmd_ready = fringeCommon_io_memStreams_stores_0_cmd_ready; // @[FringeZynq.scala 126:17:@143716.4]
  assign io_memStreams_stores_0_data_ready = fringeCommon_io_memStreams_stores_0_data_ready; // @[FringeZynq.scala 126:17:@143712.4]
  assign io_memStreams_stores_0_wresp_valid = fringeCommon_io_memStreams_stores_0_wresp_valid; // @[FringeZynq.scala 126:17:@143707.4]
  assign io_memStreams_stores_0_wresp_bits = fringeCommon_io_memStreams_stores_0_wresp_bits; // @[FringeZynq.scala 126:17:@143706.4]
  assign io_heap_0_resp_valid = fringeCommon_io_heap_0_resp_valid; // @[FringeZynq.scala 127:11:@143741.4]
  assign io_heap_0_resp_bits_allocDealloc = fringeCommon_io_heap_0_resp_bits_allocDealloc; // @[FringeZynq.scala 127:11:@143740.4]
  assign io_heap_0_resp_bits_sizeAddr = fringeCommon_io_heap_0_resp_bits_sizeAddr; // @[FringeZynq.scala 127:11:@143739.4]
  assign fringeCommon_clock = clock; // @[:@142690.4]
  assign fringeCommon_reset = reset; // @[:@142691.4 FringeZynq.scala 117:22:@143626.4]
  assign fringeCommon_io_raddr = AXI4LiteToRFBridge_io_raddr; // @[FringeZynq.scala 94:27:@143617.4]
  assign fringeCommon_io_wen = AXI4LiteToRFBridge_io_wen; // @[FringeZynq.scala 95:27:@143618.4]
  assign fringeCommon_io_waddr = AXI4LiteToRFBridge_io_waddr; // @[FringeZynq.scala 96:27:@143619.4]
  assign fringeCommon_io_wdata = {{32'd0}, AXI4LiteToRFBridge_io_wdata}; // @[FringeZynq.scala 97:27:@143620.4]
  assign fringeCommon_io_done = io_done; // @[FringeZynq.scala 116:24:@143624.4]
  assign fringeCommon_io_argOuts_0_valid = io_argOuts_0_valid; // @[FringeZynq.scala 122:27:@143631.4]
  assign fringeCommon_io_argOuts_0_bits = io_argOuts_0_bits; // @[FringeZynq.scala 122:27:@143630.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_valid = io_memStreams_stores_0_cmd_valid; // @[FringeZynq.scala 126:17:@143715.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_addr = io_memStreams_stores_0_cmd_bits_addr; // @[FringeZynq.scala 126:17:@143714.4]
  assign fringeCommon_io_memStreams_stores_0_cmd_bits_size = io_memStreams_stores_0_cmd_bits_size; // @[FringeZynq.scala 126:17:@143713.4]
  assign fringeCommon_io_memStreams_stores_0_data_valid = io_memStreams_stores_0_data_valid; // @[FringeZynq.scala 126:17:@143711.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wdata_0 = io_memStreams_stores_0_data_bits_wdata_0; // @[FringeZynq.scala 126:17:@143710.4]
  assign fringeCommon_io_memStreams_stores_0_data_bits_wstrb = io_memStreams_stores_0_data_bits_wstrb; // @[FringeZynq.scala 126:17:@143709.4]
  assign fringeCommon_io_memStreams_stores_0_wresp_ready = io_memStreams_stores_0_wresp_ready; // @[FringeZynq.scala 126:17:@143708.4]
  assign fringeCommon_io_dram_0_cmd_ready = MAGToAXI4Bridge_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@143859.4]
  assign fringeCommon_io_dram_0_wdata_ready = MAGToAXI4Bridge_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@143852.4]
  assign fringeCommon_io_dram_0_wresp_valid = MAGToAXI4Bridge_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@143749.4]
  assign fringeCommon_io_dram_0_wresp_bits_tag = MAGToAXI4Bridge_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@143748.4]
  assign fringeCommon_io_dram_1_cmd_ready = MAGToAXI4Bridge_1_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@144015.4]
  assign fringeCommon_io_dram_1_wdata_ready = MAGToAXI4Bridge_1_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@144008.4]
  assign fringeCommon_io_dram_1_wresp_valid = MAGToAXI4Bridge_1_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@143905.4]
  assign fringeCommon_io_dram_1_wresp_bits_tag = MAGToAXI4Bridge_1_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@143904.4]
  assign fringeCommon_io_dram_2_cmd_ready = MAGToAXI4Bridge_2_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@144171.4]
  assign fringeCommon_io_dram_2_wdata_ready = MAGToAXI4Bridge_2_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@144164.4]
  assign fringeCommon_io_dram_2_wresp_valid = MAGToAXI4Bridge_2_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@144061.4]
  assign fringeCommon_io_dram_2_wresp_bits_tag = MAGToAXI4Bridge_2_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@144060.4]
  assign fringeCommon_io_dram_3_cmd_ready = MAGToAXI4Bridge_3_io_in_cmd_ready; // @[FringeZynq.scala 132:21:@144327.4]
  assign fringeCommon_io_dram_3_wdata_ready = MAGToAXI4Bridge_3_io_in_wdata_ready; // @[FringeZynq.scala 132:21:@144320.4]
  assign fringeCommon_io_dram_3_wresp_valid = MAGToAXI4Bridge_3_io_in_wresp_valid; // @[FringeZynq.scala 132:21:@144217.4]
  assign fringeCommon_io_dram_3_wresp_bits_tag = MAGToAXI4Bridge_3_io_in_wresp_bits_tag; // @[FringeZynq.scala 132:21:@144216.4]
  assign fringeCommon_io_heap_0_req_valid = io_heap_0_req_valid; // @[FringeZynq.scala 127:11:@143744.4]
  assign fringeCommon_io_heap_0_req_bits_allocDealloc = io_heap_0_req_bits_allocDealloc; // @[FringeZynq.scala 127:11:@143743.4]
  assign fringeCommon_io_heap_0_req_bits_sizeAddr = io_heap_0_req_bits_sizeAddr; // @[FringeZynq.scala 127:11:@143742.4]
  assign AXI4LiteToRFBridge_clock = clock; // @[:@143596.4]
  assign AXI4LiteToRFBridge_reset = reset; // @[:@143597.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[FringeZynq.scala 91:28:@143616.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[FringeZynq.scala 91:28:@143615.4]
  assign AXI4LiteToRFBridge_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[FringeZynq.scala 91:28:@143614.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[FringeZynq.scala 91:28:@143612.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[FringeZynq.scala 91:28:@143611.4]
  assign AXI4LiteToRFBridge_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[FringeZynq.scala 91:28:@143610.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[FringeZynq.scala 91:28:@143608.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[FringeZynq.scala 91:28:@143607.4]
  assign AXI4LiteToRFBridge_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[FringeZynq.scala 91:28:@143606.4]
  assign AXI4LiteToRFBridge_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[FringeZynq.scala 91:28:@143601.4]
  assign AXI4LiteToRFBridge_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[FringeZynq.scala 91:28:@143598.4]
  assign AXI4LiteToRFBridge_io_rdata = fringeCommon_io_rdata[31:0]; // @[FringeZynq.scala 98:28:@143621.4]
  assign MAGToAXI4Bridge_io_in_cmd_valid = fringeCommon_io_dram_0_cmd_valid; // @[FringeZynq.scala 132:21:@143858.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_addr = fringeCommon_io_dram_0_cmd_bits_addr; // @[FringeZynq.scala 132:21:@143857.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_size = fringeCommon_io_dram_0_cmd_bits_size; // @[FringeZynq.scala 132:21:@143856.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_isWr = fringeCommon_io_dram_0_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@143854.4]
  assign MAGToAXI4Bridge_io_in_cmd_bits_tag = fringeCommon_io_dram_0_cmd_bits_tag; // @[FringeZynq.scala 132:21:@143853.4]
  assign MAGToAXI4Bridge_io_in_wdata_valid = fringeCommon_io_dram_0_wdata_valid; // @[FringeZynq.scala 132:21:@143851.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_0_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@143835.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_0_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@143836.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_0_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@143837.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_0_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@143838.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_0_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@143839.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_0_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@143840.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_0_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@143841.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_0_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@143842.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_0_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@143843.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_0_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@143844.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_0_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@143845.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_0_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@143846.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_0_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@143847.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_0_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@143848.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_0_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@143849.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_0_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@143850.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_0_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@143771.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_0_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@143772.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_0_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@143773.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_0_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@143774.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_0_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@143775.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_0_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@143776.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_0_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@143777.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_0_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@143778.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_0_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@143779.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_0_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@143780.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_0_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@143781.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_0_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@143782.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_0_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@143783.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_0_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@143784.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_0_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@143785.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_0_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@143786.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_0_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@143787.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_0_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@143788.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_0_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@143789.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_0_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@143790.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_0_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@143791.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_0_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@143792.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_0_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@143793.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_0_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@143794.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_0_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@143795.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_0_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@143796.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_0_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@143797.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_0_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@143798.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_0_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@143799.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_0_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@143800.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_0_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@143801.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_0_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@143802.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_0_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@143803.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_0_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@143804.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_0_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@143805.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_0_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@143806.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_0_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@143807.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_0_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@143808.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_0_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@143809.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_0_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@143810.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_0_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@143811.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_0_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@143812.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_0_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@143813.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_0_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@143814.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_0_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@143815.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_0_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@143816.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_0_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@143817.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_0_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@143818.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_0_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@143819.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_0_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@143820.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_0_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@143821.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_0_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@143822.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_0_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@143823.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_0_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@143824.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_0_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@143825.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_0_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@143826.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_0_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@143827.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_0_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@143828.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_0_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@143829.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_0_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@143830.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_0_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@143831.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_0_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@143832.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_0_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@143833.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_0_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@143834.4]
  assign MAGToAXI4Bridge_io_in_wdata_bits_wlast = fringeCommon_io_dram_0_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@143770.4]
  assign MAGToAXI4Bridge_io_in_rresp_ready = fringeCommon_io_dram_0_rresp_ready; // @[FringeZynq.scala 132:21:@143769.4]
  assign MAGToAXI4Bridge_io_in_wresp_ready = fringeCommon_io_dram_0_wresp_ready; // @[FringeZynq.scala 132:21:@143750.4]
  assign MAGToAXI4Bridge_io_M_AXI_AWREADY = io_M_AXI_0_AWREADY; // @[FringeZynq.scala 133:10:@143889.4]
  assign MAGToAXI4Bridge_io_M_AXI_ARREADY = io_M_AXI_0_ARREADY; // @[FringeZynq.scala 133:10:@143877.4]
  assign MAGToAXI4Bridge_io_M_AXI_WREADY = io_M_AXI_0_WREADY; // @[FringeZynq.scala 133:10:@143872.4]
  assign MAGToAXI4Bridge_io_M_AXI_BID = io_M_AXI_0_BID; // @[FringeZynq.scala 133:10:@143864.4]
  assign MAGToAXI4Bridge_io_M_AXI_BVALID = io_M_AXI_0_BVALID; // @[FringeZynq.scala 133:10:@143861.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_valid = fringeCommon_io_dram_1_cmd_valid; // @[FringeZynq.scala 132:21:@144014.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_addr = fringeCommon_io_dram_1_cmd_bits_addr; // @[FringeZynq.scala 132:21:@144013.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_size = fringeCommon_io_dram_1_cmd_bits_size; // @[FringeZynq.scala 132:21:@144012.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_isWr = fringeCommon_io_dram_1_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@144010.4]
  assign MAGToAXI4Bridge_1_io_in_cmd_bits_tag = fringeCommon_io_dram_1_cmd_bits_tag; // @[FringeZynq.scala 132:21:@144009.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_valid = fringeCommon_io_dram_1_wdata_valid; // @[FringeZynq.scala 132:21:@144007.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_1_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@143991.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_1_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@143992.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_1_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@143993.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_1_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@143994.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_1_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@143995.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_1_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@143996.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_1_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@143997.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_1_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@143998.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_1_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@143999.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_1_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@144000.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_1_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@144001.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_1_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@144002.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_1_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@144003.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_1_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@144004.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_1_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@144005.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_1_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@144006.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_1_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@143927.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_1_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@143928.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_1_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@143929.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_1_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@143930.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_1_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@143931.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_1_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@143932.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_1_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@143933.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_1_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@143934.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_1_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@143935.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_1_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@143936.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_1_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@143937.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_1_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@143938.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_1_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@143939.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_1_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@143940.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_1_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@143941.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_1_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@143942.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_1_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@143943.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_1_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@143944.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_1_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@143945.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_1_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@143946.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_1_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@143947.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_1_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@143948.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_1_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@143949.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_1_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@143950.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_1_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@143951.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_1_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@143952.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_1_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@143953.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_1_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@143954.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_1_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@143955.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_1_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@143956.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_1_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@143957.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_1_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@143958.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_1_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@143959.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_1_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@143960.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_1_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@143961.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_1_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@143962.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_1_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@143963.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_1_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@143964.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_1_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@143965.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_1_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@143966.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_1_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@143967.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_1_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@143968.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_1_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@143969.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_1_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@143970.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_1_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@143971.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_1_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@143972.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_1_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@143973.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_1_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@143974.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_1_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@143975.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_1_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@143976.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_1_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@143977.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_1_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@143978.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_1_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@143979.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_1_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@143980.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_1_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@143981.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_1_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@143982.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_1_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@143983.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_1_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@143984.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_1_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@143985.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_1_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@143986.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_1_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@143987.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_1_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@143988.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_1_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@143989.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_1_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@143990.4]
  assign MAGToAXI4Bridge_1_io_in_wdata_bits_wlast = fringeCommon_io_dram_1_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@143926.4]
  assign MAGToAXI4Bridge_1_io_in_rresp_ready = fringeCommon_io_dram_1_rresp_ready; // @[FringeZynq.scala 132:21:@143925.4]
  assign MAGToAXI4Bridge_1_io_in_wresp_ready = fringeCommon_io_dram_1_wresp_ready; // @[FringeZynq.scala 132:21:@143906.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_AWREADY = io_M_AXI_1_AWREADY; // @[FringeZynq.scala 133:10:@144045.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_ARREADY = io_M_AXI_1_ARREADY; // @[FringeZynq.scala 133:10:@144033.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_WREADY = io_M_AXI_1_WREADY; // @[FringeZynq.scala 133:10:@144028.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BID = io_M_AXI_1_BID; // @[FringeZynq.scala 133:10:@144020.4]
  assign MAGToAXI4Bridge_1_io_M_AXI_BVALID = io_M_AXI_1_BVALID; // @[FringeZynq.scala 133:10:@144017.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_valid = fringeCommon_io_dram_2_cmd_valid; // @[FringeZynq.scala 132:21:@144170.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_addr = fringeCommon_io_dram_2_cmd_bits_addr; // @[FringeZynq.scala 132:21:@144169.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_size = fringeCommon_io_dram_2_cmd_bits_size; // @[FringeZynq.scala 132:21:@144168.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_isWr = fringeCommon_io_dram_2_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@144166.4]
  assign MAGToAXI4Bridge_2_io_in_cmd_bits_tag = fringeCommon_io_dram_2_cmd_bits_tag; // @[FringeZynq.scala 132:21:@144165.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_valid = fringeCommon_io_dram_2_wdata_valid; // @[FringeZynq.scala 132:21:@144163.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_2_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@144147.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_2_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@144148.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_2_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@144149.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_2_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@144150.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_2_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@144151.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_2_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@144152.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_2_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@144153.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_2_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@144154.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_2_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@144155.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_2_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@144156.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_2_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@144157.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_2_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@144158.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_2_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@144159.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_2_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@144160.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_2_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@144161.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_2_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@144162.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_2_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@144083.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_2_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@144084.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_2_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@144085.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_2_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@144086.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_2_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@144087.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_2_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@144088.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_2_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@144089.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_2_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@144090.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_2_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@144091.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_2_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@144092.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_2_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@144093.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_2_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@144094.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_2_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@144095.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_2_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@144096.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_2_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@144097.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_2_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@144098.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_2_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@144099.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_2_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@144100.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_2_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@144101.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_2_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@144102.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_2_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@144103.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_2_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@144104.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_2_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@144105.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_2_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@144106.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_2_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@144107.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_2_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@144108.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_2_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@144109.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_2_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@144110.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_2_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@144111.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_2_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@144112.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_2_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@144113.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_2_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@144114.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_2_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@144115.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_2_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@144116.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_2_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@144117.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_2_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@144118.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_2_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@144119.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_2_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@144120.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_2_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@144121.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_2_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@144122.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_2_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@144123.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_2_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@144124.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_2_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@144125.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_2_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@144126.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_2_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@144127.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_2_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@144128.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_2_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@144129.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_2_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@144130.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_2_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@144131.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_2_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@144132.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_2_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@144133.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_2_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@144134.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_2_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@144135.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_2_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@144136.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_2_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@144137.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_2_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@144138.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_2_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@144139.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_2_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@144140.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_2_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@144141.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_2_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@144142.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_2_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@144143.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_2_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@144144.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_2_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@144145.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_2_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@144146.4]
  assign MAGToAXI4Bridge_2_io_in_wdata_bits_wlast = fringeCommon_io_dram_2_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@144082.4]
  assign MAGToAXI4Bridge_2_io_in_rresp_ready = fringeCommon_io_dram_2_rresp_ready; // @[FringeZynq.scala 132:21:@144081.4]
  assign MAGToAXI4Bridge_2_io_in_wresp_ready = fringeCommon_io_dram_2_wresp_ready; // @[FringeZynq.scala 132:21:@144062.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_AWREADY = io_M_AXI_2_AWREADY; // @[FringeZynq.scala 133:10:@144201.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_ARREADY = io_M_AXI_2_ARREADY; // @[FringeZynq.scala 133:10:@144189.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_WREADY = io_M_AXI_2_WREADY; // @[FringeZynq.scala 133:10:@144184.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BID = io_M_AXI_2_BID; // @[FringeZynq.scala 133:10:@144176.4]
  assign MAGToAXI4Bridge_2_io_M_AXI_BVALID = io_M_AXI_2_BVALID; // @[FringeZynq.scala 133:10:@144173.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_valid = fringeCommon_io_dram_3_cmd_valid; // @[FringeZynq.scala 132:21:@144326.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_addr = fringeCommon_io_dram_3_cmd_bits_addr; // @[FringeZynq.scala 132:21:@144325.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_size = fringeCommon_io_dram_3_cmd_bits_size; // @[FringeZynq.scala 132:21:@144324.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_isWr = fringeCommon_io_dram_3_cmd_bits_isWr; // @[FringeZynq.scala 132:21:@144322.4]
  assign MAGToAXI4Bridge_3_io_in_cmd_bits_tag = fringeCommon_io_dram_3_cmd_bits_tag; // @[FringeZynq.scala 132:21:@144321.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_valid = fringeCommon_io_dram_3_wdata_valid; // @[FringeZynq.scala 132:21:@144319.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_0 = fringeCommon_io_dram_3_wdata_bits_wdata_0; // @[FringeZynq.scala 132:21:@144303.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_1 = fringeCommon_io_dram_3_wdata_bits_wdata_1; // @[FringeZynq.scala 132:21:@144304.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_2 = fringeCommon_io_dram_3_wdata_bits_wdata_2; // @[FringeZynq.scala 132:21:@144305.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_3 = fringeCommon_io_dram_3_wdata_bits_wdata_3; // @[FringeZynq.scala 132:21:@144306.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_4 = fringeCommon_io_dram_3_wdata_bits_wdata_4; // @[FringeZynq.scala 132:21:@144307.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_5 = fringeCommon_io_dram_3_wdata_bits_wdata_5; // @[FringeZynq.scala 132:21:@144308.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_6 = fringeCommon_io_dram_3_wdata_bits_wdata_6; // @[FringeZynq.scala 132:21:@144309.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_7 = fringeCommon_io_dram_3_wdata_bits_wdata_7; // @[FringeZynq.scala 132:21:@144310.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_8 = fringeCommon_io_dram_3_wdata_bits_wdata_8; // @[FringeZynq.scala 132:21:@144311.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_9 = fringeCommon_io_dram_3_wdata_bits_wdata_9; // @[FringeZynq.scala 132:21:@144312.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_10 = fringeCommon_io_dram_3_wdata_bits_wdata_10; // @[FringeZynq.scala 132:21:@144313.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_11 = fringeCommon_io_dram_3_wdata_bits_wdata_11; // @[FringeZynq.scala 132:21:@144314.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_12 = fringeCommon_io_dram_3_wdata_bits_wdata_12; // @[FringeZynq.scala 132:21:@144315.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_13 = fringeCommon_io_dram_3_wdata_bits_wdata_13; // @[FringeZynq.scala 132:21:@144316.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_14 = fringeCommon_io_dram_3_wdata_bits_wdata_14; // @[FringeZynq.scala 132:21:@144317.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wdata_15 = fringeCommon_io_dram_3_wdata_bits_wdata_15; // @[FringeZynq.scala 132:21:@144318.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_0 = fringeCommon_io_dram_3_wdata_bits_wstrb_0; // @[FringeZynq.scala 132:21:@144239.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_1 = fringeCommon_io_dram_3_wdata_bits_wstrb_1; // @[FringeZynq.scala 132:21:@144240.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_2 = fringeCommon_io_dram_3_wdata_bits_wstrb_2; // @[FringeZynq.scala 132:21:@144241.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_3 = fringeCommon_io_dram_3_wdata_bits_wstrb_3; // @[FringeZynq.scala 132:21:@144242.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_4 = fringeCommon_io_dram_3_wdata_bits_wstrb_4; // @[FringeZynq.scala 132:21:@144243.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_5 = fringeCommon_io_dram_3_wdata_bits_wstrb_5; // @[FringeZynq.scala 132:21:@144244.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_6 = fringeCommon_io_dram_3_wdata_bits_wstrb_6; // @[FringeZynq.scala 132:21:@144245.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_7 = fringeCommon_io_dram_3_wdata_bits_wstrb_7; // @[FringeZynq.scala 132:21:@144246.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_8 = fringeCommon_io_dram_3_wdata_bits_wstrb_8; // @[FringeZynq.scala 132:21:@144247.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_9 = fringeCommon_io_dram_3_wdata_bits_wstrb_9; // @[FringeZynq.scala 132:21:@144248.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_10 = fringeCommon_io_dram_3_wdata_bits_wstrb_10; // @[FringeZynq.scala 132:21:@144249.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_11 = fringeCommon_io_dram_3_wdata_bits_wstrb_11; // @[FringeZynq.scala 132:21:@144250.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_12 = fringeCommon_io_dram_3_wdata_bits_wstrb_12; // @[FringeZynq.scala 132:21:@144251.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_13 = fringeCommon_io_dram_3_wdata_bits_wstrb_13; // @[FringeZynq.scala 132:21:@144252.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_14 = fringeCommon_io_dram_3_wdata_bits_wstrb_14; // @[FringeZynq.scala 132:21:@144253.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_15 = fringeCommon_io_dram_3_wdata_bits_wstrb_15; // @[FringeZynq.scala 132:21:@144254.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_16 = fringeCommon_io_dram_3_wdata_bits_wstrb_16; // @[FringeZynq.scala 132:21:@144255.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_17 = fringeCommon_io_dram_3_wdata_bits_wstrb_17; // @[FringeZynq.scala 132:21:@144256.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_18 = fringeCommon_io_dram_3_wdata_bits_wstrb_18; // @[FringeZynq.scala 132:21:@144257.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_19 = fringeCommon_io_dram_3_wdata_bits_wstrb_19; // @[FringeZynq.scala 132:21:@144258.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_20 = fringeCommon_io_dram_3_wdata_bits_wstrb_20; // @[FringeZynq.scala 132:21:@144259.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_21 = fringeCommon_io_dram_3_wdata_bits_wstrb_21; // @[FringeZynq.scala 132:21:@144260.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_22 = fringeCommon_io_dram_3_wdata_bits_wstrb_22; // @[FringeZynq.scala 132:21:@144261.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_23 = fringeCommon_io_dram_3_wdata_bits_wstrb_23; // @[FringeZynq.scala 132:21:@144262.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_24 = fringeCommon_io_dram_3_wdata_bits_wstrb_24; // @[FringeZynq.scala 132:21:@144263.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_25 = fringeCommon_io_dram_3_wdata_bits_wstrb_25; // @[FringeZynq.scala 132:21:@144264.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_26 = fringeCommon_io_dram_3_wdata_bits_wstrb_26; // @[FringeZynq.scala 132:21:@144265.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_27 = fringeCommon_io_dram_3_wdata_bits_wstrb_27; // @[FringeZynq.scala 132:21:@144266.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_28 = fringeCommon_io_dram_3_wdata_bits_wstrb_28; // @[FringeZynq.scala 132:21:@144267.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_29 = fringeCommon_io_dram_3_wdata_bits_wstrb_29; // @[FringeZynq.scala 132:21:@144268.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_30 = fringeCommon_io_dram_3_wdata_bits_wstrb_30; // @[FringeZynq.scala 132:21:@144269.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_31 = fringeCommon_io_dram_3_wdata_bits_wstrb_31; // @[FringeZynq.scala 132:21:@144270.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_32 = fringeCommon_io_dram_3_wdata_bits_wstrb_32; // @[FringeZynq.scala 132:21:@144271.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_33 = fringeCommon_io_dram_3_wdata_bits_wstrb_33; // @[FringeZynq.scala 132:21:@144272.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_34 = fringeCommon_io_dram_3_wdata_bits_wstrb_34; // @[FringeZynq.scala 132:21:@144273.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_35 = fringeCommon_io_dram_3_wdata_bits_wstrb_35; // @[FringeZynq.scala 132:21:@144274.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_36 = fringeCommon_io_dram_3_wdata_bits_wstrb_36; // @[FringeZynq.scala 132:21:@144275.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_37 = fringeCommon_io_dram_3_wdata_bits_wstrb_37; // @[FringeZynq.scala 132:21:@144276.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_38 = fringeCommon_io_dram_3_wdata_bits_wstrb_38; // @[FringeZynq.scala 132:21:@144277.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_39 = fringeCommon_io_dram_3_wdata_bits_wstrb_39; // @[FringeZynq.scala 132:21:@144278.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_40 = fringeCommon_io_dram_3_wdata_bits_wstrb_40; // @[FringeZynq.scala 132:21:@144279.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_41 = fringeCommon_io_dram_3_wdata_bits_wstrb_41; // @[FringeZynq.scala 132:21:@144280.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_42 = fringeCommon_io_dram_3_wdata_bits_wstrb_42; // @[FringeZynq.scala 132:21:@144281.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_43 = fringeCommon_io_dram_3_wdata_bits_wstrb_43; // @[FringeZynq.scala 132:21:@144282.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_44 = fringeCommon_io_dram_3_wdata_bits_wstrb_44; // @[FringeZynq.scala 132:21:@144283.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_45 = fringeCommon_io_dram_3_wdata_bits_wstrb_45; // @[FringeZynq.scala 132:21:@144284.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_46 = fringeCommon_io_dram_3_wdata_bits_wstrb_46; // @[FringeZynq.scala 132:21:@144285.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_47 = fringeCommon_io_dram_3_wdata_bits_wstrb_47; // @[FringeZynq.scala 132:21:@144286.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_48 = fringeCommon_io_dram_3_wdata_bits_wstrb_48; // @[FringeZynq.scala 132:21:@144287.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_49 = fringeCommon_io_dram_3_wdata_bits_wstrb_49; // @[FringeZynq.scala 132:21:@144288.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_50 = fringeCommon_io_dram_3_wdata_bits_wstrb_50; // @[FringeZynq.scala 132:21:@144289.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_51 = fringeCommon_io_dram_3_wdata_bits_wstrb_51; // @[FringeZynq.scala 132:21:@144290.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_52 = fringeCommon_io_dram_3_wdata_bits_wstrb_52; // @[FringeZynq.scala 132:21:@144291.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_53 = fringeCommon_io_dram_3_wdata_bits_wstrb_53; // @[FringeZynq.scala 132:21:@144292.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_54 = fringeCommon_io_dram_3_wdata_bits_wstrb_54; // @[FringeZynq.scala 132:21:@144293.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_55 = fringeCommon_io_dram_3_wdata_bits_wstrb_55; // @[FringeZynq.scala 132:21:@144294.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_56 = fringeCommon_io_dram_3_wdata_bits_wstrb_56; // @[FringeZynq.scala 132:21:@144295.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_57 = fringeCommon_io_dram_3_wdata_bits_wstrb_57; // @[FringeZynq.scala 132:21:@144296.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_58 = fringeCommon_io_dram_3_wdata_bits_wstrb_58; // @[FringeZynq.scala 132:21:@144297.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_59 = fringeCommon_io_dram_3_wdata_bits_wstrb_59; // @[FringeZynq.scala 132:21:@144298.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_60 = fringeCommon_io_dram_3_wdata_bits_wstrb_60; // @[FringeZynq.scala 132:21:@144299.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_61 = fringeCommon_io_dram_3_wdata_bits_wstrb_61; // @[FringeZynq.scala 132:21:@144300.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_62 = fringeCommon_io_dram_3_wdata_bits_wstrb_62; // @[FringeZynq.scala 132:21:@144301.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wstrb_63 = fringeCommon_io_dram_3_wdata_bits_wstrb_63; // @[FringeZynq.scala 132:21:@144302.4]
  assign MAGToAXI4Bridge_3_io_in_wdata_bits_wlast = fringeCommon_io_dram_3_wdata_bits_wlast; // @[FringeZynq.scala 132:21:@144238.4]
  assign MAGToAXI4Bridge_3_io_in_rresp_ready = fringeCommon_io_dram_3_rresp_ready; // @[FringeZynq.scala 132:21:@144237.4]
  assign MAGToAXI4Bridge_3_io_in_wresp_ready = fringeCommon_io_dram_3_wresp_ready; // @[FringeZynq.scala 132:21:@144218.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_AWREADY = io_M_AXI_3_AWREADY; // @[FringeZynq.scala 133:10:@144357.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_ARREADY = io_M_AXI_3_ARREADY; // @[FringeZynq.scala 133:10:@144345.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_WREADY = io_M_AXI_3_WREADY; // @[FringeZynq.scala 133:10:@144340.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BID = io_M_AXI_3_BID; // @[FringeZynq.scala 133:10:@144332.4]
  assign MAGToAXI4Bridge_3_io_M_AXI_BVALID = io_M_AXI_3_BVALID; // @[FringeZynq.scala 133:10:@144329.4]
endmodule
module SpatialIP( // @[:@144370.2]
  input          clock, // @[:@144371.4]
  input          reset, // @[:@144372.4]
  input          io_raddr, // @[:@144373.4]
  input          io_wen, // @[:@144373.4]
  input          io_waddr, // @[:@144373.4]
  input          io_wdata, // @[:@144373.4]
  output         io_rdata, // @[:@144373.4]
  input  [31:0]  io_S_AXI_AWADDR, // @[:@144373.4]
  input  [2:0]   io_S_AXI_AWPROT, // @[:@144373.4]
  input          io_S_AXI_AWVALID, // @[:@144373.4]
  output         io_S_AXI_AWREADY, // @[:@144373.4]
  input  [31:0]  io_S_AXI_ARADDR, // @[:@144373.4]
  input  [2:0]   io_S_AXI_ARPROT, // @[:@144373.4]
  input          io_S_AXI_ARVALID, // @[:@144373.4]
  output         io_S_AXI_ARREADY, // @[:@144373.4]
  input  [31:0]  io_S_AXI_WDATA, // @[:@144373.4]
  input  [3:0]   io_S_AXI_WSTRB, // @[:@144373.4]
  input          io_S_AXI_WVALID, // @[:@144373.4]
  output         io_S_AXI_WREADY, // @[:@144373.4]
  output [31:0]  io_S_AXI_RDATA, // @[:@144373.4]
  output [1:0]   io_S_AXI_RRESP, // @[:@144373.4]
  output         io_S_AXI_RVALID, // @[:@144373.4]
  input          io_S_AXI_RREADY, // @[:@144373.4]
  output [1:0]   io_S_AXI_BRESP, // @[:@144373.4]
  output         io_S_AXI_BVALID, // @[:@144373.4]
  input          io_S_AXI_BREADY, // @[:@144373.4]
  output [31:0]  io_M_AXI_0_AWID, // @[:@144373.4]
  output [31:0]  io_M_AXI_0_AWUSER, // @[:@144373.4]
  output [31:0]  io_M_AXI_0_AWADDR, // @[:@144373.4]
  output [7:0]   io_M_AXI_0_AWLEN, // @[:@144373.4]
  output [2:0]   io_M_AXI_0_AWSIZE, // @[:@144373.4]
  output [1:0]   io_M_AXI_0_AWBURST, // @[:@144373.4]
  output         io_M_AXI_0_AWLOCK, // @[:@144373.4]
  output [3:0]   io_M_AXI_0_AWCACHE, // @[:@144373.4]
  output [2:0]   io_M_AXI_0_AWPROT, // @[:@144373.4]
  output [3:0]   io_M_AXI_0_AWQOS, // @[:@144373.4]
  output         io_M_AXI_0_AWVALID, // @[:@144373.4]
  input          io_M_AXI_0_AWREADY, // @[:@144373.4]
  output [31:0]  io_M_AXI_0_ARID, // @[:@144373.4]
  output [31:0]  io_M_AXI_0_ARUSER, // @[:@144373.4]
  output [31:0]  io_M_AXI_0_ARADDR, // @[:@144373.4]
  output [7:0]   io_M_AXI_0_ARLEN, // @[:@144373.4]
  output [2:0]   io_M_AXI_0_ARSIZE, // @[:@144373.4]
  output [1:0]   io_M_AXI_0_ARBURST, // @[:@144373.4]
  output         io_M_AXI_0_ARLOCK, // @[:@144373.4]
  output [3:0]   io_M_AXI_0_ARCACHE, // @[:@144373.4]
  output [2:0]   io_M_AXI_0_ARPROT, // @[:@144373.4]
  output [3:0]   io_M_AXI_0_ARQOS, // @[:@144373.4]
  output         io_M_AXI_0_ARVALID, // @[:@144373.4]
  input          io_M_AXI_0_ARREADY, // @[:@144373.4]
  output [511:0] io_M_AXI_0_WDATA, // @[:@144373.4]
  output [63:0]  io_M_AXI_0_WSTRB, // @[:@144373.4]
  output         io_M_AXI_0_WLAST, // @[:@144373.4]
  output         io_M_AXI_0_WVALID, // @[:@144373.4]
  input          io_M_AXI_0_WREADY, // @[:@144373.4]
  input  [31:0]  io_M_AXI_0_RID, // @[:@144373.4]
  input  [31:0]  io_M_AXI_0_RUSER, // @[:@144373.4]
  input  [511:0] io_M_AXI_0_RDATA, // @[:@144373.4]
  input  [1:0]   io_M_AXI_0_RRESP, // @[:@144373.4]
  input          io_M_AXI_0_RLAST, // @[:@144373.4]
  input          io_M_AXI_0_RVALID, // @[:@144373.4]
  output         io_M_AXI_0_RREADY, // @[:@144373.4]
  input  [31:0]  io_M_AXI_0_BID, // @[:@144373.4]
  input  [31:0]  io_M_AXI_0_BUSER, // @[:@144373.4]
  input  [1:0]   io_M_AXI_0_BRESP, // @[:@144373.4]
  input          io_M_AXI_0_BVALID, // @[:@144373.4]
  output         io_M_AXI_0_BREADY, // @[:@144373.4]
  output [31:0]  io_M_AXI_1_AWID, // @[:@144373.4]
  output [31:0]  io_M_AXI_1_AWUSER, // @[:@144373.4]
  output [31:0]  io_M_AXI_1_AWADDR, // @[:@144373.4]
  output [7:0]   io_M_AXI_1_AWLEN, // @[:@144373.4]
  output [2:0]   io_M_AXI_1_AWSIZE, // @[:@144373.4]
  output [1:0]   io_M_AXI_1_AWBURST, // @[:@144373.4]
  output         io_M_AXI_1_AWLOCK, // @[:@144373.4]
  output [3:0]   io_M_AXI_1_AWCACHE, // @[:@144373.4]
  output [2:0]   io_M_AXI_1_AWPROT, // @[:@144373.4]
  output [3:0]   io_M_AXI_1_AWQOS, // @[:@144373.4]
  output         io_M_AXI_1_AWVALID, // @[:@144373.4]
  input          io_M_AXI_1_AWREADY, // @[:@144373.4]
  output [31:0]  io_M_AXI_1_ARID, // @[:@144373.4]
  output [31:0]  io_M_AXI_1_ARUSER, // @[:@144373.4]
  output [31:0]  io_M_AXI_1_ARADDR, // @[:@144373.4]
  output [7:0]   io_M_AXI_1_ARLEN, // @[:@144373.4]
  output [2:0]   io_M_AXI_1_ARSIZE, // @[:@144373.4]
  output [1:0]   io_M_AXI_1_ARBURST, // @[:@144373.4]
  output         io_M_AXI_1_ARLOCK, // @[:@144373.4]
  output [3:0]   io_M_AXI_1_ARCACHE, // @[:@144373.4]
  output [2:0]   io_M_AXI_1_ARPROT, // @[:@144373.4]
  output [3:0]   io_M_AXI_1_ARQOS, // @[:@144373.4]
  output         io_M_AXI_1_ARVALID, // @[:@144373.4]
  input          io_M_AXI_1_ARREADY, // @[:@144373.4]
  output [511:0] io_M_AXI_1_WDATA, // @[:@144373.4]
  output [63:0]  io_M_AXI_1_WSTRB, // @[:@144373.4]
  output         io_M_AXI_1_WLAST, // @[:@144373.4]
  output         io_M_AXI_1_WVALID, // @[:@144373.4]
  input          io_M_AXI_1_WREADY, // @[:@144373.4]
  input  [31:0]  io_M_AXI_1_RID, // @[:@144373.4]
  input  [31:0]  io_M_AXI_1_RUSER, // @[:@144373.4]
  input  [511:0] io_M_AXI_1_RDATA, // @[:@144373.4]
  input  [1:0]   io_M_AXI_1_RRESP, // @[:@144373.4]
  input          io_M_AXI_1_RLAST, // @[:@144373.4]
  input          io_M_AXI_1_RVALID, // @[:@144373.4]
  output         io_M_AXI_1_RREADY, // @[:@144373.4]
  input  [31:0]  io_M_AXI_1_BID, // @[:@144373.4]
  input  [31:0]  io_M_AXI_1_BUSER, // @[:@144373.4]
  input  [1:0]   io_M_AXI_1_BRESP, // @[:@144373.4]
  input          io_M_AXI_1_BVALID, // @[:@144373.4]
  output         io_M_AXI_1_BREADY, // @[:@144373.4]
  output [31:0]  io_M_AXI_2_AWID, // @[:@144373.4]
  output [31:0]  io_M_AXI_2_AWUSER, // @[:@144373.4]
  output [31:0]  io_M_AXI_2_AWADDR, // @[:@144373.4]
  output [7:0]   io_M_AXI_2_AWLEN, // @[:@144373.4]
  output [2:0]   io_M_AXI_2_AWSIZE, // @[:@144373.4]
  output [1:0]   io_M_AXI_2_AWBURST, // @[:@144373.4]
  output         io_M_AXI_2_AWLOCK, // @[:@144373.4]
  output [3:0]   io_M_AXI_2_AWCACHE, // @[:@144373.4]
  output [2:0]   io_M_AXI_2_AWPROT, // @[:@144373.4]
  output [3:0]   io_M_AXI_2_AWQOS, // @[:@144373.4]
  output         io_M_AXI_2_AWVALID, // @[:@144373.4]
  input          io_M_AXI_2_AWREADY, // @[:@144373.4]
  output [31:0]  io_M_AXI_2_ARID, // @[:@144373.4]
  output [31:0]  io_M_AXI_2_ARUSER, // @[:@144373.4]
  output [31:0]  io_M_AXI_2_ARADDR, // @[:@144373.4]
  output [7:0]   io_M_AXI_2_ARLEN, // @[:@144373.4]
  output [2:0]   io_M_AXI_2_ARSIZE, // @[:@144373.4]
  output [1:0]   io_M_AXI_2_ARBURST, // @[:@144373.4]
  output         io_M_AXI_2_ARLOCK, // @[:@144373.4]
  output [3:0]   io_M_AXI_2_ARCACHE, // @[:@144373.4]
  output [2:0]   io_M_AXI_2_ARPROT, // @[:@144373.4]
  output [3:0]   io_M_AXI_2_ARQOS, // @[:@144373.4]
  output         io_M_AXI_2_ARVALID, // @[:@144373.4]
  input          io_M_AXI_2_ARREADY, // @[:@144373.4]
  output [511:0] io_M_AXI_2_WDATA, // @[:@144373.4]
  output [63:0]  io_M_AXI_2_WSTRB, // @[:@144373.4]
  output         io_M_AXI_2_WLAST, // @[:@144373.4]
  output         io_M_AXI_2_WVALID, // @[:@144373.4]
  input          io_M_AXI_2_WREADY, // @[:@144373.4]
  input  [31:0]  io_M_AXI_2_RID, // @[:@144373.4]
  input  [31:0]  io_M_AXI_2_RUSER, // @[:@144373.4]
  input  [511:0] io_M_AXI_2_RDATA, // @[:@144373.4]
  input  [1:0]   io_M_AXI_2_RRESP, // @[:@144373.4]
  input          io_M_AXI_2_RLAST, // @[:@144373.4]
  input          io_M_AXI_2_RVALID, // @[:@144373.4]
  output         io_M_AXI_2_RREADY, // @[:@144373.4]
  input  [31:0]  io_M_AXI_2_BID, // @[:@144373.4]
  input  [31:0]  io_M_AXI_2_BUSER, // @[:@144373.4]
  input  [1:0]   io_M_AXI_2_BRESP, // @[:@144373.4]
  input          io_M_AXI_2_BVALID, // @[:@144373.4]
  output         io_M_AXI_2_BREADY, // @[:@144373.4]
  output [31:0]  io_M_AXI_3_AWID, // @[:@144373.4]
  output [31:0]  io_M_AXI_3_AWUSER, // @[:@144373.4]
  output [31:0]  io_M_AXI_3_AWADDR, // @[:@144373.4]
  output [7:0]   io_M_AXI_3_AWLEN, // @[:@144373.4]
  output [2:0]   io_M_AXI_3_AWSIZE, // @[:@144373.4]
  output [1:0]   io_M_AXI_3_AWBURST, // @[:@144373.4]
  output         io_M_AXI_3_AWLOCK, // @[:@144373.4]
  output [3:0]   io_M_AXI_3_AWCACHE, // @[:@144373.4]
  output [2:0]   io_M_AXI_3_AWPROT, // @[:@144373.4]
  output [3:0]   io_M_AXI_3_AWQOS, // @[:@144373.4]
  output         io_M_AXI_3_AWVALID, // @[:@144373.4]
  input          io_M_AXI_3_AWREADY, // @[:@144373.4]
  output [31:0]  io_M_AXI_3_ARID, // @[:@144373.4]
  output [31:0]  io_M_AXI_3_ARUSER, // @[:@144373.4]
  output [31:0]  io_M_AXI_3_ARADDR, // @[:@144373.4]
  output [7:0]   io_M_AXI_3_ARLEN, // @[:@144373.4]
  output [2:0]   io_M_AXI_3_ARSIZE, // @[:@144373.4]
  output [1:0]   io_M_AXI_3_ARBURST, // @[:@144373.4]
  output         io_M_AXI_3_ARLOCK, // @[:@144373.4]
  output [3:0]   io_M_AXI_3_ARCACHE, // @[:@144373.4]
  output [2:0]   io_M_AXI_3_ARPROT, // @[:@144373.4]
  output [3:0]   io_M_AXI_3_ARQOS, // @[:@144373.4]
  output         io_M_AXI_3_ARVALID, // @[:@144373.4]
  input          io_M_AXI_3_ARREADY, // @[:@144373.4]
  output [511:0] io_M_AXI_3_WDATA, // @[:@144373.4]
  output [63:0]  io_M_AXI_3_WSTRB, // @[:@144373.4]
  output         io_M_AXI_3_WLAST, // @[:@144373.4]
  output         io_M_AXI_3_WVALID, // @[:@144373.4]
  input          io_M_AXI_3_WREADY, // @[:@144373.4]
  input  [31:0]  io_M_AXI_3_RID, // @[:@144373.4]
  input  [31:0]  io_M_AXI_3_RUSER, // @[:@144373.4]
  input  [511:0] io_M_AXI_3_RDATA, // @[:@144373.4]
  input  [1:0]   io_M_AXI_3_RRESP, // @[:@144373.4]
  input          io_M_AXI_3_RLAST, // @[:@144373.4]
  input          io_M_AXI_3_RVALID, // @[:@144373.4]
  output         io_M_AXI_3_RREADY, // @[:@144373.4]
  input  [31:0]  io_M_AXI_3_BID, // @[:@144373.4]
  input  [31:0]  io_M_AXI_3_BUSER, // @[:@144373.4]
  input  [1:0]   io_M_AXI_3_BRESP, // @[:@144373.4]
  input          io_M_AXI_3_BVALID, // @[:@144373.4]
  output         io_M_AXI_3_BREADY, // @[:@144373.4]
  input          io_TOP_AXI_AWID, // @[:@144373.4]
  input          io_TOP_AXI_AWUSER, // @[:@144373.4]
  input  [31:0]  io_TOP_AXI_AWADDR, // @[:@144373.4]
  input  [7:0]   io_TOP_AXI_AWLEN, // @[:@144373.4]
  input  [2:0]   io_TOP_AXI_AWSIZE, // @[:@144373.4]
  input  [1:0]   io_TOP_AXI_AWBURST, // @[:@144373.4]
  input          io_TOP_AXI_AWLOCK, // @[:@144373.4]
  input  [3:0]   io_TOP_AXI_AWCACHE, // @[:@144373.4]
  input  [2:0]   io_TOP_AXI_AWPROT, // @[:@144373.4]
  input  [3:0]   io_TOP_AXI_AWQOS, // @[:@144373.4]
  input          io_TOP_AXI_AWVALID, // @[:@144373.4]
  input          io_TOP_AXI_AWREADY, // @[:@144373.4]
  input          io_TOP_AXI_ARID, // @[:@144373.4]
  input          io_TOP_AXI_ARUSER, // @[:@144373.4]
  input  [31:0]  io_TOP_AXI_ARADDR, // @[:@144373.4]
  input  [7:0]   io_TOP_AXI_ARLEN, // @[:@144373.4]
  input  [2:0]   io_TOP_AXI_ARSIZE, // @[:@144373.4]
  input  [1:0]   io_TOP_AXI_ARBURST, // @[:@144373.4]
  input          io_TOP_AXI_ARLOCK, // @[:@144373.4]
  input  [3:0]   io_TOP_AXI_ARCACHE, // @[:@144373.4]
  input  [2:0]   io_TOP_AXI_ARPROT, // @[:@144373.4]
  input  [3:0]   io_TOP_AXI_ARQOS, // @[:@144373.4]
  input          io_TOP_AXI_ARVALID, // @[:@144373.4]
  input          io_TOP_AXI_ARREADY, // @[:@144373.4]
  input  [31:0]  io_TOP_AXI_WDATA, // @[:@144373.4]
  input  [63:0]  io_TOP_AXI_WSTRB, // @[:@144373.4]
  input          io_TOP_AXI_WLAST, // @[:@144373.4]
  input          io_TOP_AXI_WVALID, // @[:@144373.4]
  input          io_TOP_AXI_WREADY, // @[:@144373.4]
  input          io_TOP_AXI_RID, // @[:@144373.4]
  input          io_TOP_AXI_RUSER, // @[:@144373.4]
  input  [31:0]  io_TOP_AXI_RDATA, // @[:@144373.4]
  input  [1:0]   io_TOP_AXI_RRESP, // @[:@144373.4]
  input          io_TOP_AXI_RLAST, // @[:@144373.4]
  input          io_TOP_AXI_RVALID, // @[:@144373.4]
  input          io_TOP_AXI_RREADY, // @[:@144373.4]
  input          io_TOP_AXI_BID, // @[:@144373.4]
  input          io_TOP_AXI_BUSER, // @[:@144373.4]
  input  [1:0]   io_TOP_AXI_BRESP, // @[:@144373.4]
  input          io_TOP_AXI_BVALID, // @[:@144373.4]
  input          io_TOP_AXI_BREADY, // @[:@144373.4]
  input          io_DWIDTH_AXI_AWID, // @[:@144373.4]
  input          io_DWIDTH_AXI_AWUSER, // @[:@144373.4]
  input  [31:0]  io_DWIDTH_AXI_AWADDR, // @[:@144373.4]
  input  [7:0]   io_DWIDTH_AXI_AWLEN, // @[:@144373.4]
  input  [2:0]   io_DWIDTH_AXI_AWSIZE, // @[:@144373.4]
  input  [1:0]   io_DWIDTH_AXI_AWBURST, // @[:@144373.4]
  input          io_DWIDTH_AXI_AWLOCK, // @[:@144373.4]
  input  [3:0]   io_DWIDTH_AXI_AWCACHE, // @[:@144373.4]
  input  [2:0]   io_DWIDTH_AXI_AWPROT, // @[:@144373.4]
  input  [3:0]   io_DWIDTH_AXI_AWQOS, // @[:@144373.4]
  input          io_DWIDTH_AXI_AWVALID, // @[:@144373.4]
  input          io_DWIDTH_AXI_AWREADY, // @[:@144373.4]
  input          io_DWIDTH_AXI_ARID, // @[:@144373.4]
  input          io_DWIDTH_AXI_ARUSER, // @[:@144373.4]
  input  [31:0]  io_DWIDTH_AXI_ARADDR, // @[:@144373.4]
  input  [7:0]   io_DWIDTH_AXI_ARLEN, // @[:@144373.4]
  input  [2:0]   io_DWIDTH_AXI_ARSIZE, // @[:@144373.4]
  input  [1:0]   io_DWIDTH_AXI_ARBURST, // @[:@144373.4]
  input          io_DWIDTH_AXI_ARLOCK, // @[:@144373.4]
  input  [3:0]   io_DWIDTH_AXI_ARCACHE, // @[:@144373.4]
  input  [2:0]   io_DWIDTH_AXI_ARPROT, // @[:@144373.4]
  input  [3:0]   io_DWIDTH_AXI_ARQOS, // @[:@144373.4]
  input          io_DWIDTH_AXI_ARVALID, // @[:@144373.4]
  input          io_DWIDTH_AXI_ARREADY, // @[:@144373.4]
  input  [31:0]  io_DWIDTH_AXI_WDATA, // @[:@144373.4]
  input  [63:0]  io_DWIDTH_AXI_WSTRB, // @[:@144373.4]
  input          io_DWIDTH_AXI_WLAST, // @[:@144373.4]
  input          io_DWIDTH_AXI_WVALID, // @[:@144373.4]
  input          io_DWIDTH_AXI_WREADY, // @[:@144373.4]
  input          io_DWIDTH_AXI_RID, // @[:@144373.4]
  input          io_DWIDTH_AXI_RUSER, // @[:@144373.4]
  input  [31:0]  io_DWIDTH_AXI_RDATA, // @[:@144373.4]
  input  [1:0]   io_DWIDTH_AXI_RRESP, // @[:@144373.4]
  input          io_DWIDTH_AXI_RLAST, // @[:@144373.4]
  input          io_DWIDTH_AXI_RVALID, // @[:@144373.4]
  input          io_DWIDTH_AXI_RREADY, // @[:@144373.4]
  input          io_DWIDTH_AXI_BID, // @[:@144373.4]
  input          io_DWIDTH_AXI_BUSER, // @[:@144373.4]
  input  [1:0]   io_DWIDTH_AXI_BRESP, // @[:@144373.4]
  input          io_DWIDTH_AXI_BVALID, // @[:@144373.4]
  input          io_DWIDTH_AXI_BREADY, // @[:@144373.4]
  input          io_PROTOCOL_AXI_AWID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_AWUSER, // @[:@144373.4]
  input  [31:0]  io_PROTOCOL_AXI_AWADDR, // @[:@144373.4]
  input  [7:0]   io_PROTOCOL_AXI_AWLEN, // @[:@144373.4]
  input  [2:0]   io_PROTOCOL_AXI_AWSIZE, // @[:@144373.4]
  input  [1:0]   io_PROTOCOL_AXI_AWBURST, // @[:@144373.4]
  input          io_PROTOCOL_AXI_AWLOCK, // @[:@144373.4]
  input  [3:0]   io_PROTOCOL_AXI_AWCACHE, // @[:@144373.4]
  input  [2:0]   io_PROTOCOL_AXI_AWPROT, // @[:@144373.4]
  input  [3:0]   io_PROTOCOL_AXI_AWQOS, // @[:@144373.4]
  input          io_PROTOCOL_AXI_AWVALID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_AWREADY, // @[:@144373.4]
  input          io_PROTOCOL_AXI_ARID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_ARUSER, // @[:@144373.4]
  input  [31:0]  io_PROTOCOL_AXI_ARADDR, // @[:@144373.4]
  input  [7:0]   io_PROTOCOL_AXI_ARLEN, // @[:@144373.4]
  input  [2:0]   io_PROTOCOL_AXI_ARSIZE, // @[:@144373.4]
  input  [1:0]   io_PROTOCOL_AXI_ARBURST, // @[:@144373.4]
  input          io_PROTOCOL_AXI_ARLOCK, // @[:@144373.4]
  input  [3:0]   io_PROTOCOL_AXI_ARCACHE, // @[:@144373.4]
  input  [2:0]   io_PROTOCOL_AXI_ARPROT, // @[:@144373.4]
  input  [3:0]   io_PROTOCOL_AXI_ARQOS, // @[:@144373.4]
  input          io_PROTOCOL_AXI_ARVALID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_ARREADY, // @[:@144373.4]
  input  [31:0]  io_PROTOCOL_AXI_WDATA, // @[:@144373.4]
  input  [63:0]  io_PROTOCOL_AXI_WSTRB, // @[:@144373.4]
  input          io_PROTOCOL_AXI_WLAST, // @[:@144373.4]
  input          io_PROTOCOL_AXI_WVALID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_WREADY, // @[:@144373.4]
  input          io_PROTOCOL_AXI_RID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_RUSER, // @[:@144373.4]
  input  [31:0]  io_PROTOCOL_AXI_RDATA, // @[:@144373.4]
  input  [1:0]   io_PROTOCOL_AXI_RRESP, // @[:@144373.4]
  input          io_PROTOCOL_AXI_RLAST, // @[:@144373.4]
  input          io_PROTOCOL_AXI_RVALID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_RREADY, // @[:@144373.4]
  input          io_PROTOCOL_AXI_BID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_BUSER, // @[:@144373.4]
  input  [1:0]   io_PROTOCOL_AXI_BRESP, // @[:@144373.4]
  input          io_PROTOCOL_AXI_BVALID, // @[:@144373.4]
  input          io_PROTOCOL_AXI_BREADY, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_AWID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_AWUSER, // @[:@144373.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_AWADDR, // @[:@144373.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_AWLEN, // @[:@144373.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWSIZE, // @[:@144373.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_AWBURST, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_AWLOCK, // @[:@144373.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWCACHE, // @[:@144373.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_AWPROT, // @[:@144373.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_AWQOS, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_AWVALID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_AWREADY, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_ARID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_ARUSER, // @[:@144373.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_ARADDR, // @[:@144373.4]
  input  [7:0]   io_CLOCKCONVERT_AXI_ARLEN, // @[:@144373.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARSIZE, // @[:@144373.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_ARBURST, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_ARLOCK, // @[:@144373.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARCACHE, // @[:@144373.4]
  input  [2:0]   io_CLOCKCONVERT_AXI_ARPROT, // @[:@144373.4]
  input  [3:0]   io_CLOCKCONVERT_AXI_ARQOS, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_ARVALID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_ARREADY, // @[:@144373.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_WDATA, // @[:@144373.4]
  input  [63:0]  io_CLOCKCONVERT_AXI_WSTRB, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_WLAST, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_WVALID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_WREADY, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_RID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_RUSER, // @[:@144373.4]
  input  [31:0]  io_CLOCKCONVERT_AXI_RDATA, // @[:@144373.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_RRESP, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_RLAST, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_RVALID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_RREADY, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_BID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_BUSER, // @[:@144373.4]
  input  [1:0]   io_CLOCKCONVERT_AXI_BRESP, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_BVALID, // @[:@144373.4]
  input          io_CLOCKCONVERT_AXI_BREADY // @[:@144373.4]
);
  wire  accel_clock; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_reset; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_enable; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_done; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_reset; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_loads_0_cmd_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_loads_0_cmd_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_loads_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_cmd_bits_size; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_loads_0_data_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_loads_0_data_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_0; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_1; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_2; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_3; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_4; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_5; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_6; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_7; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_8; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_9; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_10; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_11; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_12; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_13; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_14; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_loads_0_data_bits_rdata_15; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_stores_0_cmd_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_stores_0_cmd_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_stores_0_cmd_bits_addr; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_stores_0_cmd_bits_size; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_stores_0_data_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_stores_0_data_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_stores_0_data_bits_wstrb; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_stores_0_wresp_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_stores_0_wresp_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_stores_0_wresp_bits; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_gathers_0_cmd_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_gathers_0_cmd_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_0; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_1; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_2; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_3; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_4; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_5; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_6; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_7; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_8; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_9; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_10; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_11; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_12; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_13; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_14; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_gathers_0_cmd_bits_addr_15; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_gathers_0_data_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_gathers_0_data_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_0; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_1; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_2; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_3; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_4; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_5; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_6; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_7; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_8; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_9; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_10; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_11; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_12; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_13; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_14; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_gathers_0_data_bits_15; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_scatters_0_cmd_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_scatters_0_cmd_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_0; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_1; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_2; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_3; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_4; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_5; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_6; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_7; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_8; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_9; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_10; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_11; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_12; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_13; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_14; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_memStreams_scatters_0_cmd_bits_wdata_15; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_scatters_0_wresp_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_scatters_0_wresp_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_memStreams_scatters_0_wresp_bits; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_axiStreamsIn_0_TVALID; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_axiStreamsIn_0_TREADY; // @[Instantiator.scala 53:44:@144375.4]
  wire [255:0] accel_io_axiStreamsIn_0_TDATA; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_axiStreamsIn_0_TSTRB; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_axiStreamsIn_0_TKEEP; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_axiStreamsIn_0_TLAST; // @[Instantiator.scala 53:44:@144375.4]
  wire [7:0] accel_io_axiStreamsIn_0_TID; // @[Instantiator.scala 53:44:@144375.4]
  wire [7:0] accel_io_axiStreamsIn_0_TDEST; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_axiStreamsIn_0_TUSER; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_axiStreamsOut_0_TVALID; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_axiStreamsOut_0_TREADY; // @[Instantiator.scala 53:44:@144375.4]
  wire [255:0] accel_io_axiStreamsOut_0_TDATA; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_axiStreamsOut_0_TSTRB; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_axiStreamsOut_0_TKEEP; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_axiStreamsOut_0_TLAST; // @[Instantiator.scala 53:44:@144375.4]
  wire [7:0] accel_io_axiStreamsOut_0_TID; // @[Instantiator.scala 53:44:@144375.4]
  wire [7:0] accel_io_axiStreamsOut_0_TDEST; // @[Instantiator.scala 53:44:@144375.4]
  wire [31:0] accel_io_axiStreamsOut_0_TUSER; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_heap_0_req_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_heap_0_req_bits_allocDealloc; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_heap_0_req_bits_sizeAddr; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_heap_0_resp_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_heap_0_resp_bits_allocDealloc; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_heap_0_resp_bits_sizeAddr; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_argIns_0; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_argIns_1; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_argOuts_0_port_ready; // @[Instantiator.scala 53:44:@144375.4]
  wire  accel_io_argOuts_0_port_valid; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_argOuts_0_port_bits; // @[Instantiator.scala 53:44:@144375.4]
  wire [63:0] accel_io_argOuts_0_echo; // @[Instantiator.scala 53:44:@144375.4]
  wire  FringeZynq_clock; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_reset; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_S_AXI_AWADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [2:0] FringeZynq_io_S_AXI_AWPROT; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_AWVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_S_AXI_ARADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [2:0] FringeZynq_io_S_AXI_ARPROT; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_ARVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_S_AXI_WDATA; // @[Zynq.scala 18:24:@144517.4]
  wire [3:0] FringeZynq_io_S_AXI_WSTRB; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_WVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 18:24:@144517.4]
  wire [1:0] FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_RREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [1:0] FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_S_AXI_BREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [7:0] FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_AWREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [7:0] FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_ARREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [511:0] FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_WREADY; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_0_BID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_BVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [7:0] FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_AWREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [7:0] FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_ARREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [511:0] FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_WREADY; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_1_BID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_BVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [7:0] FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_AWREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [7:0] FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_ARREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [511:0] FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_WREADY; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_2_BID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_BVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [7:0] FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_AWREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 18:24:@144517.4]
  wire [7:0] FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_ARREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [511:0] FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_WREADY; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_M_AXI_3_BID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_BVALID; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_enable; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_done; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_reset; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_argIns_0; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_argIns_1; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_argOuts_0_valid; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_argOuts_0_bits; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_memStreams_stores_0_data_valid; // @[Zynq.scala 18:24:@144517.4]
  wire [31:0] FringeZynq_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_heap_0_req_valid; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 18:24:@144517.4]
  wire  FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 18:24:@144517.4]
  wire [63:0] FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 18:24:@144517.4]
  AccelUnit accel ( // @[Instantiator.scala 53:44:@144375.4]
    .clock(accel_clock),
    .reset(accel_reset),
    .io_enable(accel_io_enable),
    .io_done(accel_io_done),
    .io_reset(accel_io_reset),
    .io_memStreams_loads_0_cmd_ready(accel_io_memStreams_loads_0_cmd_ready),
    .io_memStreams_loads_0_cmd_valid(accel_io_memStreams_loads_0_cmd_valid),
    .io_memStreams_loads_0_cmd_bits_addr(accel_io_memStreams_loads_0_cmd_bits_addr),
    .io_memStreams_loads_0_cmd_bits_size(accel_io_memStreams_loads_0_cmd_bits_size),
    .io_memStreams_loads_0_data_ready(accel_io_memStreams_loads_0_data_ready),
    .io_memStreams_loads_0_data_valid(accel_io_memStreams_loads_0_data_valid),
    .io_memStreams_loads_0_data_bits_rdata_0(accel_io_memStreams_loads_0_data_bits_rdata_0),
    .io_memStreams_loads_0_data_bits_rdata_1(accel_io_memStreams_loads_0_data_bits_rdata_1),
    .io_memStreams_loads_0_data_bits_rdata_2(accel_io_memStreams_loads_0_data_bits_rdata_2),
    .io_memStreams_loads_0_data_bits_rdata_3(accel_io_memStreams_loads_0_data_bits_rdata_3),
    .io_memStreams_loads_0_data_bits_rdata_4(accel_io_memStreams_loads_0_data_bits_rdata_4),
    .io_memStreams_loads_0_data_bits_rdata_5(accel_io_memStreams_loads_0_data_bits_rdata_5),
    .io_memStreams_loads_0_data_bits_rdata_6(accel_io_memStreams_loads_0_data_bits_rdata_6),
    .io_memStreams_loads_0_data_bits_rdata_7(accel_io_memStreams_loads_0_data_bits_rdata_7),
    .io_memStreams_loads_0_data_bits_rdata_8(accel_io_memStreams_loads_0_data_bits_rdata_8),
    .io_memStreams_loads_0_data_bits_rdata_9(accel_io_memStreams_loads_0_data_bits_rdata_9),
    .io_memStreams_loads_0_data_bits_rdata_10(accel_io_memStreams_loads_0_data_bits_rdata_10),
    .io_memStreams_loads_0_data_bits_rdata_11(accel_io_memStreams_loads_0_data_bits_rdata_11),
    .io_memStreams_loads_0_data_bits_rdata_12(accel_io_memStreams_loads_0_data_bits_rdata_12),
    .io_memStreams_loads_0_data_bits_rdata_13(accel_io_memStreams_loads_0_data_bits_rdata_13),
    .io_memStreams_loads_0_data_bits_rdata_14(accel_io_memStreams_loads_0_data_bits_rdata_14),
    .io_memStreams_loads_0_data_bits_rdata_15(accel_io_memStreams_loads_0_data_bits_rdata_15),
    .io_memStreams_stores_0_cmd_ready(accel_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(accel_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(accel_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(accel_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(accel_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(accel_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(accel_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(accel_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(accel_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(accel_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(accel_io_memStreams_stores_0_wresp_bits),
    .io_memStreams_gathers_0_cmd_ready(accel_io_memStreams_gathers_0_cmd_ready),
    .io_memStreams_gathers_0_cmd_valid(accel_io_memStreams_gathers_0_cmd_valid),
    .io_memStreams_gathers_0_cmd_bits_addr_0(accel_io_memStreams_gathers_0_cmd_bits_addr_0),
    .io_memStreams_gathers_0_cmd_bits_addr_1(accel_io_memStreams_gathers_0_cmd_bits_addr_1),
    .io_memStreams_gathers_0_cmd_bits_addr_2(accel_io_memStreams_gathers_0_cmd_bits_addr_2),
    .io_memStreams_gathers_0_cmd_bits_addr_3(accel_io_memStreams_gathers_0_cmd_bits_addr_3),
    .io_memStreams_gathers_0_cmd_bits_addr_4(accel_io_memStreams_gathers_0_cmd_bits_addr_4),
    .io_memStreams_gathers_0_cmd_bits_addr_5(accel_io_memStreams_gathers_0_cmd_bits_addr_5),
    .io_memStreams_gathers_0_cmd_bits_addr_6(accel_io_memStreams_gathers_0_cmd_bits_addr_6),
    .io_memStreams_gathers_0_cmd_bits_addr_7(accel_io_memStreams_gathers_0_cmd_bits_addr_7),
    .io_memStreams_gathers_0_cmd_bits_addr_8(accel_io_memStreams_gathers_0_cmd_bits_addr_8),
    .io_memStreams_gathers_0_cmd_bits_addr_9(accel_io_memStreams_gathers_0_cmd_bits_addr_9),
    .io_memStreams_gathers_0_cmd_bits_addr_10(accel_io_memStreams_gathers_0_cmd_bits_addr_10),
    .io_memStreams_gathers_0_cmd_bits_addr_11(accel_io_memStreams_gathers_0_cmd_bits_addr_11),
    .io_memStreams_gathers_0_cmd_bits_addr_12(accel_io_memStreams_gathers_0_cmd_bits_addr_12),
    .io_memStreams_gathers_0_cmd_bits_addr_13(accel_io_memStreams_gathers_0_cmd_bits_addr_13),
    .io_memStreams_gathers_0_cmd_bits_addr_14(accel_io_memStreams_gathers_0_cmd_bits_addr_14),
    .io_memStreams_gathers_0_cmd_bits_addr_15(accel_io_memStreams_gathers_0_cmd_bits_addr_15),
    .io_memStreams_gathers_0_data_ready(accel_io_memStreams_gathers_0_data_ready),
    .io_memStreams_gathers_0_data_valid(accel_io_memStreams_gathers_0_data_valid),
    .io_memStreams_gathers_0_data_bits_0(accel_io_memStreams_gathers_0_data_bits_0),
    .io_memStreams_gathers_0_data_bits_1(accel_io_memStreams_gathers_0_data_bits_1),
    .io_memStreams_gathers_0_data_bits_2(accel_io_memStreams_gathers_0_data_bits_2),
    .io_memStreams_gathers_0_data_bits_3(accel_io_memStreams_gathers_0_data_bits_3),
    .io_memStreams_gathers_0_data_bits_4(accel_io_memStreams_gathers_0_data_bits_4),
    .io_memStreams_gathers_0_data_bits_5(accel_io_memStreams_gathers_0_data_bits_5),
    .io_memStreams_gathers_0_data_bits_6(accel_io_memStreams_gathers_0_data_bits_6),
    .io_memStreams_gathers_0_data_bits_7(accel_io_memStreams_gathers_0_data_bits_7),
    .io_memStreams_gathers_0_data_bits_8(accel_io_memStreams_gathers_0_data_bits_8),
    .io_memStreams_gathers_0_data_bits_9(accel_io_memStreams_gathers_0_data_bits_9),
    .io_memStreams_gathers_0_data_bits_10(accel_io_memStreams_gathers_0_data_bits_10),
    .io_memStreams_gathers_0_data_bits_11(accel_io_memStreams_gathers_0_data_bits_11),
    .io_memStreams_gathers_0_data_bits_12(accel_io_memStreams_gathers_0_data_bits_12),
    .io_memStreams_gathers_0_data_bits_13(accel_io_memStreams_gathers_0_data_bits_13),
    .io_memStreams_gathers_0_data_bits_14(accel_io_memStreams_gathers_0_data_bits_14),
    .io_memStreams_gathers_0_data_bits_15(accel_io_memStreams_gathers_0_data_bits_15),
    .io_memStreams_scatters_0_cmd_ready(accel_io_memStreams_scatters_0_cmd_ready),
    .io_memStreams_scatters_0_cmd_valid(accel_io_memStreams_scatters_0_cmd_valid),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_0(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_0),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_1(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_1),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_2(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_2),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_3(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_3),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_4(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_4),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_5(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_5),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_6(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_6),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_7(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_7),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_8(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_8),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_9(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_9),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_10(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_10),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_11(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_11),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_12(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_12),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_13(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_13),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_14(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_14),
    .io_memStreams_scatters_0_cmd_bits_addr_addr_15(accel_io_memStreams_scatters_0_cmd_bits_addr_addr_15),
    .io_memStreams_scatters_0_cmd_bits_wdata_0(accel_io_memStreams_scatters_0_cmd_bits_wdata_0),
    .io_memStreams_scatters_0_cmd_bits_wdata_1(accel_io_memStreams_scatters_0_cmd_bits_wdata_1),
    .io_memStreams_scatters_0_cmd_bits_wdata_2(accel_io_memStreams_scatters_0_cmd_bits_wdata_2),
    .io_memStreams_scatters_0_cmd_bits_wdata_3(accel_io_memStreams_scatters_0_cmd_bits_wdata_3),
    .io_memStreams_scatters_0_cmd_bits_wdata_4(accel_io_memStreams_scatters_0_cmd_bits_wdata_4),
    .io_memStreams_scatters_0_cmd_bits_wdata_5(accel_io_memStreams_scatters_0_cmd_bits_wdata_5),
    .io_memStreams_scatters_0_cmd_bits_wdata_6(accel_io_memStreams_scatters_0_cmd_bits_wdata_6),
    .io_memStreams_scatters_0_cmd_bits_wdata_7(accel_io_memStreams_scatters_0_cmd_bits_wdata_7),
    .io_memStreams_scatters_0_cmd_bits_wdata_8(accel_io_memStreams_scatters_0_cmd_bits_wdata_8),
    .io_memStreams_scatters_0_cmd_bits_wdata_9(accel_io_memStreams_scatters_0_cmd_bits_wdata_9),
    .io_memStreams_scatters_0_cmd_bits_wdata_10(accel_io_memStreams_scatters_0_cmd_bits_wdata_10),
    .io_memStreams_scatters_0_cmd_bits_wdata_11(accel_io_memStreams_scatters_0_cmd_bits_wdata_11),
    .io_memStreams_scatters_0_cmd_bits_wdata_12(accel_io_memStreams_scatters_0_cmd_bits_wdata_12),
    .io_memStreams_scatters_0_cmd_bits_wdata_13(accel_io_memStreams_scatters_0_cmd_bits_wdata_13),
    .io_memStreams_scatters_0_cmd_bits_wdata_14(accel_io_memStreams_scatters_0_cmd_bits_wdata_14),
    .io_memStreams_scatters_0_cmd_bits_wdata_15(accel_io_memStreams_scatters_0_cmd_bits_wdata_15),
    .io_memStreams_scatters_0_wresp_ready(accel_io_memStreams_scatters_0_wresp_ready),
    .io_memStreams_scatters_0_wresp_valid(accel_io_memStreams_scatters_0_wresp_valid),
    .io_memStreams_scatters_0_wresp_bits(accel_io_memStreams_scatters_0_wresp_bits),
    .io_axiStreamsIn_0_TVALID(accel_io_axiStreamsIn_0_TVALID),
    .io_axiStreamsIn_0_TREADY(accel_io_axiStreamsIn_0_TREADY),
    .io_axiStreamsIn_0_TDATA(accel_io_axiStreamsIn_0_TDATA),
    .io_axiStreamsIn_0_TSTRB(accel_io_axiStreamsIn_0_TSTRB),
    .io_axiStreamsIn_0_TKEEP(accel_io_axiStreamsIn_0_TKEEP),
    .io_axiStreamsIn_0_TLAST(accel_io_axiStreamsIn_0_TLAST),
    .io_axiStreamsIn_0_TID(accel_io_axiStreamsIn_0_TID),
    .io_axiStreamsIn_0_TDEST(accel_io_axiStreamsIn_0_TDEST),
    .io_axiStreamsIn_0_TUSER(accel_io_axiStreamsIn_0_TUSER),
    .io_axiStreamsOut_0_TVALID(accel_io_axiStreamsOut_0_TVALID),
    .io_axiStreamsOut_0_TREADY(accel_io_axiStreamsOut_0_TREADY),
    .io_axiStreamsOut_0_TDATA(accel_io_axiStreamsOut_0_TDATA),
    .io_axiStreamsOut_0_TSTRB(accel_io_axiStreamsOut_0_TSTRB),
    .io_axiStreamsOut_0_TKEEP(accel_io_axiStreamsOut_0_TKEEP),
    .io_axiStreamsOut_0_TLAST(accel_io_axiStreamsOut_0_TLAST),
    .io_axiStreamsOut_0_TID(accel_io_axiStreamsOut_0_TID),
    .io_axiStreamsOut_0_TDEST(accel_io_axiStreamsOut_0_TDEST),
    .io_axiStreamsOut_0_TUSER(accel_io_axiStreamsOut_0_TUSER),
    .io_heap_0_req_valid(accel_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(accel_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(accel_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(accel_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(accel_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(accel_io_heap_0_resp_bits_sizeAddr),
    .io_argIns_0(accel_io_argIns_0),
    .io_argIns_1(accel_io_argIns_1),
    .io_argOuts_0_port_ready(accel_io_argOuts_0_port_ready),
    .io_argOuts_0_port_valid(accel_io_argOuts_0_port_valid),
    .io_argOuts_0_port_bits(accel_io_argOuts_0_port_bits),
    .io_argOuts_0_echo(accel_io_argOuts_0_echo)
  );
  FringeZynq FringeZynq ( // @[Zynq.scala 18:24:@144517.4]
    .clock(FringeZynq_clock),
    .reset(FringeZynq_reset),
    .io_S_AXI_AWADDR(FringeZynq_io_S_AXI_AWADDR),
    .io_S_AXI_AWPROT(FringeZynq_io_S_AXI_AWPROT),
    .io_S_AXI_AWVALID(FringeZynq_io_S_AXI_AWVALID),
    .io_S_AXI_AWREADY(FringeZynq_io_S_AXI_AWREADY),
    .io_S_AXI_ARADDR(FringeZynq_io_S_AXI_ARADDR),
    .io_S_AXI_ARPROT(FringeZynq_io_S_AXI_ARPROT),
    .io_S_AXI_ARVALID(FringeZynq_io_S_AXI_ARVALID),
    .io_S_AXI_ARREADY(FringeZynq_io_S_AXI_ARREADY),
    .io_S_AXI_WDATA(FringeZynq_io_S_AXI_WDATA),
    .io_S_AXI_WSTRB(FringeZynq_io_S_AXI_WSTRB),
    .io_S_AXI_WVALID(FringeZynq_io_S_AXI_WVALID),
    .io_S_AXI_WREADY(FringeZynq_io_S_AXI_WREADY),
    .io_S_AXI_RDATA(FringeZynq_io_S_AXI_RDATA),
    .io_S_AXI_RRESP(FringeZynq_io_S_AXI_RRESP),
    .io_S_AXI_RVALID(FringeZynq_io_S_AXI_RVALID),
    .io_S_AXI_RREADY(FringeZynq_io_S_AXI_RREADY),
    .io_S_AXI_BRESP(FringeZynq_io_S_AXI_BRESP),
    .io_S_AXI_BVALID(FringeZynq_io_S_AXI_BVALID),
    .io_S_AXI_BREADY(FringeZynq_io_S_AXI_BREADY),
    .io_M_AXI_0_AWID(FringeZynq_io_M_AXI_0_AWID),
    .io_M_AXI_0_AWADDR(FringeZynq_io_M_AXI_0_AWADDR),
    .io_M_AXI_0_AWLEN(FringeZynq_io_M_AXI_0_AWLEN),
    .io_M_AXI_0_AWVALID(FringeZynq_io_M_AXI_0_AWVALID),
    .io_M_AXI_0_AWREADY(FringeZynq_io_M_AXI_0_AWREADY),
    .io_M_AXI_0_ARID(FringeZynq_io_M_AXI_0_ARID),
    .io_M_AXI_0_ARADDR(FringeZynq_io_M_AXI_0_ARADDR),
    .io_M_AXI_0_ARLEN(FringeZynq_io_M_AXI_0_ARLEN),
    .io_M_AXI_0_ARVALID(FringeZynq_io_M_AXI_0_ARVALID),
    .io_M_AXI_0_ARREADY(FringeZynq_io_M_AXI_0_ARREADY),
    .io_M_AXI_0_WDATA(FringeZynq_io_M_AXI_0_WDATA),
    .io_M_AXI_0_WSTRB(FringeZynq_io_M_AXI_0_WSTRB),
    .io_M_AXI_0_WLAST(FringeZynq_io_M_AXI_0_WLAST),
    .io_M_AXI_0_WVALID(FringeZynq_io_M_AXI_0_WVALID),
    .io_M_AXI_0_WREADY(FringeZynq_io_M_AXI_0_WREADY),
    .io_M_AXI_0_RREADY(FringeZynq_io_M_AXI_0_RREADY),
    .io_M_AXI_0_BID(FringeZynq_io_M_AXI_0_BID),
    .io_M_AXI_0_BVALID(FringeZynq_io_M_AXI_0_BVALID),
    .io_M_AXI_0_BREADY(FringeZynq_io_M_AXI_0_BREADY),
    .io_M_AXI_1_AWID(FringeZynq_io_M_AXI_1_AWID),
    .io_M_AXI_1_AWADDR(FringeZynq_io_M_AXI_1_AWADDR),
    .io_M_AXI_1_AWLEN(FringeZynq_io_M_AXI_1_AWLEN),
    .io_M_AXI_1_AWVALID(FringeZynq_io_M_AXI_1_AWVALID),
    .io_M_AXI_1_AWREADY(FringeZynq_io_M_AXI_1_AWREADY),
    .io_M_AXI_1_ARID(FringeZynq_io_M_AXI_1_ARID),
    .io_M_AXI_1_ARADDR(FringeZynq_io_M_AXI_1_ARADDR),
    .io_M_AXI_1_ARLEN(FringeZynq_io_M_AXI_1_ARLEN),
    .io_M_AXI_1_ARVALID(FringeZynq_io_M_AXI_1_ARVALID),
    .io_M_AXI_1_ARREADY(FringeZynq_io_M_AXI_1_ARREADY),
    .io_M_AXI_1_WDATA(FringeZynq_io_M_AXI_1_WDATA),
    .io_M_AXI_1_WSTRB(FringeZynq_io_M_AXI_1_WSTRB),
    .io_M_AXI_1_WLAST(FringeZynq_io_M_AXI_1_WLAST),
    .io_M_AXI_1_WVALID(FringeZynq_io_M_AXI_1_WVALID),
    .io_M_AXI_1_WREADY(FringeZynq_io_M_AXI_1_WREADY),
    .io_M_AXI_1_RREADY(FringeZynq_io_M_AXI_1_RREADY),
    .io_M_AXI_1_BID(FringeZynq_io_M_AXI_1_BID),
    .io_M_AXI_1_BVALID(FringeZynq_io_M_AXI_1_BVALID),
    .io_M_AXI_1_BREADY(FringeZynq_io_M_AXI_1_BREADY),
    .io_M_AXI_2_AWID(FringeZynq_io_M_AXI_2_AWID),
    .io_M_AXI_2_AWADDR(FringeZynq_io_M_AXI_2_AWADDR),
    .io_M_AXI_2_AWLEN(FringeZynq_io_M_AXI_2_AWLEN),
    .io_M_AXI_2_AWVALID(FringeZynq_io_M_AXI_2_AWVALID),
    .io_M_AXI_2_AWREADY(FringeZynq_io_M_AXI_2_AWREADY),
    .io_M_AXI_2_ARID(FringeZynq_io_M_AXI_2_ARID),
    .io_M_AXI_2_ARADDR(FringeZynq_io_M_AXI_2_ARADDR),
    .io_M_AXI_2_ARLEN(FringeZynq_io_M_AXI_2_ARLEN),
    .io_M_AXI_2_ARVALID(FringeZynq_io_M_AXI_2_ARVALID),
    .io_M_AXI_2_ARREADY(FringeZynq_io_M_AXI_2_ARREADY),
    .io_M_AXI_2_WDATA(FringeZynq_io_M_AXI_2_WDATA),
    .io_M_AXI_2_WSTRB(FringeZynq_io_M_AXI_2_WSTRB),
    .io_M_AXI_2_WLAST(FringeZynq_io_M_AXI_2_WLAST),
    .io_M_AXI_2_WVALID(FringeZynq_io_M_AXI_2_WVALID),
    .io_M_AXI_2_WREADY(FringeZynq_io_M_AXI_2_WREADY),
    .io_M_AXI_2_RREADY(FringeZynq_io_M_AXI_2_RREADY),
    .io_M_AXI_2_BID(FringeZynq_io_M_AXI_2_BID),
    .io_M_AXI_2_BVALID(FringeZynq_io_M_AXI_2_BVALID),
    .io_M_AXI_2_BREADY(FringeZynq_io_M_AXI_2_BREADY),
    .io_M_AXI_3_AWID(FringeZynq_io_M_AXI_3_AWID),
    .io_M_AXI_3_AWADDR(FringeZynq_io_M_AXI_3_AWADDR),
    .io_M_AXI_3_AWLEN(FringeZynq_io_M_AXI_3_AWLEN),
    .io_M_AXI_3_AWVALID(FringeZynq_io_M_AXI_3_AWVALID),
    .io_M_AXI_3_AWREADY(FringeZynq_io_M_AXI_3_AWREADY),
    .io_M_AXI_3_ARID(FringeZynq_io_M_AXI_3_ARID),
    .io_M_AXI_3_ARADDR(FringeZynq_io_M_AXI_3_ARADDR),
    .io_M_AXI_3_ARLEN(FringeZynq_io_M_AXI_3_ARLEN),
    .io_M_AXI_3_ARVALID(FringeZynq_io_M_AXI_3_ARVALID),
    .io_M_AXI_3_ARREADY(FringeZynq_io_M_AXI_3_ARREADY),
    .io_M_AXI_3_WDATA(FringeZynq_io_M_AXI_3_WDATA),
    .io_M_AXI_3_WSTRB(FringeZynq_io_M_AXI_3_WSTRB),
    .io_M_AXI_3_WLAST(FringeZynq_io_M_AXI_3_WLAST),
    .io_M_AXI_3_WVALID(FringeZynq_io_M_AXI_3_WVALID),
    .io_M_AXI_3_WREADY(FringeZynq_io_M_AXI_3_WREADY),
    .io_M_AXI_3_RREADY(FringeZynq_io_M_AXI_3_RREADY),
    .io_M_AXI_3_BID(FringeZynq_io_M_AXI_3_BID),
    .io_M_AXI_3_BVALID(FringeZynq_io_M_AXI_3_BVALID),
    .io_M_AXI_3_BREADY(FringeZynq_io_M_AXI_3_BREADY),
    .io_enable(FringeZynq_io_enable),
    .io_done(FringeZynq_io_done),
    .io_reset(FringeZynq_io_reset),
    .io_argIns_0(FringeZynq_io_argIns_0),
    .io_argIns_1(FringeZynq_io_argIns_1),
    .io_argOuts_0_valid(FringeZynq_io_argOuts_0_valid),
    .io_argOuts_0_bits(FringeZynq_io_argOuts_0_bits),
    .io_memStreams_stores_0_cmd_ready(FringeZynq_io_memStreams_stores_0_cmd_ready),
    .io_memStreams_stores_0_cmd_valid(FringeZynq_io_memStreams_stores_0_cmd_valid),
    .io_memStreams_stores_0_cmd_bits_addr(FringeZynq_io_memStreams_stores_0_cmd_bits_addr),
    .io_memStreams_stores_0_cmd_bits_size(FringeZynq_io_memStreams_stores_0_cmd_bits_size),
    .io_memStreams_stores_0_data_ready(FringeZynq_io_memStreams_stores_0_data_ready),
    .io_memStreams_stores_0_data_valid(FringeZynq_io_memStreams_stores_0_data_valid),
    .io_memStreams_stores_0_data_bits_wdata_0(FringeZynq_io_memStreams_stores_0_data_bits_wdata_0),
    .io_memStreams_stores_0_data_bits_wstrb(FringeZynq_io_memStreams_stores_0_data_bits_wstrb),
    .io_memStreams_stores_0_wresp_ready(FringeZynq_io_memStreams_stores_0_wresp_ready),
    .io_memStreams_stores_0_wresp_valid(FringeZynq_io_memStreams_stores_0_wresp_valid),
    .io_memStreams_stores_0_wresp_bits(FringeZynq_io_memStreams_stores_0_wresp_bits),
    .io_heap_0_req_valid(FringeZynq_io_heap_0_req_valid),
    .io_heap_0_req_bits_allocDealloc(FringeZynq_io_heap_0_req_bits_allocDealloc),
    .io_heap_0_req_bits_sizeAddr(FringeZynq_io_heap_0_req_bits_sizeAddr),
    .io_heap_0_resp_valid(FringeZynq_io_heap_0_resp_valid),
    .io_heap_0_resp_bits_allocDealloc(FringeZynq_io_heap_0_resp_bits_allocDealloc),
    .io_heap_0_resp_bits_sizeAddr(FringeZynq_io_heap_0_resp_bits_sizeAddr)
  );
  assign io_rdata = 1'h0;
  assign io_S_AXI_AWREADY = FringeZynq_io_S_AXI_AWREADY; // @[Zynq.scala 21:21:@144535.4]
  assign io_S_AXI_ARREADY = FringeZynq_io_S_AXI_ARREADY; // @[Zynq.scala 21:21:@144531.4]
  assign io_S_AXI_WREADY = FringeZynq_io_S_AXI_WREADY; // @[Zynq.scala 21:21:@144527.4]
  assign io_S_AXI_RDATA = FringeZynq_io_S_AXI_RDATA; // @[Zynq.scala 21:21:@144526.4]
  assign io_S_AXI_RRESP = FringeZynq_io_S_AXI_RRESP; // @[Zynq.scala 21:21:@144525.4]
  assign io_S_AXI_RVALID = FringeZynq_io_S_AXI_RVALID; // @[Zynq.scala 21:21:@144524.4]
  assign io_S_AXI_BRESP = FringeZynq_io_S_AXI_BRESP; // @[Zynq.scala 21:21:@144522.4]
  assign io_S_AXI_BVALID = FringeZynq_io_S_AXI_BVALID; // @[Zynq.scala 21:21:@144521.4]
  assign io_M_AXI_0_AWID = FringeZynq_io_M_AXI_0_AWID; // @[Zynq.scala 24:14:@144579.4]
  assign io_M_AXI_0_AWUSER = 32'h0; // @[Zynq.scala 24:14:@144578.4]
  assign io_M_AXI_0_AWADDR = FringeZynq_io_M_AXI_0_AWADDR; // @[Zynq.scala 24:14:@144577.4]
  assign io_M_AXI_0_AWLEN = FringeZynq_io_M_AXI_0_AWLEN; // @[Zynq.scala 24:14:@144576.4]
  assign io_M_AXI_0_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@144575.4]
  assign io_M_AXI_0_AWBURST = 2'h1; // @[Zynq.scala 24:14:@144574.4]
  assign io_M_AXI_0_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@144573.4]
  assign io_M_AXI_0_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@144572.4]
  assign io_M_AXI_0_AWPROT = 3'h0; // @[Zynq.scala 24:14:@144571.4]
  assign io_M_AXI_0_AWQOS = 4'h0; // @[Zynq.scala 24:14:@144570.4]
  assign io_M_AXI_0_AWVALID = FringeZynq_io_M_AXI_0_AWVALID; // @[Zynq.scala 24:14:@144569.4]
  assign io_M_AXI_0_ARID = FringeZynq_io_M_AXI_0_ARID; // @[Zynq.scala 24:14:@144567.4]
  assign io_M_AXI_0_ARUSER = 32'h0; // @[Zynq.scala 24:14:@144566.4]
  assign io_M_AXI_0_ARADDR = FringeZynq_io_M_AXI_0_ARADDR; // @[Zynq.scala 24:14:@144565.4]
  assign io_M_AXI_0_ARLEN = FringeZynq_io_M_AXI_0_ARLEN; // @[Zynq.scala 24:14:@144564.4]
  assign io_M_AXI_0_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@144563.4]
  assign io_M_AXI_0_ARBURST = 2'h1; // @[Zynq.scala 24:14:@144562.4]
  assign io_M_AXI_0_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@144561.4]
  assign io_M_AXI_0_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@144560.4]
  assign io_M_AXI_0_ARPROT = 3'h0; // @[Zynq.scala 24:14:@144559.4]
  assign io_M_AXI_0_ARQOS = 4'h0; // @[Zynq.scala 24:14:@144558.4]
  assign io_M_AXI_0_ARVALID = FringeZynq_io_M_AXI_0_ARVALID; // @[Zynq.scala 24:14:@144557.4]
  assign io_M_AXI_0_WDATA = FringeZynq_io_M_AXI_0_WDATA; // @[Zynq.scala 24:14:@144555.4]
  assign io_M_AXI_0_WSTRB = FringeZynq_io_M_AXI_0_WSTRB; // @[Zynq.scala 24:14:@144554.4]
  assign io_M_AXI_0_WLAST = FringeZynq_io_M_AXI_0_WLAST; // @[Zynq.scala 24:14:@144553.4]
  assign io_M_AXI_0_WVALID = FringeZynq_io_M_AXI_0_WVALID; // @[Zynq.scala 24:14:@144552.4]
  assign io_M_AXI_0_RREADY = FringeZynq_io_M_AXI_0_RREADY; // @[Zynq.scala 24:14:@144544.4]
  assign io_M_AXI_0_BREADY = FringeZynq_io_M_AXI_0_BREADY; // @[Zynq.scala 24:14:@144539.4]
  assign io_M_AXI_1_AWID = FringeZynq_io_M_AXI_1_AWID; // @[Zynq.scala 24:14:@144620.4]
  assign io_M_AXI_1_AWUSER = 32'h0; // @[Zynq.scala 24:14:@144619.4]
  assign io_M_AXI_1_AWADDR = FringeZynq_io_M_AXI_1_AWADDR; // @[Zynq.scala 24:14:@144618.4]
  assign io_M_AXI_1_AWLEN = FringeZynq_io_M_AXI_1_AWLEN; // @[Zynq.scala 24:14:@144617.4]
  assign io_M_AXI_1_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@144616.4]
  assign io_M_AXI_1_AWBURST = 2'h1; // @[Zynq.scala 24:14:@144615.4]
  assign io_M_AXI_1_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@144614.4]
  assign io_M_AXI_1_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@144613.4]
  assign io_M_AXI_1_AWPROT = 3'h0; // @[Zynq.scala 24:14:@144612.4]
  assign io_M_AXI_1_AWQOS = 4'h0; // @[Zynq.scala 24:14:@144611.4]
  assign io_M_AXI_1_AWVALID = FringeZynq_io_M_AXI_1_AWVALID; // @[Zynq.scala 24:14:@144610.4]
  assign io_M_AXI_1_ARID = FringeZynq_io_M_AXI_1_ARID; // @[Zynq.scala 24:14:@144608.4]
  assign io_M_AXI_1_ARUSER = 32'h0; // @[Zynq.scala 24:14:@144607.4]
  assign io_M_AXI_1_ARADDR = FringeZynq_io_M_AXI_1_ARADDR; // @[Zynq.scala 24:14:@144606.4]
  assign io_M_AXI_1_ARLEN = FringeZynq_io_M_AXI_1_ARLEN; // @[Zynq.scala 24:14:@144605.4]
  assign io_M_AXI_1_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@144604.4]
  assign io_M_AXI_1_ARBURST = 2'h1; // @[Zynq.scala 24:14:@144603.4]
  assign io_M_AXI_1_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@144602.4]
  assign io_M_AXI_1_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@144601.4]
  assign io_M_AXI_1_ARPROT = 3'h0; // @[Zynq.scala 24:14:@144600.4]
  assign io_M_AXI_1_ARQOS = 4'h0; // @[Zynq.scala 24:14:@144599.4]
  assign io_M_AXI_1_ARVALID = FringeZynq_io_M_AXI_1_ARVALID; // @[Zynq.scala 24:14:@144598.4]
  assign io_M_AXI_1_WDATA = FringeZynq_io_M_AXI_1_WDATA; // @[Zynq.scala 24:14:@144596.4]
  assign io_M_AXI_1_WSTRB = FringeZynq_io_M_AXI_1_WSTRB; // @[Zynq.scala 24:14:@144595.4]
  assign io_M_AXI_1_WLAST = FringeZynq_io_M_AXI_1_WLAST; // @[Zynq.scala 24:14:@144594.4]
  assign io_M_AXI_1_WVALID = FringeZynq_io_M_AXI_1_WVALID; // @[Zynq.scala 24:14:@144593.4]
  assign io_M_AXI_1_RREADY = FringeZynq_io_M_AXI_1_RREADY; // @[Zynq.scala 24:14:@144585.4]
  assign io_M_AXI_1_BREADY = FringeZynq_io_M_AXI_1_BREADY; // @[Zynq.scala 24:14:@144580.4]
  assign io_M_AXI_2_AWID = FringeZynq_io_M_AXI_2_AWID; // @[Zynq.scala 24:14:@144661.4]
  assign io_M_AXI_2_AWUSER = 32'h0; // @[Zynq.scala 24:14:@144660.4]
  assign io_M_AXI_2_AWADDR = FringeZynq_io_M_AXI_2_AWADDR; // @[Zynq.scala 24:14:@144659.4]
  assign io_M_AXI_2_AWLEN = FringeZynq_io_M_AXI_2_AWLEN; // @[Zynq.scala 24:14:@144658.4]
  assign io_M_AXI_2_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@144657.4]
  assign io_M_AXI_2_AWBURST = 2'h1; // @[Zynq.scala 24:14:@144656.4]
  assign io_M_AXI_2_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@144655.4]
  assign io_M_AXI_2_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@144654.4]
  assign io_M_AXI_2_AWPROT = 3'h0; // @[Zynq.scala 24:14:@144653.4]
  assign io_M_AXI_2_AWQOS = 4'h0; // @[Zynq.scala 24:14:@144652.4]
  assign io_M_AXI_2_AWVALID = FringeZynq_io_M_AXI_2_AWVALID; // @[Zynq.scala 24:14:@144651.4]
  assign io_M_AXI_2_ARID = FringeZynq_io_M_AXI_2_ARID; // @[Zynq.scala 24:14:@144649.4]
  assign io_M_AXI_2_ARUSER = 32'h0; // @[Zynq.scala 24:14:@144648.4]
  assign io_M_AXI_2_ARADDR = FringeZynq_io_M_AXI_2_ARADDR; // @[Zynq.scala 24:14:@144647.4]
  assign io_M_AXI_2_ARLEN = FringeZynq_io_M_AXI_2_ARLEN; // @[Zynq.scala 24:14:@144646.4]
  assign io_M_AXI_2_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@144645.4]
  assign io_M_AXI_2_ARBURST = 2'h1; // @[Zynq.scala 24:14:@144644.4]
  assign io_M_AXI_2_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@144643.4]
  assign io_M_AXI_2_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@144642.4]
  assign io_M_AXI_2_ARPROT = 3'h0; // @[Zynq.scala 24:14:@144641.4]
  assign io_M_AXI_2_ARQOS = 4'h0; // @[Zynq.scala 24:14:@144640.4]
  assign io_M_AXI_2_ARVALID = FringeZynq_io_M_AXI_2_ARVALID; // @[Zynq.scala 24:14:@144639.4]
  assign io_M_AXI_2_WDATA = FringeZynq_io_M_AXI_2_WDATA; // @[Zynq.scala 24:14:@144637.4]
  assign io_M_AXI_2_WSTRB = FringeZynq_io_M_AXI_2_WSTRB; // @[Zynq.scala 24:14:@144636.4]
  assign io_M_AXI_2_WLAST = FringeZynq_io_M_AXI_2_WLAST; // @[Zynq.scala 24:14:@144635.4]
  assign io_M_AXI_2_WVALID = FringeZynq_io_M_AXI_2_WVALID; // @[Zynq.scala 24:14:@144634.4]
  assign io_M_AXI_2_RREADY = FringeZynq_io_M_AXI_2_RREADY; // @[Zynq.scala 24:14:@144626.4]
  assign io_M_AXI_2_BREADY = FringeZynq_io_M_AXI_2_BREADY; // @[Zynq.scala 24:14:@144621.4]
  assign io_M_AXI_3_AWID = FringeZynq_io_M_AXI_3_AWID; // @[Zynq.scala 24:14:@144702.4]
  assign io_M_AXI_3_AWUSER = 32'h0; // @[Zynq.scala 24:14:@144701.4]
  assign io_M_AXI_3_AWADDR = FringeZynq_io_M_AXI_3_AWADDR; // @[Zynq.scala 24:14:@144700.4]
  assign io_M_AXI_3_AWLEN = FringeZynq_io_M_AXI_3_AWLEN; // @[Zynq.scala 24:14:@144699.4]
  assign io_M_AXI_3_AWSIZE = 3'h6; // @[Zynq.scala 24:14:@144698.4]
  assign io_M_AXI_3_AWBURST = 2'h1; // @[Zynq.scala 24:14:@144697.4]
  assign io_M_AXI_3_AWLOCK = 1'h0; // @[Zynq.scala 24:14:@144696.4]
  assign io_M_AXI_3_AWCACHE = 4'h3; // @[Zynq.scala 24:14:@144695.4]
  assign io_M_AXI_3_AWPROT = 3'h0; // @[Zynq.scala 24:14:@144694.4]
  assign io_M_AXI_3_AWQOS = 4'h0; // @[Zynq.scala 24:14:@144693.4]
  assign io_M_AXI_3_AWVALID = FringeZynq_io_M_AXI_3_AWVALID; // @[Zynq.scala 24:14:@144692.4]
  assign io_M_AXI_3_ARID = FringeZynq_io_M_AXI_3_ARID; // @[Zynq.scala 24:14:@144690.4]
  assign io_M_AXI_3_ARUSER = 32'h0; // @[Zynq.scala 24:14:@144689.4]
  assign io_M_AXI_3_ARADDR = FringeZynq_io_M_AXI_3_ARADDR; // @[Zynq.scala 24:14:@144688.4]
  assign io_M_AXI_3_ARLEN = FringeZynq_io_M_AXI_3_ARLEN; // @[Zynq.scala 24:14:@144687.4]
  assign io_M_AXI_3_ARSIZE = 3'h6; // @[Zynq.scala 24:14:@144686.4]
  assign io_M_AXI_3_ARBURST = 2'h1; // @[Zynq.scala 24:14:@144685.4]
  assign io_M_AXI_3_ARLOCK = 1'h0; // @[Zynq.scala 24:14:@144684.4]
  assign io_M_AXI_3_ARCACHE = 4'h3; // @[Zynq.scala 24:14:@144683.4]
  assign io_M_AXI_3_ARPROT = 3'h0; // @[Zynq.scala 24:14:@144682.4]
  assign io_M_AXI_3_ARQOS = 4'h0; // @[Zynq.scala 24:14:@144681.4]
  assign io_M_AXI_3_ARVALID = FringeZynq_io_M_AXI_3_ARVALID; // @[Zynq.scala 24:14:@144680.4]
  assign io_M_AXI_3_WDATA = FringeZynq_io_M_AXI_3_WDATA; // @[Zynq.scala 24:14:@144678.4]
  assign io_M_AXI_3_WSTRB = FringeZynq_io_M_AXI_3_WSTRB; // @[Zynq.scala 24:14:@144677.4]
  assign io_M_AXI_3_WLAST = FringeZynq_io_M_AXI_3_WLAST; // @[Zynq.scala 24:14:@144676.4]
  assign io_M_AXI_3_WVALID = FringeZynq_io_M_AXI_3_WVALID; // @[Zynq.scala 24:14:@144675.4]
  assign io_M_AXI_3_RREADY = FringeZynq_io_M_AXI_3_RREADY; // @[Zynq.scala 24:14:@144667.4]
  assign io_M_AXI_3_BREADY = FringeZynq_io_M_AXI_3_BREADY; // @[Zynq.scala 24:14:@144662.4]
  assign accel_clock = clock; // @[:@144376.4]
  assign accel_reset = FringeZynq_io_reset; // @[:@144377.4 Zynq.scala 54:17:@144991.4]
  assign accel_io_enable = FringeZynq_io_enable; // @[Zynq.scala 51:21:@144986.4]
  assign accel_io_reset = 1'h0;
  assign accel_io_memStreams_loads_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@144979.4]
  assign accel_io_memStreams_loads_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@144974.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_0 = 32'h0; // @[Zynq.scala 49:26:@144958.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_1 = 32'h0; // @[Zynq.scala 49:26:@144959.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_2 = 32'h0; // @[Zynq.scala 49:26:@144960.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_3 = 32'h0; // @[Zynq.scala 49:26:@144961.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_4 = 32'h0; // @[Zynq.scala 49:26:@144962.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_5 = 32'h0; // @[Zynq.scala 49:26:@144963.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_6 = 32'h0; // @[Zynq.scala 49:26:@144964.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_7 = 32'h0; // @[Zynq.scala 49:26:@144965.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_8 = 32'h0; // @[Zynq.scala 49:26:@144966.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_9 = 32'h0; // @[Zynq.scala 49:26:@144967.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_10 = 32'h0; // @[Zynq.scala 49:26:@144968.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_11 = 32'h0; // @[Zynq.scala 49:26:@144969.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_12 = 32'h0; // @[Zynq.scala 49:26:@144970.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_13 = 32'h0; // @[Zynq.scala 49:26:@144971.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_14 = 32'h0; // @[Zynq.scala 49:26:@144972.4]
  assign accel_io_memStreams_loads_0_data_bits_rdata_15 = 32'h0; // @[Zynq.scala 49:26:@144973.4]
  assign accel_io_memStreams_stores_0_cmd_ready = FringeZynq_io_memStreams_stores_0_cmd_ready; // @[Zynq.scala 49:26:@144957.4]
  assign accel_io_memStreams_stores_0_data_ready = FringeZynq_io_memStreams_stores_0_data_ready; // @[Zynq.scala 49:26:@144953.4]
  assign accel_io_memStreams_stores_0_wresp_valid = FringeZynq_io_memStreams_stores_0_wresp_valid; // @[Zynq.scala 49:26:@144948.4]
  assign accel_io_memStreams_stores_0_wresp_bits = FringeZynq_io_memStreams_stores_0_wresp_bits; // @[Zynq.scala 49:26:@144947.4]
  assign accel_io_memStreams_gathers_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@144946.4]
  assign accel_io_memStreams_gathers_0_data_valid = 1'h0; // @[Zynq.scala 49:26:@144927.4]
  assign accel_io_memStreams_gathers_0_data_bits_0 = 32'h0; // @[Zynq.scala 49:26:@144911.4]
  assign accel_io_memStreams_gathers_0_data_bits_1 = 32'h0; // @[Zynq.scala 49:26:@144912.4]
  assign accel_io_memStreams_gathers_0_data_bits_2 = 32'h0; // @[Zynq.scala 49:26:@144913.4]
  assign accel_io_memStreams_gathers_0_data_bits_3 = 32'h0; // @[Zynq.scala 49:26:@144914.4]
  assign accel_io_memStreams_gathers_0_data_bits_4 = 32'h0; // @[Zynq.scala 49:26:@144915.4]
  assign accel_io_memStreams_gathers_0_data_bits_5 = 32'h0; // @[Zynq.scala 49:26:@144916.4]
  assign accel_io_memStreams_gathers_0_data_bits_6 = 32'h0; // @[Zynq.scala 49:26:@144917.4]
  assign accel_io_memStreams_gathers_0_data_bits_7 = 32'h0; // @[Zynq.scala 49:26:@144918.4]
  assign accel_io_memStreams_gathers_0_data_bits_8 = 32'h0; // @[Zynq.scala 49:26:@144919.4]
  assign accel_io_memStreams_gathers_0_data_bits_9 = 32'h0; // @[Zynq.scala 49:26:@144920.4]
  assign accel_io_memStreams_gathers_0_data_bits_10 = 32'h0; // @[Zynq.scala 49:26:@144921.4]
  assign accel_io_memStreams_gathers_0_data_bits_11 = 32'h0; // @[Zynq.scala 49:26:@144922.4]
  assign accel_io_memStreams_gathers_0_data_bits_12 = 32'h0; // @[Zynq.scala 49:26:@144923.4]
  assign accel_io_memStreams_gathers_0_data_bits_13 = 32'h0; // @[Zynq.scala 49:26:@144924.4]
  assign accel_io_memStreams_gathers_0_data_bits_14 = 32'h0; // @[Zynq.scala 49:26:@144925.4]
  assign accel_io_memStreams_gathers_0_data_bits_15 = 32'h0; // @[Zynq.scala 49:26:@144926.4]
  assign accel_io_memStreams_scatters_0_cmd_ready = 1'h0; // @[Zynq.scala 49:26:@144910.4]
  assign accel_io_memStreams_scatters_0_wresp_valid = 1'h0; // @[Zynq.scala 49:26:@144875.4]
  assign accel_io_memStreams_scatters_0_wresp_bits = 1'h0; // @[Zynq.scala 49:26:@144874.4]
  assign accel_io_axiStreamsIn_0_TVALID = 1'h0;
  assign accel_io_axiStreamsIn_0_TDATA = 256'h0;
  assign accel_io_axiStreamsIn_0_TSTRB = 32'h0;
  assign accel_io_axiStreamsIn_0_TKEEP = 32'h0;
  assign accel_io_axiStreamsIn_0_TLAST = 1'h0;
  assign accel_io_axiStreamsIn_0_TID = 8'h0;
  assign accel_io_axiStreamsIn_0_TDEST = 8'h0;
  assign accel_io_axiStreamsIn_0_TUSER = 32'h0;
  assign accel_io_axiStreamsOut_0_TREADY = 1'h0;
  assign accel_io_heap_0_resp_valid = FringeZynq_io_heap_0_resp_valid; // @[Zynq.scala 50:20:@144982.4]
  assign accel_io_heap_0_resp_bits_allocDealloc = FringeZynq_io_heap_0_resp_bits_allocDealloc; // @[Zynq.scala 50:20:@144981.4]
  assign accel_io_heap_0_resp_bits_sizeAddr = FringeZynq_io_heap_0_resp_bits_sizeAddr; // @[Zynq.scala 50:20:@144980.4]
  assign accel_io_argIns_0 = FringeZynq_io_argIns_0; // @[Zynq.scala 34:21:@144868.4]
  assign accel_io_argIns_1 = FringeZynq_io_argIns_1; // @[Zynq.scala 34:21:@144869.4]
  assign accel_io_argOuts_0_port_ready = 1'h0;
  assign accel_io_argOuts_0_echo = 64'h0; // @[Zynq.scala 40:24:@144872.4]
  assign FringeZynq_clock = clock; // @[:@144518.4]
  assign FringeZynq_reset = reset == 1'h0; // @[:@144519.4 Zynq.scala 53:18:@144990.4]
  assign FringeZynq_io_S_AXI_AWADDR = io_S_AXI_AWADDR; // @[Zynq.scala 21:21:@144538.4]
  assign FringeZynq_io_S_AXI_AWPROT = io_S_AXI_AWPROT; // @[Zynq.scala 21:21:@144537.4]
  assign FringeZynq_io_S_AXI_AWVALID = io_S_AXI_AWVALID; // @[Zynq.scala 21:21:@144536.4]
  assign FringeZynq_io_S_AXI_ARADDR = io_S_AXI_ARADDR; // @[Zynq.scala 21:21:@144534.4]
  assign FringeZynq_io_S_AXI_ARPROT = io_S_AXI_ARPROT; // @[Zynq.scala 21:21:@144533.4]
  assign FringeZynq_io_S_AXI_ARVALID = io_S_AXI_ARVALID; // @[Zynq.scala 21:21:@144532.4]
  assign FringeZynq_io_S_AXI_WDATA = io_S_AXI_WDATA; // @[Zynq.scala 21:21:@144530.4]
  assign FringeZynq_io_S_AXI_WSTRB = io_S_AXI_WSTRB; // @[Zynq.scala 21:21:@144529.4]
  assign FringeZynq_io_S_AXI_WVALID = io_S_AXI_WVALID; // @[Zynq.scala 21:21:@144528.4]
  assign FringeZynq_io_S_AXI_RREADY = io_S_AXI_RREADY; // @[Zynq.scala 21:21:@144523.4]
  assign FringeZynq_io_S_AXI_BREADY = io_S_AXI_BREADY; // @[Zynq.scala 21:21:@144520.4]
  assign FringeZynq_io_M_AXI_0_AWREADY = io_M_AXI_0_AWREADY; // @[Zynq.scala 24:14:@144568.4]
  assign FringeZynq_io_M_AXI_0_ARREADY = io_M_AXI_0_ARREADY; // @[Zynq.scala 24:14:@144556.4]
  assign FringeZynq_io_M_AXI_0_WREADY = io_M_AXI_0_WREADY; // @[Zynq.scala 24:14:@144551.4]
  assign FringeZynq_io_M_AXI_0_BID = io_M_AXI_0_BID; // @[Zynq.scala 24:14:@144543.4]
  assign FringeZynq_io_M_AXI_0_BVALID = io_M_AXI_0_BVALID; // @[Zynq.scala 24:14:@144540.4]
  assign FringeZynq_io_M_AXI_1_AWREADY = io_M_AXI_1_AWREADY; // @[Zynq.scala 24:14:@144609.4]
  assign FringeZynq_io_M_AXI_1_ARREADY = io_M_AXI_1_ARREADY; // @[Zynq.scala 24:14:@144597.4]
  assign FringeZynq_io_M_AXI_1_WREADY = io_M_AXI_1_WREADY; // @[Zynq.scala 24:14:@144592.4]
  assign FringeZynq_io_M_AXI_1_BID = io_M_AXI_1_BID; // @[Zynq.scala 24:14:@144584.4]
  assign FringeZynq_io_M_AXI_1_BVALID = io_M_AXI_1_BVALID; // @[Zynq.scala 24:14:@144581.4]
  assign FringeZynq_io_M_AXI_2_AWREADY = io_M_AXI_2_AWREADY; // @[Zynq.scala 24:14:@144650.4]
  assign FringeZynq_io_M_AXI_2_ARREADY = io_M_AXI_2_ARREADY; // @[Zynq.scala 24:14:@144638.4]
  assign FringeZynq_io_M_AXI_2_WREADY = io_M_AXI_2_WREADY; // @[Zynq.scala 24:14:@144633.4]
  assign FringeZynq_io_M_AXI_2_BID = io_M_AXI_2_BID; // @[Zynq.scala 24:14:@144625.4]
  assign FringeZynq_io_M_AXI_2_BVALID = io_M_AXI_2_BVALID; // @[Zynq.scala 24:14:@144622.4]
  assign FringeZynq_io_M_AXI_3_AWREADY = io_M_AXI_3_AWREADY; // @[Zynq.scala 24:14:@144691.4]
  assign FringeZynq_io_M_AXI_3_ARREADY = io_M_AXI_3_ARREADY; // @[Zynq.scala 24:14:@144679.4]
  assign FringeZynq_io_M_AXI_3_WREADY = io_M_AXI_3_WREADY; // @[Zynq.scala 24:14:@144674.4]
  assign FringeZynq_io_M_AXI_3_BID = io_M_AXI_3_BID; // @[Zynq.scala 24:14:@144666.4]
  assign FringeZynq_io_M_AXI_3_BVALID = io_M_AXI_3_BVALID; // @[Zynq.scala 24:14:@144663.4]
  assign FringeZynq_io_done = accel_io_done; // @[Zynq.scala 52:20:@144987.4]
  assign FringeZynq_io_argOuts_0_valid = accel_io_argOuts_0_port_valid; // @[Zynq.scala 37:26:@144871.4]
  assign FringeZynq_io_argOuts_0_bits = accel_io_argOuts_0_port_bits; // @[Zynq.scala 36:25:@144870.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_valid = accel_io_memStreams_stores_0_cmd_valid; // @[Zynq.scala 49:26:@144956.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_addr = accel_io_memStreams_stores_0_cmd_bits_addr; // @[Zynq.scala 49:26:@144955.4]
  assign FringeZynq_io_memStreams_stores_0_cmd_bits_size = accel_io_memStreams_stores_0_cmd_bits_size; // @[Zynq.scala 49:26:@144954.4]
  assign FringeZynq_io_memStreams_stores_0_data_valid = accel_io_memStreams_stores_0_data_valid; // @[Zynq.scala 49:26:@144952.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wdata_0 = accel_io_memStreams_stores_0_data_bits_wdata_0; // @[Zynq.scala 49:26:@144951.4]
  assign FringeZynq_io_memStreams_stores_0_data_bits_wstrb = accel_io_memStreams_stores_0_data_bits_wstrb; // @[Zynq.scala 49:26:@144950.4]
  assign FringeZynq_io_memStreams_stores_0_wresp_ready = accel_io_memStreams_stores_0_wresp_ready; // @[Zynq.scala 49:26:@144949.4]
  assign FringeZynq_io_heap_0_req_valid = accel_io_heap_0_req_valid; // @[Zynq.scala 50:20:@144985.4]
  assign FringeZynq_io_heap_0_req_bits_allocDealloc = accel_io_heap_0_req_bits_allocDealloc; // @[Zynq.scala 50:20:@144984.4]
  assign FringeZynq_io_heap_0_req_bits_sizeAddr = accel_io_heap_0_req_bits_sizeAddr; // @[Zynq.scala 50:20:@144983.4]
endmodule
module SRAMVerilogAWS
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr,
    input [AWIDTH-1:0] waddr,
    input raddrEn,
    input waddrEn,
    input wen,
    input [DWIDTH-1:0] wdata,
    input backpressure,
    output reg [DWIDTH-1:0] rdata
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk) begin
      if (wen) mem[waddr] <= wdata;
      if (backpressure) rdata <= mem[raddr];
    end

endmodule
module SRAMVerilogDualRead
#(
    parameter WORDS = 1024,
    parameter AWIDTH = 10,
    parameter DWIDTH = 32)
(
    input clk,
    input [AWIDTH-1:0] raddr0,
    input [AWIDTH-1:0] raddr1,
    input [AWIDTH-1:0] waddr,
    input raddrEn0,
    input raddrEn1,
    input waddrEn,
    input wen,
    input backpressure0,
    input backpressure1,
    input [DWIDTH-1:0] wdata,
    output reg [DWIDTH-1:0] rdata0,
    output reg [DWIDTH-1:0] rdata1
);

    reg [DWIDTH-1:0] mem [0:WORDS-1];

    always @(posedge clk)
    begin
            if (wen)
            begin
                mem[waddr] <= wdata;
            end
            if (backpressure0) rdata0 <= mem[raddr0];
    end


    always @(posedge clk)
    begin
        if (backpressure1) rdata1 <= mem[raddr1];
    end
endmodule




