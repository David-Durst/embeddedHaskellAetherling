module corebit_and (input in0/*verilator public*/, input in1/*verilator public*/, output out/*verilator public*/);
  assign out = in0 & in1;
endmodule

module atomTupleCreator_t0Int_t1Int (input [7:0] I0/*verilator public*/, input [7:0] I1/*verilator public*/, output [7:0] O__0/*verilator public*/, output [7:0] O__1/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
assign O__0 = I0;
assign O__1 = I1;
assign valid_down = valid_up;
endmodule

module coreir_term #(parameter width = 1) (input [width-1:0] in/*verilator public*/);

endmodule

module coreir_reg #(parameter width = 1, parameter clk_posedge = 1, parameter init = 1) (input clk/*verilator public*/, input [width-1:0] in/*verilator public*/, output [width-1:0] out/*verilator public*/);
  reg [width-1:0] outReg/*verilator public*/=init;
  wire real_clk;
  assign real_clk = clk_posedge ? clk : ~clk;
  always @(posedge real_clk) begin
    outReg <= in;
  end
  assign out = outReg;
endmodule

module coreir_const #(parameter width = 1, parameter value = 1) (output [width-1:0] out/*verilator public*/);
  assign out = value;
endmodule

module coreir_add #(parameter width = 1) (input [width-1:0] in0/*verilator public*/, input [width-1:0] in1/*verilator public*/, output [width-1:0] out/*verilator public*/);
  assign out = in0 + in1;
endmodule

module lutN #(parameter N = 1, parameter init = 1) (input [N-1:0] in/*verilator public*/, output out/*verilator public*/);
  assign out = init[in];
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit8200 (input [1599:0] in/*verilator public*/, output [7:0] out_0/*verilator public*/, output [7:0] out_1/*verilator public*/, output [7:0] out_10/*verilator public*/, output [7:0] out_100/*verilator public*/, output [7:0] out_101/*verilator public*/, output [7:0] out_102/*verilator public*/, output [7:0] out_103/*verilator public*/, output [7:0] out_104/*verilator public*/, output [7:0] out_105/*verilator public*/, output [7:0] out_106/*verilator public*/, output [7:0] out_107/*verilator public*/, output [7:0] out_108/*verilator public*/, output [7:0] out_109/*verilator public*/, output [7:0] out_11/*verilator public*/, output [7:0] out_110/*verilator public*/, output [7:0] out_111/*verilator public*/, output [7:0] out_112/*verilator public*/, output [7:0] out_113/*verilator public*/, output [7:0] out_114/*verilator public*/, output [7:0] out_115/*verilator public*/, output [7:0] out_116/*verilator public*/, output [7:0] out_117/*verilator public*/, output [7:0] out_118/*verilator public*/, output [7:0] out_119/*verilator public*/, output [7:0] out_12/*verilator public*/, output [7:0] out_120/*verilator public*/, output [7:0] out_121/*verilator public*/, output [7:0] out_122/*verilator public*/, output [7:0] out_123/*verilator public*/, output [7:0] out_124/*verilator public*/, output [7:0] out_125/*verilator public*/, output [7:0] out_126/*verilator public*/, output [7:0] out_127/*verilator public*/, output [7:0] out_128/*verilator public*/, output [7:0] out_129/*verilator public*/, output [7:0] out_13/*verilator public*/, output [7:0] out_130/*verilator public*/, output [7:0] out_131/*verilator public*/, output [7:0] out_132/*verilator public*/, output [7:0] out_133/*verilator public*/, output [7:0] out_134/*verilator public*/, output [7:0] out_135/*verilator public*/, output [7:0] out_136/*verilator public*/, output [7:0] out_137/*verilator public*/, output [7:0] out_138/*verilator public*/, output [7:0] out_139/*verilator public*/, output [7:0] out_14/*verilator public*/, output [7:0] out_140/*verilator public*/, output [7:0] out_141/*verilator public*/, output [7:0] out_142/*verilator public*/, output [7:0] out_143/*verilator public*/, output [7:0] out_144/*verilator public*/, output [7:0] out_145/*verilator public*/, output [7:0] out_146/*verilator public*/, output [7:0] out_147/*verilator public*/, output [7:0] out_148/*verilator public*/, output [7:0] out_149/*verilator public*/, output [7:0] out_15/*verilator public*/, output [7:0] out_150/*verilator public*/, output [7:0] out_151/*verilator public*/, output [7:0] out_152/*verilator public*/, output [7:0] out_153/*verilator public*/, output [7:0] out_154/*verilator public*/, output [7:0] out_155/*verilator public*/, output [7:0] out_156/*verilator public*/, output [7:0] out_157/*verilator public*/, output [7:0] out_158/*verilator public*/, output [7:0] out_159/*verilator public*/, output [7:0] out_16/*verilator public*/, output [7:0] out_160/*verilator public*/, output [7:0] out_161/*verilator public*/, output [7:0] out_162/*verilator public*/, output [7:0] out_163/*verilator public*/, output [7:0] out_164/*verilator public*/, output [7:0] out_165/*verilator public*/, output [7:0] out_166/*verilator public*/, output [7:0] out_167/*verilator public*/, output [7:0] out_168/*verilator public*/, output [7:0] out_169/*verilator public*/, output [7:0] out_17/*verilator public*/, output [7:0] out_170/*verilator public*/, output [7:0] out_171/*verilator public*/, output [7:0] out_172/*verilator public*/, output [7:0] out_173/*verilator public*/, output [7:0] out_174/*verilator public*/, output [7:0] out_175/*verilator public*/, output [7:0] out_176/*verilator public*/, output [7:0] out_177/*verilator public*/, output [7:0] out_178/*verilator public*/, output [7:0] out_179/*verilator public*/, output [7:0] out_18/*verilator public*/, output [7:0] out_180/*verilator public*/, output [7:0] out_181/*verilator public*/, output [7:0] out_182/*verilator public*/, output [7:0] out_183/*verilator public*/, output [7:0] out_184/*verilator public*/, output [7:0] out_185/*verilator public*/, output [7:0] out_186/*verilator public*/, output [7:0] out_187/*verilator public*/, output [7:0] out_188/*verilator public*/, output [7:0] out_189/*verilator public*/, output [7:0] out_19/*verilator public*/, output [7:0] out_190/*verilator public*/, output [7:0] out_191/*verilator public*/, output [7:0] out_192/*verilator public*/, output [7:0] out_193/*verilator public*/, output [7:0] out_194/*verilator public*/, output [7:0] out_195/*verilator public*/, output [7:0] out_196/*verilator public*/, output [7:0] out_197/*verilator public*/, output [7:0] out_198/*verilator public*/, output [7:0] out_199/*verilator public*/, output [7:0] out_2/*verilator public*/, output [7:0] out_20/*verilator public*/, output [7:0] out_21/*verilator public*/, output [7:0] out_22/*verilator public*/, output [7:0] out_23/*verilator public*/, output [7:0] out_24/*verilator public*/, output [7:0] out_25/*verilator public*/, output [7:0] out_26/*verilator public*/, output [7:0] out_27/*verilator public*/, output [7:0] out_28/*verilator public*/, output [7:0] out_29/*verilator public*/, output [7:0] out_3/*verilator public*/, output [7:0] out_30/*verilator public*/, output [7:0] out_31/*verilator public*/, output [7:0] out_32/*verilator public*/, output [7:0] out_33/*verilator public*/, output [7:0] out_34/*verilator public*/, output [7:0] out_35/*verilator public*/, output [7:0] out_36/*verilator public*/, output [7:0] out_37/*verilator public*/, output [7:0] out_38/*verilator public*/, output [7:0] out_39/*verilator public*/, output [7:0] out_4/*verilator public*/, output [7:0] out_40/*verilator public*/, output [7:0] out_41/*verilator public*/, output [7:0] out_42/*verilator public*/, output [7:0] out_43/*verilator public*/, output [7:0] out_44/*verilator public*/, output [7:0] out_45/*verilator public*/, output [7:0] out_46/*verilator public*/, output [7:0] out_47/*verilator public*/, output [7:0] out_48/*verilator public*/, output [7:0] out_49/*verilator public*/, output [7:0] out_5/*verilator public*/, output [7:0] out_50/*verilator public*/, output [7:0] out_51/*verilator public*/, output [7:0] out_52/*verilator public*/, output [7:0] out_53/*verilator public*/, output [7:0] out_54/*verilator public*/, output [7:0] out_55/*verilator public*/, output [7:0] out_56/*verilator public*/, output [7:0] out_57/*verilator public*/, output [7:0] out_58/*verilator public*/, output [7:0] out_59/*verilator public*/, output [7:0] out_6/*verilator public*/, output [7:0] out_60/*verilator public*/, output [7:0] out_61/*verilator public*/, output [7:0] out_62/*verilator public*/, output [7:0] out_63/*verilator public*/, output [7:0] out_64/*verilator public*/, output [7:0] out_65/*verilator public*/, output [7:0] out_66/*verilator public*/, output [7:0] out_67/*verilator public*/, output [7:0] out_68/*verilator public*/, output [7:0] out_69/*verilator public*/, output [7:0] out_7/*verilator public*/, output [7:0] out_70/*verilator public*/, output [7:0] out_71/*verilator public*/, output [7:0] out_72/*verilator public*/, output [7:0] out_73/*verilator public*/, output [7:0] out_74/*verilator public*/, output [7:0] out_75/*verilator public*/, output [7:0] out_76/*verilator public*/, output [7:0] out_77/*verilator public*/, output [7:0] out_78/*verilator public*/, output [7:0] out_79/*verilator public*/, output [7:0] out_8/*verilator public*/, output [7:0] out_80/*verilator public*/, output [7:0] out_81/*verilator public*/, output [7:0] out_82/*verilator public*/, output [7:0] out_83/*verilator public*/, output [7:0] out_84/*verilator public*/, output [7:0] out_85/*verilator public*/, output [7:0] out_86/*verilator public*/, output [7:0] out_87/*verilator public*/, output [7:0] out_88/*verilator public*/, output [7:0] out_89/*verilator public*/, output [7:0] out_9/*verilator public*/, output [7:0] out_90/*verilator public*/, output [7:0] out_91/*verilator public*/, output [7:0] out_92/*verilator public*/, output [7:0] out_93/*verilator public*/, output [7:0] out_94/*verilator public*/, output [7:0] out_95/*verilator public*/, output [7:0] out_96/*verilator public*/, output [7:0] out_97/*verilator public*/, output [7:0] out_98/*verilator public*/, output [7:0] out_99/*verilator public*/);
assign out_0 = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
assign out_1 = {in[15],in[14],in[13],in[12],in[11],in[10],in[9],in[8]};
assign out_10 = {in[87],in[86],in[85],in[84],in[83],in[82],in[81],in[80]};
assign out_100 = {in[807],in[806],in[805],in[804],in[803],in[802],in[801],in[800]};
assign out_101 = {in[815],in[814],in[813],in[812],in[811],in[810],in[809],in[808]};
assign out_102 = {in[823],in[822],in[821],in[820],in[819],in[818],in[817],in[816]};
assign out_103 = {in[831],in[830],in[829],in[828],in[827],in[826],in[825],in[824]};
assign out_104 = {in[839],in[838],in[837],in[836],in[835],in[834],in[833],in[832]};
assign out_105 = {in[847],in[846],in[845],in[844],in[843],in[842],in[841],in[840]};
assign out_106 = {in[855],in[854],in[853],in[852],in[851],in[850],in[849],in[848]};
assign out_107 = {in[863],in[862],in[861],in[860],in[859],in[858],in[857],in[856]};
assign out_108 = {in[871],in[870],in[869],in[868],in[867],in[866],in[865],in[864]};
assign out_109 = {in[879],in[878],in[877],in[876],in[875],in[874],in[873],in[872]};
assign out_11 = {in[95],in[94],in[93],in[92],in[91],in[90],in[89],in[88]};
assign out_110 = {in[887],in[886],in[885],in[884],in[883],in[882],in[881],in[880]};
assign out_111 = {in[895],in[894],in[893],in[892],in[891],in[890],in[889],in[888]};
assign out_112 = {in[903],in[902],in[901],in[900],in[899],in[898],in[897],in[896]};
assign out_113 = {in[911],in[910],in[909],in[908],in[907],in[906],in[905],in[904]};
assign out_114 = {in[919],in[918],in[917],in[916],in[915],in[914],in[913],in[912]};
assign out_115 = {in[927],in[926],in[925],in[924],in[923],in[922],in[921],in[920]};
assign out_116 = {in[935],in[934],in[933],in[932],in[931],in[930],in[929],in[928]};
assign out_117 = {in[943],in[942],in[941],in[940],in[939],in[938],in[937],in[936]};
assign out_118 = {in[951],in[950],in[949],in[948],in[947],in[946],in[945],in[944]};
assign out_119 = {in[959],in[958],in[957],in[956],in[955],in[954],in[953],in[952]};
assign out_12 = {in[103],in[102],in[101],in[100],in[99],in[98],in[97],in[96]};
assign out_120 = {in[967],in[966],in[965],in[964],in[963],in[962],in[961],in[960]};
assign out_121 = {in[975],in[974],in[973],in[972],in[971],in[970],in[969],in[968]};
assign out_122 = {in[983],in[982],in[981],in[980],in[979],in[978],in[977],in[976]};
assign out_123 = {in[991],in[990],in[989],in[988],in[987],in[986],in[985],in[984]};
assign out_124 = {in[999],in[998],in[997],in[996],in[995],in[994],in[993],in[992]};
assign out_125 = {in[1007],in[1006],in[1005],in[1004],in[1003],in[1002],in[1001],in[1000]};
assign out_126 = {in[1015],in[1014],in[1013],in[1012],in[1011],in[1010],in[1009],in[1008]};
assign out_127 = {in[1023],in[1022],in[1021],in[1020],in[1019],in[1018],in[1017],in[1016]};
assign out_128 = {in[1031],in[1030],in[1029],in[1028],in[1027],in[1026],in[1025],in[1024]};
assign out_129 = {in[1039],in[1038],in[1037],in[1036],in[1035],in[1034],in[1033],in[1032]};
assign out_13 = {in[111],in[110],in[109],in[108],in[107],in[106],in[105],in[104]};
assign out_130 = {in[1047],in[1046],in[1045],in[1044],in[1043],in[1042],in[1041],in[1040]};
assign out_131 = {in[1055],in[1054],in[1053],in[1052],in[1051],in[1050],in[1049],in[1048]};
assign out_132 = {in[1063],in[1062],in[1061],in[1060],in[1059],in[1058],in[1057],in[1056]};
assign out_133 = {in[1071],in[1070],in[1069],in[1068],in[1067],in[1066],in[1065],in[1064]};
assign out_134 = {in[1079],in[1078],in[1077],in[1076],in[1075],in[1074],in[1073],in[1072]};
assign out_135 = {in[1087],in[1086],in[1085],in[1084],in[1083],in[1082],in[1081],in[1080]};
assign out_136 = {in[1095],in[1094],in[1093],in[1092],in[1091],in[1090],in[1089],in[1088]};
assign out_137 = {in[1103],in[1102],in[1101],in[1100],in[1099],in[1098],in[1097],in[1096]};
assign out_138 = {in[1111],in[1110],in[1109],in[1108],in[1107],in[1106],in[1105],in[1104]};
assign out_139 = {in[1119],in[1118],in[1117],in[1116],in[1115],in[1114],in[1113],in[1112]};
assign out_14 = {in[119],in[118],in[117],in[116],in[115],in[114],in[113],in[112]};
assign out_140 = {in[1127],in[1126],in[1125],in[1124],in[1123],in[1122],in[1121],in[1120]};
assign out_141 = {in[1135],in[1134],in[1133],in[1132],in[1131],in[1130],in[1129],in[1128]};
assign out_142 = {in[1143],in[1142],in[1141],in[1140],in[1139],in[1138],in[1137],in[1136]};
assign out_143 = {in[1151],in[1150],in[1149],in[1148],in[1147],in[1146],in[1145],in[1144]};
assign out_144 = {in[1159],in[1158],in[1157],in[1156],in[1155],in[1154],in[1153],in[1152]};
assign out_145 = {in[1167],in[1166],in[1165],in[1164],in[1163],in[1162],in[1161],in[1160]};
assign out_146 = {in[1175],in[1174],in[1173],in[1172],in[1171],in[1170],in[1169],in[1168]};
assign out_147 = {in[1183],in[1182],in[1181],in[1180],in[1179],in[1178],in[1177],in[1176]};
assign out_148 = {in[1191],in[1190],in[1189],in[1188],in[1187],in[1186],in[1185],in[1184]};
assign out_149 = {in[1199],in[1198],in[1197],in[1196],in[1195],in[1194],in[1193],in[1192]};
assign out_15 = {in[127],in[126],in[125],in[124],in[123],in[122],in[121],in[120]};
assign out_150 = {in[1207],in[1206],in[1205],in[1204],in[1203],in[1202],in[1201],in[1200]};
assign out_151 = {in[1215],in[1214],in[1213],in[1212],in[1211],in[1210],in[1209],in[1208]};
assign out_152 = {in[1223],in[1222],in[1221],in[1220],in[1219],in[1218],in[1217],in[1216]};
assign out_153 = {in[1231],in[1230],in[1229],in[1228],in[1227],in[1226],in[1225],in[1224]};
assign out_154 = {in[1239],in[1238],in[1237],in[1236],in[1235],in[1234],in[1233],in[1232]};
assign out_155 = {in[1247],in[1246],in[1245],in[1244],in[1243],in[1242],in[1241],in[1240]};
assign out_156 = {in[1255],in[1254],in[1253],in[1252],in[1251],in[1250],in[1249],in[1248]};
assign out_157 = {in[1263],in[1262],in[1261],in[1260],in[1259],in[1258],in[1257],in[1256]};
assign out_158 = {in[1271],in[1270],in[1269],in[1268],in[1267],in[1266],in[1265],in[1264]};
assign out_159 = {in[1279],in[1278],in[1277],in[1276],in[1275],in[1274],in[1273],in[1272]};
assign out_16 = {in[135],in[134],in[133],in[132],in[131],in[130],in[129],in[128]};
assign out_160 = {in[1287],in[1286],in[1285],in[1284],in[1283],in[1282],in[1281],in[1280]};
assign out_161 = {in[1295],in[1294],in[1293],in[1292],in[1291],in[1290],in[1289],in[1288]};
assign out_162 = {in[1303],in[1302],in[1301],in[1300],in[1299],in[1298],in[1297],in[1296]};
assign out_163 = {in[1311],in[1310],in[1309],in[1308],in[1307],in[1306],in[1305],in[1304]};
assign out_164 = {in[1319],in[1318],in[1317],in[1316],in[1315],in[1314],in[1313],in[1312]};
assign out_165 = {in[1327],in[1326],in[1325],in[1324],in[1323],in[1322],in[1321],in[1320]};
assign out_166 = {in[1335],in[1334],in[1333],in[1332],in[1331],in[1330],in[1329],in[1328]};
assign out_167 = {in[1343],in[1342],in[1341],in[1340],in[1339],in[1338],in[1337],in[1336]};
assign out_168 = {in[1351],in[1350],in[1349],in[1348],in[1347],in[1346],in[1345],in[1344]};
assign out_169 = {in[1359],in[1358],in[1357],in[1356],in[1355],in[1354],in[1353],in[1352]};
assign out_17 = {in[143],in[142],in[141],in[140],in[139],in[138],in[137],in[136]};
assign out_170 = {in[1367],in[1366],in[1365],in[1364],in[1363],in[1362],in[1361],in[1360]};
assign out_171 = {in[1375],in[1374],in[1373],in[1372],in[1371],in[1370],in[1369],in[1368]};
assign out_172 = {in[1383],in[1382],in[1381],in[1380],in[1379],in[1378],in[1377],in[1376]};
assign out_173 = {in[1391],in[1390],in[1389],in[1388],in[1387],in[1386],in[1385],in[1384]};
assign out_174 = {in[1399],in[1398],in[1397],in[1396],in[1395],in[1394],in[1393],in[1392]};
assign out_175 = {in[1407],in[1406],in[1405],in[1404],in[1403],in[1402],in[1401],in[1400]};
assign out_176 = {in[1415],in[1414],in[1413],in[1412],in[1411],in[1410],in[1409],in[1408]};
assign out_177 = {in[1423],in[1422],in[1421],in[1420],in[1419],in[1418],in[1417],in[1416]};
assign out_178 = {in[1431],in[1430],in[1429],in[1428],in[1427],in[1426],in[1425],in[1424]};
assign out_179 = {in[1439],in[1438],in[1437],in[1436],in[1435],in[1434],in[1433],in[1432]};
assign out_18 = {in[151],in[150],in[149],in[148],in[147],in[146],in[145],in[144]};
assign out_180 = {in[1447],in[1446],in[1445],in[1444],in[1443],in[1442],in[1441],in[1440]};
assign out_181 = {in[1455],in[1454],in[1453],in[1452],in[1451],in[1450],in[1449],in[1448]};
assign out_182 = {in[1463],in[1462],in[1461],in[1460],in[1459],in[1458],in[1457],in[1456]};
assign out_183 = {in[1471],in[1470],in[1469],in[1468],in[1467],in[1466],in[1465],in[1464]};
assign out_184 = {in[1479],in[1478],in[1477],in[1476],in[1475],in[1474],in[1473],in[1472]};
assign out_185 = {in[1487],in[1486],in[1485],in[1484],in[1483],in[1482],in[1481],in[1480]};
assign out_186 = {in[1495],in[1494],in[1493],in[1492],in[1491],in[1490],in[1489],in[1488]};
assign out_187 = {in[1503],in[1502],in[1501],in[1500],in[1499],in[1498],in[1497],in[1496]};
assign out_188 = {in[1511],in[1510],in[1509],in[1508],in[1507],in[1506],in[1505],in[1504]};
assign out_189 = {in[1519],in[1518],in[1517],in[1516],in[1515],in[1514],in[1513],in[1512]};
assign out_19 = {in[159],in[158],in[157],in[156],in[155],in[154],in[153],in[152]};
assign out_190 = {in[1527],in[1526],in[1525],in[1524],in[1523],in[1522],in[1521],in[1520]};
assign out_191 = {in[1535],in[1534],in[1533],in[1532],in[1531],in[1530],in[1529],in[1528]};
assign out_192 = {in[1543],in[1542],in[1541],in[1540],in[1539],in[1538],in[1537],in[1536]};
assign out_193 = {in[1551],in[1550],in[1549],in[1548],in[1547],in[1546],in[1545],in[1544]};
assign out_194 = {in[1559],in[1558],in[1557],in[1556],in[1555],in[1554],in[1553],in[1552]};
assign out_195 = {in[1567],in[1566],in[1565],in[1564],in[1563],in[1562],in[1561],in[1560]};
assign out_196 = {in[1575],in[1574],in[1573],in[1572],in[1571],in[1570],in[1569],in[1568]};
assign out_197 = {in[1583],in[1582],in[1581],in[1580],in[1579],in[1578],in[1577],in[1576]};
assign out_198 = {in[1591],in[1590],in[1589],in[1588],in[1587],in[1586],in[1585],in[1584]};
assign out_199 = {in[1599],in[1598],in[1597],in[1596],in[1595],in[1594],in[1593],in[1592]};
assign out_2 = {in[23],in[22],in[21],in[20],in[19],in[18],in[17],in[16]};
assign out_20 = {in[167],in[166],in[165],in[164],in[163],in[162],in[161],in[160]};
assign out_21 = {in[175],in[174],in[173],in[172],in[171],in[170],in[169],in[168]};
assign out_22 = {in[183],in[182],in[181],in[180],in[179],in[178],in[177],in[176]};
assign out_23 = {in[191],in[190],in[189],in[188],in[187],in[186],in[185],in[184]};
assign out_24 = {in[199],in[198],in[197],in[196],in[195],in[194],in[193],in[192]};
assign out_25 = {in[207],in[206],in[205],in[204],in[203],in[202],in[201],in[200]};
assign out_26 = {in[215],in[214],in[213],in[212],in[211],in[210],in[209],in[208]};
assign out_27 = {in[223],in[222],in[221],in[220],in[219],in[218],in[217],in[216]};
assign out_28 = {in[231],in[230],in[229],in[228],in[227],in[226],in[225],in[224]};
assign out_29 = {in[239],in[238],in[237],in[236],in[235],in[234],in[233],in[232]};
assign out_3 = {in[31],in[30],in[29],in[28],in[27],in[26],in[25],in[24]};
assign out_30 = {in[247],in[246],in[245],in[244],in[243],in[242],in[241],in[240]};
assign out_31 = {in[255],in[254],in[253],in[252],in[251],in[250],in[249],in[248]};
assign out_32 = {in[263],in[262],in[261],in[260],in[259],in[258],in[257],in[256]};
assign out_33 = {in[271],in[270],in[269],in[268],in[267],in[266],in[265],in[264]};
assign out_34 = {in[279],in[278],in[277],in[276],in[275],in[274],in[273],in[272]};
assign out_35 = {in[287],in[286],in[285],in[284],in[283],in[282],in[281],in[280]};
assign out_36 = {in[295],in[294],in[293],in[292],in[291],in[290],in[289],in[288]};
assign out_37 = {in[303],in[302],in[301],in[300],in[299],in[298],in[297],in[296]};
assign out_38 = {in[311],in[310],in[309],in[308],in[307],in[306],in[305],in[304]};
assign out_39 = {in[319],in[318],in[317],in[316],in[315],in[314],in[313],in[312]};
assign out_4 = {in[39],in[38],in[37],in[36],in[35],in[34],in[33],in[32]};
assign out_40 = {in[327],in[326],in[325],in[324],in[323],in[322],in[321],in[320]};
assign out_41 = {in[335],in[334],in[333],in[332],in[331],in[330],in[329],in[328]};
assign out_42 = {in[343],in[342],in[341],in[340],in[339],in[338],in[337],in[336]};
assign out_43 = {in[351],in[350],in[349],in[348],in[347],in[346],in[345],in[344]};
assign out_44 = {in[359],in[358],in[357],in[356],in[355],in[354],in[353],in[352]};
assign out_45 = {in[367],in[366],in[365],in[364],in[363],in[362],in[361],in[360]};
assign out_46 = {in[375],in[374],in[373],in[372],in[371],in[370],in[369],in[368]};
assign out_47 = {in[383],in[382],in[381],in[380],in[379],in[378],in[377],in[376]};
assign out_48 = {in[391],in[390],in[389],in[388],in[387],in[386],in[385],in[384]};
assign out_49 = {in[399],in[398],in[397],in[396],in[395],in[394],in[393],in[392]};
assign out_5 = {in[47],in[46],in[45],in[44],in[43],in[42],in[41],in[40]};
assign out_50 = {in[407],in[406],in[405],in[404],in[403],in[402],in[401],in[400]};
assign out_51 = {in[415],in[414],in[413],in[412],in[411],in[410],in[409],in[408]};
assign out_52 = {in[423],in[422],in[421],in[420],in[419],in[418],in[417],in[416]};
assign out_53 = {in[431],in[430],in[429],in[428],in[427],in[426],in[425],in[424]};
assign out_54 = {in[439],in[438],in[437],in[436],in[435],in[434],in[433],in[432]};
assign out_55 = {in[447],in[446],in[445],in[444],in[443],in[442],in[441],in[440]};
assign out_56 = {in[455],in[454],in[453],in[452],in[451],in[450],in[449],in[448]};
assign out_57 = {in[463],in[462],in[461],in[460],in[459],in[458],in[457],in[456]};
assign out_58 = {in[471],in[470],in[469],in[468],in[467],in[466],in[465],in[464]};
assign out_59 = {in[479],in[478],in[477],in[476],in[475],in[474],in[473],in[472]};
assign out_6 = {in[55],in[54],in[53],in[52],in[51],in[50],in[49],in[48]};
assign out_60 = {in[487],in[486],in[485],in[484],in[483],in[482],in[481],in[480]};
assign out_61 = {in[495],in[494],in[493],in[492],in[491],in[490],in[489],in[488]};
assign out_62 = {in[503],in[502],in[501],in[500],in[499],in[498],in[497],in[496]};
assign out_63 = {in[511],in[510],in[509],in[508],in[507],in[506],in[505],in[504]};
assign out_64 = {in[519],in[518],in[517],in[516],in[515],in[514],in[513],in[512]};
assign out_65 = {in[527],in[526],in[525],in[524],in[523],in[522],in[521],in[520]};
assign out_66 = {in[535],in[534],in[533],in[532],in[531],in[530],in[529],in[528]};
assign out_67 = {in[543],in[542],in[541],in[540],in[539],in[538],in[537],in[536]};
assign out_68 = {in[551],in[550],in[549],in[548],in[547],in[546],in[545],in[544]};
assign out_69 = {in[559],in[558],in[557],in[556],in[555],in[554],in[553],in[552]};
assign out_7 = {in[63],in[62],in[61],in[60],in[59],in[58],in[57],in[56]};
assign out_70 = {in[567],in[566],in[565],in[564],in[563],in[562],in[561],in[560]};
assign out_71 = {in[575],in[574],in[573],in[572],in[571],in[570],in[569],in[568]};
assign out_72 = {in[583],in[582],in[581],in[580],in[579],in[578],in[577],in[576]};
assign out_73 = {in[591],in[590],in[589],in[588],in[587],in[586],in[585],in[584]};
assign out_74 = {in[599],in[598],in[597],in[596],in[595],in[594],in[593],in[592]};
assign out_75 = {in[607],in[606],in[605],in[604],in[603],in[602],in[601],in[600]};
assign out_76 = {in[615],in[614],in[613],in[612],in[611],in[610],in[609],in[608]};
assign out_77 = {in[623],in[622],in[621],in[620],in[619],in[618],in[617],in[616]};
assign out_78 = {in[631],in[630],in[629],in[628],in[627],in[626],in[625],in[624]};
assign out_79 = {in[639],in[638],in[637],in[636],in[635],in[634],in[633],in[632]};
assign out_8 = {in[71],in[70],in[69],in[68],in[67],in[66],in[65],in[64]};
assign out_80 = {in[647],in[646],in[645],in[644],in[643],in[642],in[641],in[640]};
assign out_81 = {in[655],in[654],in[653],in[652],in[651],in[650],in[649],in[648]};
assign out_82 = {in[663],in[662],in[661],in[660],in[659],in[658],in[657],in[656]};
assign out_83 = {in[671],in[670],in[669],in[668],in[667],in[666],in[665],in[664]};
assign out_84 = {in[679],in[678],in[677],in[676],in[675],in[674],in[673],in[672]};
assign out_85 = {in[687],in[686],in[685],in[684],in[683],in[682],in[681],in[680]};
assign out_86 = {in[695],in[694],in[693],in[692],in[691],in[690],in[689],in[688]};
assign out_87 = {in[703],in[702],in[701],in[700],in[699],in[698],in[697],in[696]};
assign out_88 = {in[711],in[710],in[709],in[708],in[707],in[706],in[705],in[704]};
assign out_89 = {in[719],in[718],in[717],in[716],in[715],in[714],in[713],in[712]};
assign out_9 = {in[79],in[78],in[77],in[76],in[75],in[74],in[73],in[72]};
assign out_90 = {in[727],in[726],in[725],in[724],in[723],in[722],in[721],in[720]};
assign out_91 = {in[735],in[734],in[733],in[732],in[731],in[730],in[729],in[728]};
assign out_92 = {in[743],in[742],in[741],in[740],in[739],in[738],in[737],in[736]};
assign out_93 = {in[751],in[750],in[749],in[748],in[747],in[746],in[745],in[744]};
assign out_94 = {in[759],in[758],in[757],in[756],in[755],in[754],in[753],in[752]};
assign out_95 = {in[767],in[766],in[765],in[764],in[763],in[762],in[761],in[760]};
assign out_96 = {in[775],in[774],in[773],in[772],in[771],in[770],in[769],in[768]};
assign out_97 = {in[783],in[782],in[781],in[780],in[779],in[778],in[777],in[776]};
assign out_98 = {in[791],in[790],in[789],in[788],in[787],in[786],in[785],in[784]};
assign out_99 = {in[799],in[798],in[797],in[796],in[795],in[794],in[793],in[792]};
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit8 (input [7:0] in/*verilator public*/, output [7:0] out/*verilator public*/);
assign out = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
endmodule

module \aetherlinglib_hydrate__hydratedTypeBit (input [0:0] in/*verilator public*/, output out/*verilator public*/);
assign out = in[0];
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit8200 (input [7:0] in_0/*verilator public*/, input [7:0] in_1/*verilator public*/, input [7:0] in_10/*verilator public*/, input [7:0] in_100/*verilator public*/, input [7:0] in_101/*verilator public*/, input [7:0] in_102/*verilator public*/, input [7:0] in_103/*verilator public*/, input [7:0] in_104/*verilator public*/, input [7:0] in_105/*verilator public*/, input [7:0] in_106/*verilator public*/, input [7:0] in_107/*verilator public*/, input [7:0] in_108/*verilator public*/, input [7:0] in_109/*verilator public*/, input [7:0] in_11/*verilator public*/, input [7:0] in_110/*verilator public*/, input [7:0] in_111/*verilator public*/, input [7:0] in_112/*verilator public*/, input [7:0] in_113/*verilator public*/, input [7:0] in_114/*verilator public*/, input [7:0] in_115/*verilator public*/, input [7:0] in_116/*verilator public*/, input [7:0] in_117/*verilator public*/, input [7:0] in_118/*verilator public*/, input [7:0] in_119/*verilator public*/, input [7:0] in_12/*verilator public*/, input [7:0] in_120/*verilator public*/, input [7:0] in_121/*verilator public*/, input [7:0] in_122/*verilator public*/, input [7:0] in_123/*verilator public*/, input [7:0] in_124/*verilator public*/, input [7:0] in_125/*verilator public*/, input [7:0] in_126/*verilator public*/, input [7:0] in_127/*verilator public*/, input [7:0] in_128/*verilator public*/, input [7:0] in_129/*verilator public*/, input [7:0] in_13/*verilator public*/, input [7:0] in_130/*verilator public*/, input [7:0] in_131/*verilator public*/, input [7:0] in_132/*verilator public*/, input [7:0] in_133/*verilator public*/, input [7:0] in_134/*verilator public*/, input [7:0] in_135/*verilator public*/, input [7:0] in_136/*verilator public*/, input [7:0] in_137/*verilator public*/, input [7:0] in_138/*verilator public*/, input [7:0] in_139/*verilator public*/, input [7:0] in_14/*verilator public*/, input [7:0] in_140/*verilator public*/, input [7:0] in_141/*verilator public*/, input [7:0] in_142/*verilator public*/, input [7:0] in_143/*verilator public*/, input [7:0] in_144/*verilator public*/, input [7:0] in_145/*verilator public*/, input [7:0] in_146/*verilator public*/, input [7:0] in_147/*verilator public*/, input [7:0] in_148/*verilator public*/, input [7:0] in_149/*verilator public*/, input [7:0] in_15/*verilator public*/, input [7:0] in_150/*verilator public*/, input [7:0] in_151/*verilator public*/, input [7:0] in_152/*verilator public*/, input [7:0] in_153/*verilator public*/, input [7:0] in_154/*verilator public*/, input [7:0] in_155/*verilator public*/, input [7:0] in_156/*verilator public*/, input [7:0] in_157/*verilator public*/, input [7:0] in_158/*verilator public*/, input [7:0] in_159/*verilator public*/, input [7:0] in_16/*verilator public*/, input [7:0] in_160/*verilator public*/, input [7:0] in_161/*verilator public*/, input [7:0] in_162/*verilator public*/, input [7:0] in_163/*verilator public*/, input [7:0] in_164/*verilator public*/, input [7:0] in_165/*verilator public*/, input [7:0] in_166/*verilator public*/, input [7:0] in_167/*verilator public*/, input [7:0] in_168/*verilator public*/, input [7:0] in_169/*verilator public*/, input [7:0] in_17/*verilator public*/, input [7:0] in_170/*verilator public*/, input [7:0] in_171/*verilator public*/, input [7:0] in_172/*verilator public*/, input [7:0] in_173/*verilator public*/, input [7:0] in_174/*verilator public*/, input [7:0] in_175/*verilator public*/, input [7:0] in_176/*verilator public*/, input [7:0] in_177/*verilator public*/, input [7:0] in_178/*verilator public*/, input [7:0] in_179/*verilator public*/, input [7:0] in_18/*verilator public*/, input [7:0] in_180/*verilator public*/, input [7:0] in_181/*verilator public*/, input [7:0] in_182/*verilator public*/, input [7:0] in_183/*verilator public*/, input [7:0] in_184/*verilator public*/, input [7:0] in_185/*verilator public*/, input [7:0] in_186/*verilator public*/, input [7:0] in_187/*verilator public*/, input [7:0] in_188/*verilator public*/, input [7:0] in_189/*verilator public*/, input [7:0] in_19/*verilator public*/, input [7:0] in_190/*verilator public*/, input [7:0] in_191/*verilator public*/, input [7:0] in_192/*verilator public*/, input [7:0] in_193/*verilator public*/, input [7:0] in_194/*verilator public*/, input [7:0] in_195/*verilator public*/, input [7:0] in_196/*verilator public*/, input [7:0] in_197/*verilator public*/, input [7:0] in_198/*verilator public*/, input [7:0] in_199/*verilator public*/, input [7:0] in_2/*verilator public*/, input [7:0] in_20/*verilator public*/, input [7:0] in_21/*verilator public*/, input [7:0] in_22/*verilator public*/, input [7:0] in_23/*verilator public*/, input [7:0] in_24/*verilator public*/, input [7:0] in_25/*verilator public*/, input [7:0] in_26/*verilator public*/, input [7:0] in_27/*verilator public*/, input [7:0] in_28/*verilator public*/, input [7:0] in_29/*verilator public*/, input [7:0] in_3/*verilator public*/, input [7:0] in_30/*verilator public*/, input [7:0] in_31/*verilator public*/, input [7:0] in_32/*verilator public*/, input [7:0] in_33/*verilator public*/, input [7:0] in_34/*verilator public*/, input [7:0] in_35/*verilator public*/, input [7:0] in_36/*verilator public*/, input [7:0] in_37/*verilator public*/, input [7:0] in_38/*verilator public*/, input [7:0] in_39/*verilator public*/, input [7:0] in_4/*verilator public*/, input [7:0] in_40/*verilator public*/, input [7:0] in_41/*verilator public*/, input [7:0] in_42/*verilator public*/, input [7:0] in_43/*verilator public*/, input [7:0] in_44/*verilator public*/, input [7:0] in_45/*verilator public*/, input [7:0] in_46/*verilator public*/, input [7:0] in_47/*verilator public*/, input [7:0] in_48/*verilator public*/, input [7:0] in_49/*verilator public*/, input [7:0] in_5/*verilator public*/, input [7:0] in_50/*verilator public*/, input [7:0] in_51/*verilator public*/, input [7:0] in_52/*verilator public*/, input [7:0] in_53/*verilator public*/, input [7:0] in_54/*verilator public*/, input [7:0] in_55/*verilator public*/, input [7:0] in_56/*verilator public*/, input [7:0] in_57/*verilator public*/, input [7:0] in_58/*verilator public*/, input [7:0] in_59/*verilator public*/, input [7:0] in_6/*verilator public*/, input [7:0] in_60/*verilator public*/, input [7:0] in_61/*verilator public*/, input [7:0] in_62/*verilator public*/, input [7:0] in_63/*verilator public*/, input [7:0] in_64/*verilator public*/, input [7:0] in_65/*verilator public*/, input [7:0] in_66/*verilator public*/, input [7:0] in_67/*verilator public*/, input [7:0] in_68/*verilator public*/, input [7:0] in_69/*verilator public*/, input [7:0] in_7/*verilator public*/, input [7:0] in_70/*verilator public*/, input [7:0] in_71/*verilator public*/, input [7:0] in_72/*verilator public*/, input [7:0] in_73/*verilator public*/, input [7:0] in_74/*verilator public*/, input [7:0] in_75/*verilator public*/, input [7:0] in_76/*verilator public*/, input [7:0] in_77/*verilator public*/, input [7:0] in_78/*verilator public*/, input [7:0] in_79/*verilator public*/, input [7:0] in_8/*verilator public*/, input [7:0] in_80/*verilator public*/, input [7:0] in_81/*verilator public*/, input [7:0] in_82/*verilator public*/, input [7:0] in_83/*verilator public*/, input [7:0] in_84/*verilator public*/, input [7:0] in_85/*verilator public*/, input [7:0] in_86/*verilator public*/, input [7:0] in_87/*verilator public*/, input [7:0] in_88/*verilator public*/, input [7:0] in_89/*verilator public*/, input [7:0] in_9/*verilator public*/, input [7:0] in_90/*verilator public*/, input [7:0] in_91/*verilator public*/, input [7:0] in_92/*verilator public*/, input [7:0] in_93/*verilator public*/, input [7:0] in_94/*verilator public*/, input [7:0] in_95/*verilator public*/, input [7:0] in_96/*verilator public*/, input [7:0] in_97/*verilator public*/, input [7:0] in_98/*verilator public*/, input [7:0] in_99/*verilator public*/, output [1599:0] out/*verilator public*/);
assign out = {in_199[7],in_199[6],in_199[5],in_199[4],in_199[3],in_199[2],in_199[1],in_199[0],in_198[7],in_198[6],in_198[5],in_198[4],in_198[3],in_198[2],in_198[1],in_198[0],in_197[7],in_197[6],in_197[5],in_197[4],in_197[3],in_197[2],in_197[1],in_197[0],in_196[7],in_196[6],in_196[5],in_196[4],in_196[3],in_196[2],in_196[1],in_196[0],in_195[7],in_195[6],in_195[5],in_195[4],in_195[3],in_195[2],in_195[1],in_195[0],in_194[7],in_194[6],in_194[5],in_194[4],in_194[3],in_194[2],in_194[1],in_194[0],in_193[7],in_193[6],in_193[5],in_193[4],in_193[3],in_193[2],in_193[1],in_193[0],in_192[7],in_192[6],in_192[5],in_192[4],in_192[3],in_192[2],in_192[1],in_192[0],in_191[7],in_191[6],in_191[5],in_191[4],in_191[3],in_191[2],in_191[1],in_191[0],in_190[7],in_190[6],in_190[5],in_190[4],in_190[3],in_190[2],in_190[1],in_190[0],in_189[7],in_189[6],in_189[5],in_189[4],in_189[3],in_189[2],in_189[1],in_189[0],in_188[7],in_188[6],in_188[5],in_188[4],in_188[3],in_188[2],in_188[1],in_188[0],in_187[7],in_187[6],in_187[5],in_187[4],in_187[3],in_187[2],in_187[1],in_187[0],in_186[7],in_186[6],in_186[5],in_186[4],in_186[3],in_186[2],in_186[1],in_186[0],in_185[7],in_185[6],in_185[5],in_185[4],in_185[3],in_185[2],in_185[1],in_185[0],in_184[7],in_184[6],in_184[5],in_184[4],in_184[3],in_184[2],in_184[1],in_184[0],in_183[7],in_183[6],in_183[5],in_183[4],in_183[3],in_183[2],in_183[1],in_183[0],in_182[7],in_182[6],in_182[5],in_182[4],in_182[3],in_182[2],in_182[1],in_182[0],in_181[7],in_181[6],in_181[5],in_181[4],in_181[3],in_181[2],in_181[1],in_181[0],in_180[7],in_180[6],in_180[5],in_180[4],in_180[3],in_180[2],in_180[1],in_180[0],in_179[7],in_179[6],in_179[5],in_179[4],in_179[3],in_179[2],in_179[1],in_179[0],in_178[7],in_178[6],in_178[5],in_178[4],in_178[3],in_178[2],in_178[1],in_178[0],in_177[7],in_177[6],in_177[5],in_177[4],in_177[3],in_177[2],in_177[1],in_177[0],in_176[7],in_176[6],in_176[5],in_176[4],in_176[3],in_176[2],in_176[1],in_176[0],in_175[7],in_175[6],in_175[5],in_175[4],in_175[3],in_175[2],in_175[1],in_175[0],in_174[7],in_174[6],in_174[5],in_174[4],in_174[3],in_174[2],in_174[1],in_174[0],in_173[7],in_173[6],in_173[5],in_173[4],in_173[3],in_173[2],in_173[1],in_173[0],in_172[7],in_172[6],in_172[5],in_172[4],in_172[3],in_172[2],in_172[1],in_172[0],in_171[7],in_171[6],in_171[5],in_171[4],in_171[3],in_171[2],in_171[1],in_171[0],in_170[7],in_170[6],in_170[5],in_170[4],in_170[3],in_170[2],in_170[1],in_170[0],in_169[7],in_169[6],in_169[5],in_169[4],in_169[3],in_169[2],in_169[1],in_169[0],in_168[7],in_168[6],in_168[5],in_168[4],in_168[3],in_168[2],in_168[1],in_168[0],in_167[7],in_167[6],in_167[5],in_167[4],in_167[3],in_167[2],in_167[1],in_167[0],in_166[7],in_166[6],in_166[5],in_166[4],in_166[3],in_166[2],in_166[1],in_166[0],in_165[7],in_165[6],in_165[5],in_165[4],in_165[3],in_165[2],in_165[1],in_165[0],in_164[7],in_164[6],in_164[5],in_164[4],in_164[3],in_164[2],in_164[1],in_164[0],in_163[7],in_163[6],in_163[5],in_163[4],in_163[3],in_163[2],in_163[1],in_163[0],in_162[7],in_162[6],in_162[5],in_162[4],in_162[3],in_162[2],in_162[1],in_162[0],in_161[7],in_161[6],in_161[5],in_161[4],in_161[3],in_161[2],in_161[1],in_161[0],in_160[7],in_160[6],in_160[5],in_160[4],in_160[3],in_160[2],in_160[1],in_160[0],in_159[7],in_159[6],in_159[5],in_159[4],in_159[3],in_159[2],in_159[1],in_159[0],in_158[7],in_158[6],in_158[5],in_158[4],in_158[3],in_158[2],in_158[1],in_158[0],in_157[7],in_157[6],in_157[5],in_157[4],in_157[3],in_157[2],in_157[1],in_157[0],in_156[7],in_156[6],in_156[5],in_156[4],in_156[3],in_156[2],in_156[1],in_156[0],in_155[7],in_155[6],in_155[5],in_155[4],in_155[3],in_155[2],in_155[1],in_155[0],in_154[7],in_154[6],in_154[5],in_154[4],in_154[3],in_154[2],in_154[1],in_154[0],in_153[7],in_153[6],in_153[5],in_153[4],in_153[3],in_153[2],in_153[1],in_153[0],in_152[7],in_152[6],in_152[5],in_152[4],in_152[3],in_152[2],in_152[1],in_152[0],in_151[7],in_151[6],in_151[5],in_151[4],in_151[3],in_151[2],in_151[1],in_151[0],in_150[7],in_150[6],in_150[5],in_150[4],in_150[3],in_150[2],in_150[1],in_150[0],in_149[7],in_149[6],in_149[5],in_149[4],in_149[3],in_149[2],in_149[1],in_149[0],in_148[7],in_148[6],in_148[5],in_148[4],in_148[3],in_148[2],in_148[1],in_148[0],in_147[7],in_147[6],in_147[5],in_147[4],in_147[3],in_147[2],in_147[1],in_147[0],in_146[7],in_146[6],in_146[5],in_146[4],in_146[3],in_146[2],in_146[1],in_146[0],in_145[7],in_145[6],in_145[5],in_145[4],in_145[3],in_145[2],in_145[1],in_145[0],in_144[7],in_144[6],in_144[5],in_144[4],in_144[3],in_144[2],in_144[1],in_144[0],in_143[7],in_143[6],in_143[5],in_143[4],in_143[3],in_143[2],in_143[1],in_143[0],in_142[7],in_142[6],in_142[5],in_142[4],in_142[3],in_142[2],in_142[1],in_142[0],in_141[7],in_141[6],in_141[5],in_141[4],in_141[3],in_141[2],in_141[1],in_141[0],in_140[7],in_140[6],in_140[5],in_140[4],in_140[3],in_140[2],in_140[1],in_140[0],in_139[7],in_139[6],in_139[5],in_139[4],in_139[3],in_139[2],in_139[1],in_139[0],in_138[7],in_138[6],in_138[5],in_138[4],in_138[3],in_138[2],in_138[1],in_138[0],in_137[7],in_137[6],in_137[5],in_137[4],in_137[3],in_137[2],in_137[1],in_137[0],in_136[7],in_136[6],in_136[5],in_136[4],in_136[3],in_136[2],in_136[1],in_136[0],in_135[7],in_135[6],in_135[5],in_135[4],in_135[3],in_135[2],in_135[1],in_135[0],in_134[7],in_134[6],in_134[5],in_134[4],in_134[3],in_134[2],in_134[1],in_134[0],in_133[7],in_133[6],in_133[5],in_133[4],in_133[3],in_133[2],in_133[1],in_133[0],in_132[7],in_132[6],in_132[5],in_132[4],in_132[3],in_132[2],in_132[1],in_132[0],in_131[7],in_131[6],in_131[5],in_131[4],in_131[3],in_131[2],in_131[1],in_131[0],in_130[7],in_130[6],in_130[5],in_130[4],in_130[3],in_130[2],in_130[1],in_130[0],in_129[7],in_129[6],in_129[5],in_129[4],in_129[3],in_129[2],in_129[1],in_129[0],in_128[7],in_128[6],in_128[5],in_128[4],in_128[3],in_128[2],in_128[1],in_128[0],in_127[7],in_127[6],in_127[5],in_127[4],in_127[3],in_127[2],in_127[1],in_127[0],in_126[7],in_126[6],in_126[5],in_126[4],in_126[3],in_126[2],in_126[1],in_126[0],in_125[7],in_125[6],in_125[5],in_125[4],in_125[3],in_125[2],in_125[1],in_125[0],in_124[7],in_124[6],in_124[5],in_124[4],in_124[3],in_124[2],in_124[1],in_124[0],in_123[7],in_123[6],in_123[5],in_123[4],in_123[3],in_123[2],in_123[1],in_123[0],in_122[7],in_122[6],in_122[5],in_122[4],in_122[3],in_122[2],in_122[1],in_122[0],in_121[7],in_121[6],in_121[5],in_121[4],in_121[3],in_121[2],in_121[1],in_121[0],in_120[7],in_120[6],in_120[5],in_120[4],in_120[3],in_120[2],in_120[1],in_120[0],in_119[7],in_119[6],in_119[5],in_119[4],in_119[3],in_119[2],in_119[1],in_119[0],in_118[7],in_118[6],in_118[5],in_118[4],in_118[3],in_118[2],in_118[1],in_118[0],in_117[7],in_117[6],in_117[5],in_117[4],in_117[3],in_117[2],in_117[1],in_117[0],in_116[7],in_116[6],in_116[5],in_116[4],in_116[3],in_116[2],in_116[1],in_116[0],in_115[7],in_115[6],in_115[5],in_115[4],in_115[3],in_115[2],in_115[1],in_115[0],in_114[7],in_114[6],in_114[5],in_114[4],in_114[3],in_114[2],in_114[1],in_114[0],in_113[7],in_113[6],in_113[5],in_113[4],in_113[3],in_113[2],in_113[1],in_113[0],in_112[7],in_112[6],in_112[5],in_112[4],in_112[3],in_112[2],in_112[1],in_112[0],in_111[7],in_111[6],in_111[5],in_111[4],in_111[3],in_111[2],in_111[1],in_111[0],in_110[7],in_110[6],in_110[5],in_110[4],in_110[3],in_110[2],in_110[1],in_110[0],in_109[7],in_109[6],in_109[5],in_109[4],in_109[3],in_109[2],in_109[1],in_109[0],in_108[7],in_108[6],in_108[5],in_108[4],in_108[3],in_108[2],in_108[1],in_108[0],in_107[7],in_107[6],in_107[5],in_107[4],in_107[3],in_107[2],in_107[1],in_107[0],in_106[7],in_106[6],in_106[5],in_106[4],in_106[3],in_106[2],in_106[1],in_106[0],in_105[7],in_105[6],in_105[5],in_105[4],in_105[3],in_105[2],in_105[1],in_105[0],in_104[7],in_104[6],in_104[5],in_104[4],in_104[3],in_104[2],in_104[1],in_104[0],in_103[7],in_103[6],in_103[5],in_103[4],in_103[3],in_103[2],in_103[1],in_103[0],in_102[7],in_102[6],in_102[5],in_102[4],in_102[3],in_102[2],in_102[1],in_102[0],in_101[7],in_101[6],in_101[5],in_101[4],in_101[3],in_101[2],in_101[1],in_101[0],in_100[7],in_100[6],in_100[5],in_100[4],in_100[3],in_100[2],in_100[1],in_100[0],in_99[7],in_99[6],in_99[5],in_99[4],in_99[3],in_99[2],in_99[1],in_99[0],in_98[7],in_98[6],in_98[5],in_98[4],in_98[3],in_98[2],in_98[1],in_98[0],in_97[7],in_97[6],in_97[5],in_97[4],in_97[3],in_97[2],in_97[1],in_97[0],in_96[7],in_96[6],in_96[5],in_96[4],in_96[3],in_96[2],in_96[1],in_96[0],in_95[7],in_95[6],in_95[5],in_95[4],in_95[3],in_95[2],in_95[1],in_95[0],in_94[7],in_94[6],in_94[5],in_94[4],in_94[3],in_94[2],in_94[1],in_94[0],in_93[7],in_93[6],in_93[5],in_93[4],in_93[3],in_93[2],in_93[1],in_93[0],in_92[7],in_92[6],in_92[5],in_92[4],in_92[3],in_92[2],in_92[1],in_92[0],in_91[7],in_91[6],in_91[5],in_91[4],in_91[3],in_91[2],in_91[1],in_91[0],in_90[7],in_90[6],in_90[5],in_90[4],in_90[3],in_90[2],in_90[1],in_90[0],in_89[7],in_89[6],in_89[5],in_89[4],in_89[3],in_89[2],in_89[1],in_89[0],in_88[7],in_88[6],in_88[5],in_88[4],in_88[3],in_88[2],in_88[1],in_88[0],in_87[7],in_87[6],in_87[5],in_87[4],in_87[3],in_87[2],in_87[1],in_87[0],in_86[7],in_86[6],in_86[5],in_86[4],in_86[3],in_86[2],in_86[1],in_86[0],in_85[7],in_85[6],in_85[5],in_85[4],in_85[3],in_85[2],in_85[1],in_85[0],in_84[7],in_84[6],in_84[5],in_84[4],in_84[3],in_84[2],in_84[1],in_84[0],in_83[7],in_83[6],in_83[5],in_83[4],in_83[3],in_83[2],in_83[1],in_83[0],in_82[7],in_82[6],in_82[5],in_82[4],in_82[3],in_82[2],in_82[1],in_82[0],in_81[7],in_81[6],in_81[5],in_81[4],in_81[3],in_81[2],in_81[1],in_81[0],in_80[7],in_80[6],in_80[5],in_80[4],in_80[3],in_80[2],in_80[1],in_80[0],in_79[7],in_79[6],in_79[5],in_79[4],in_79[3],in_79[2],in_79[1],in_79[0],in_78[7],in_78[6],in_78[5],in_78[4],in_78[3],in_78[2],in_78[1],in_78[0],in_77[7],in_77[6],in_77[5],in_77[4],in_77[3],in_77[2],in_77[1],in_77[0],in_76[7],in_76[6],in_76[5],in_76[4],in_76[3],in_76[2],in_76[1],in_76[0],in_75[7],in_75[6],in_75[5],in_75[4],in_75[3],in_75[2],in_75[1],in_75[0],in_74[7],in_74[6],in_74[5],in_74[4],in_74[3],in_74[2],in_74[1],in_74[0],in_73[7],in_73[6],in_73[5],in_73[4],in_73[3],in_73[2],in_73[1],in_73[0],in_72[7],in_72[6],in_72[5],in_72[4],in_72[3],in_72[2],in_72[1],in_72[0],in_71[7],in_71[6],in_71[5],in_71[4],in_71[3],in_71[2],in_71[1],in_71[0],in_70[7],in_70[6],in_70[5],in_70[4],in_70[3],in_70[2],in_70[1],in_70[0],in_69[7],in_69[6],in_69[5],in_69[4],in_69[3],in_69[2],in_69[1],in_69[0],in_68[7],in_68[6],in_68[5],in_68[4],in_68[3],in_68[2],in_68[1],in_68[0],in_67[7],in_67[6],in_67[5],in_67[4],in_67[3],in_67[2],in_67[1],in_67[0],in_66[7],in_66[6],in_66[5],in_66[4],in_66[3],in_66[2],in_66[1],in_66[0],in_65[7],in_65[6],in_65[5],in_65[4],in_65[3],in_65[2],in_65[1],in_65[0],in_64[7],in_64[6],in_64[5],in_64[4],in_64[3],in_64[2],in_64[1],in_64[0],in_63[7],in_63[6],in_63[5],in_63[4],in_63[3],in_63[2],in_63[1],in_63[0],in_62[7],in_62[6],in_62[5],in_62[4],in_62[3],in_62[2],in_62[1],in_62[0],in_61[7],in_61[6],in_61[5],in_61[4],in_61[3],in_61[2],in_61[1],in_61[0],in_60[7],in_60[6],in_60[5],in_60[4],in_60[3],in_60[2],in_60[1],in_60[0],in_59[7],in_59[6],in_59[5],in_59[4],in_59[3],in_59[2],in_59[1],in_59[0],in_58[7],in_58[6],in_58[5],in_58[4],in_58[3],in_58[2],in_58[1],in_58[0],in_57[7],in_57[6],in_57[5],in_57[4],in_57[3],in_57[2],in_57[1],in_57[0],in_56[7],in_56[6],in_56[5],in_56[4],in_56[3],in_56[2],in_56[1],in_56[0],in_55[7],in_55[6],in_55[5],in_55[4],in_55[3],in_55[2],in_55[1],in_55[0],in_54[7],in_54[6],in_54[5],in_54[4],in_54[3],in_54[2],in_54[1],in_54[0],in_53[7],in_53[6],in_53[5],in_53[4],in_53[3],in_53[2],in_53[1],in_53[0],in_52[7],in_52[6],in_52[5],in_52[4],in_52[3],in_52[2],in_52[1],in_52[0],in_51[7],in_51[6],in_51[5],in_51[4],in_51[3],in_51[2],in_51[1],in_51[0],in_50[7],in_50[6],in_50[5],in_50[4],in_50[3],in_50[2],in_50[1],in_50[0],in_49[7],in_49[6],in_49[5],in_49[4],in_49[3],in_49[2],in_49[1],in_49[0],in_48[7],in_48[6],in_48[5],in_48[4],in_48[3],in_48[2],in_48[1],in_48[0],in_47[7],in_47[6],in_47[5],in_47[4],in_47[3],in_47[2],in_47[1],in_47[0],in_46[7],in_46[6],in_46[5],in_46[4],in_46[3],in_46[2],in_46[1],in_46[0],in_45[7],in_45[6],in_45[5],in_45[4],in_45[3],in_45[2],in_45[1],in_45[0],in_44[7],in_44[6],in_44[5],in_44[4],in_44[3],in_44[2],in_44[1],in_44[0],in_43[7],in_43[6],in_43[5],in_43[4],in_43[3],in_43[2],in_43[1],in_43[0],in_42[7],in_42[6],in_42[5],in_42[4],in_42[3],in_42[2],in_42[1],in_42[0],in_41[7],in_41[6],in_41[5],in_41[4],in_41[3],in_41[2],in_41[1],in_41[0],in_40[7],in_40[6],in_40[5],in_40[4],in_40[3],in_40[2],in_40[1],in_40[0],in_39[7],in_39[6],in_39[5],in_39[4],in_39[3],in_39[2],in_39[1],in_39[0],in_38[7],in_38[6],in_38[5],in_38[4],in_38[3],in_38[2],in_38[1],in_38[0],in_37[7],in_37[6],in_37[5],in_37[4],in_37[3],in_37[2],in_37[1],in_37[0],in_36[7],in_36[6],in_36[5],in_36[4],in_36[3],in_36[2],in_36[1],in_36[0],in_35[7],in_35[6],in_35[5],in_35[4],in_35[3],in_35[2],in_35[1],in_35[0],in_34[7],in_34[6],in_34[5],in_34[4],in_34[3],in_34[2],in_34[1],in_34[0],in_33[7],in_33[6],in_33[5],in_33[4],in_33[3],in_33[2],in_33[1],in_33[0],in_32[7],in_32[6],in_32[5],in_32[4],in_32[3],in_32[2],in_32[1],in_32[0],in_31[7],in_31[6],in_31[5],in_31[4],in_31[3],in_31[2],in_31[1],in_31[0],in_30[7],in_30[6],in_30[5],in_30[4],in_30[3],in_30[2],in_30[1],in_30[0],in_29[7],in_29[6],in_29[5],in_29[4],in_29[3],in_29[2],in_29[1],in_29[0],in_28[7],in_28[6],in_28[5],in_28[4],in_28[3],in_28[2],in_28[1],in_28[0],in_27[7],in_27[6],in_27[5],in_27[4],in_27[3],in_27[2],in_27[1],in_27[0],in_26[7],in_26[6],in_26[5],in_26[4],in_26[3],in_26[2],in_26[1],in_26[0],in_25[7],in_25[6],in_25[5],in_25[4],in_25[3],in_25[2],in_25[1],in_25[0],in_24[7],in_24[6],in_24[5],in_24[4],in_24[3],in_24[2],in_24[1],in_24[0],in_23[7],in_23[6],in_23[5],in_23[4],in_23[3],in_23[2],in_23[1],in_23[0],in_22[7],in_22[6],in_22[5],in_22[4],in_22[3],in_22[2],in_22[1],in_22[0],in_21[7],in_21[6],in_21[5],in_21[4],in_21[3],in_21[2],in_21[1],in_21[0],in_20[7],in_20[6],in_20[5],in_20[4],in_20[3],in_20[2],in_20[1],in_20[0],in_19[7],in_19[6],in_19[5],in_19[4],in_19[3],in_19[2],in_19[1],in_19[0],in_18[7],in_18[6],in_18[5],in_18[4],in_18[3],in_18[2],in_18[1],in_18[0],in_17[7],in_17[6],in_17[5],in_17[4],in_17[3],in_17[2],in_17[1],in_17[0],in_16[7],in_16[6],in_16[5],in_16[4],in_16[3],in_16[2],in_16[1],in_16[0],in_15[7],in_15[6],in_15[5],in_15[4],in_15[3],in_15[2],in_15[1],in_15[0],in_14[7],in_14[6],in_14[5],in_14[4],in_14[3],in_14[2],in_14[1],in_14[0],in_13[7],in_13[6],in_13[5],in_13[4],in_13[3],in_13[2],in_13[1],in_13[0],in_12[7],in_12[6],in_12[5],in_12[4],in_12[3],in_12[2],in_12[1],in_12[0],in_11[7],in_11[6],in_11[5],in_11[4],in_11[3],in_11[2],in_11[1],in_11[0],in_10[7],in_10[6],in_10[5],in_10[4],in_10[3],in_10[2],in_10[1],in_10[0],in_9[7],in_9[6],in_9[5],in_9[4],in_9[3],in_9[2],in_9[1],in_9[0],in_8[7],in_8[6],in_8[5],in_8[4],in_8[3],in_8[2],in_8[1],in_8[0],in_7[7],in_7[6],in_7[5],in_7[4],in_7[3],in_7[2],in_7[1],in_7[0],in_6[7],in_6[6],in_6[5],in_6[4],in_6[3],in_6[2],in_6[1],in_6[0],in_5[7],in_5[6],in_5[5],in_5[4],in_5[3],in_5[2],in_5[1],in_5[0],in_4[7],in_4[6],in_4[5],in_4[4],in_4[3],in_4[2],in_4[1],in_4[0],in_3[7],in_3[6],in_3[5],in_3[4],in_3[3],in_3[2],in_3[1],in_3[0],in_2[7],in_2[6],in_2[5],in_2[4],in_2[3],in_2[2],in_2[1],in_2[0],in_1[7],in_1[6],in_1[5],in_1[4],in_1[3],in_1[2],in_1[1],in_1[0],in_0[7],in_0[6],in_0[5],in_0[4],in_0[3],in_0[2],in_0[1],in_0[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit8 (input [7:0] in/*verilator public*/, output [7:0] out/*verilator public*/);
assign out = {in[7],in[6],in[5],in[4],in[3],in[2],in[1],in[0]};
endmodule

module \aetherlinglib_dehydrate__hydratedTypeBit (input in/*verilator public*/, output [0:0] out/*verilator public*/);
assign out = in;
endmodule

module Term_Bitt (input I/*verilator public*/);
wire [0:0] dehydrate_tBit_inst0_out;
\aetherlinglib_dehydrate__hydratedTypeBit dehydrate_tBit_inst0(.in(I), .out(dehydrate_tBit_inst0_out));
coreir_term #(.width(1)) term_w1_inst0(.in(dehydrate_tBit_inst0_out));
endmodule

module SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse (input CE/*verilator public*/, input CLK/*verilator public*/, output [0:0] O/*verilator public*/);
wire [0:0] const_0_1_out;
Term_Bitt Term_Bitt_inst0(.I(CE));
coreir_const #(.value(1'h0), .width(1)) const_0_1(.out(const_0_1_out));
assign O = const_0_1_out;
endmodule

module LUT1_1 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h1), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT1_0 (input I0/*verilator public*/, output O/*verilator public*/);
wire coreir_lut1_inst0_out;
lutN #(.init(2'h0), .N(1)) coreir_lut1_inst0(.in(I0), .out(coreir_lut1_inst0_out));
assign O = coreir_lut1_inst0_out;
endmodule

module LUT_Array_8_Bit_t_1n (input CLK/*verilator public*/, input [0:0] addr/*verilator public*/, output [7:0] data/*verilator public*/);
wire LUT1_0_inst0_O;
wire LUT1_0_inst1_O;
wire LUT1_0_inst2_O;
wire LUT1_0_inst3_O;
wire LUT1_0_inst4_O;
wire LUT1_0_inst5_O;
wire LUT1_1_inst0_O;
wire LUT1_1_inst1_O;
wire [7:0] hydrate_tArray_8_Bit__inst0_out;
LUT1_0 LUT1_0_inst0(.I0(addr[0]), .O(LUT1_0_inst0_O));
LUT1_0 LUT1_0_inst1(.I0(addr[0]), .O(LUT1_0_inst1_O));
LUT1_0 LUT1_0_inst2(.I0(addr[0]), .O(LUT1_0_inst2_O));
LUT1_0 LUT1_0_inst3(.I0(addr[0]), .O(LUT1_0_inst3_O));
LUT1_0 LUT1_0_inst4(.I0(addr[0]), .O(LUT1_0_inst4_O));
LUT1_0 LUT1_0_inst5(.I0(addr[0]), .O(LUT1_0_inst5_O));
LUT1_1 LUT1_1_inst0(.I0(addr[0]), .O(LUT1_1_inst0_O));
LUT1_1 LUT1_1_inst1(.I0(addr[0]), .O(LUT1_1_inst1_O));
\aetherlinglib_hydrate__hydratedTypeBit8 hydrate_tArray_8_Bit__inst0(.in({LUT1_0_inst5_O,LUT1_0_inst4_O,LUT1_0_inst3_O,LUT1_0_inst2_O,LUT1_0_inst1_O,LUT1_1_inst1_O,LUT1_0_inst0_O,LUT1_1_inst0_O}), .out(hydrate_tArray_8_Bit__inst0_out));
assign data = hydrate_tArray_8_Bit__inst0_out;
endmodule

module DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] reg_P_inst0_out;
coreir_reg #(.clk_posedge(1), .init(1'h0), .width(1)) reg_P_inst0(.clk(CLK), .in(I), .out(reg_P_inst0_out));
assign O = reg_P_inst0_out[0];
endmodule

module Register8 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7(.CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_8_Bit_t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/);
wire [7:0] Register8_inst0_O;
wire [7:0] dehydrate_tArray_8_Bit__inst0_out;
wire [7:0] hydrate_tArray_8_Bit__inst0_out;
Register8 Register8_inst0(.CLK(CLK), .I(dehydrate_tArray_8_Bit__inst0_out), .O(Register8_inst0_O));
\aetherlinglib_dehydrate__hydratedTypeBit8 dehydrate_tArray_8_Bit__inst0(.in(I), .out(dehydrate_tArray_8_Bit__inst0_out));
\aetherlinglib_hydrate__hydratedTypeBit8 hydrate_tArray_8_Bit__inst0(.in(Register8_inst0_O), .out(hydrate_tArray_8_Bit__inst0_out));
assign O = hydrate_tArray_8_Bit__inst0_out;
endmodule

module Register1600 (input CLK/*verilator public*/, input [1599:0] I/*verilator public*/, output [1599:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst100_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1000_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1001_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1002_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1003_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1004_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1005_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1006_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1007_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1008_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1009_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst101_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1010_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1011_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1012_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1013_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1014_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1015_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1016_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1017_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1018_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1019_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst102_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1020_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1021_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1022_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1023_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1024_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1025_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1026_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1027_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1028_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1029_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst103_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1030_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1031_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1032_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1033_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1034_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1035_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1036_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1037_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1038_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1039_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst104_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1040_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1041_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1042_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1043_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1044_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1045_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1046_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1047_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1048_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1049_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst105_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1050_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1051_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1052_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1053_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1054_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1055_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1056_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1057_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1058_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1059_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst106_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1060_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1061_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1062_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1063_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1064_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1065_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1066_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1067_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1068_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1069_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst107_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1070_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1071_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1072_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1073_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1074_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1075_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1076_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1077_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1078_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1079_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst108_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1080_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1081_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1082_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1083_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1084_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1085_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1086_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1087_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1088_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1089_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst109_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1090_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1091_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1092_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1093_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1094_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1095_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1096_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1097_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1098_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1099_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst110_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1100_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1101_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1102_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1103_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1104_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1105_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1106_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1107_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1108_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1109_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst111_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1110_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1111_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1112_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1113_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1114_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1115_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1116_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1117_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1118_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1119_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst112_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1120_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1121_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1122_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1123_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1124_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1125_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1126_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1127_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1128_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1129_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst113_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1130_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1131_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1132_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1133_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1134_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1135_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1136_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1137_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1138_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1139_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst114_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1140_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1141_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1142_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1143_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1144_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1145_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1146_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1147_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1148_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1149_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst115_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1150_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1151_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1152_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1153_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1154_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1155_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1156_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1157_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1158_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1159_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst116_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1160_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1161_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1162_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1163_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1164_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1165_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1166_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1167_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1168_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1169_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst117_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1170_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1171_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1172_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1173_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1174_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1175_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1176_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1177_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1178_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1179_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst118_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1180_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1181_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1182_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1183_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1184_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1185_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1186_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1187_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1188_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1189_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst119_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1190_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1191_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1192_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1193_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1194_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1195_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1196_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1197_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1198_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1199_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst120_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1200_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1201_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1202_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1203_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1204_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1205_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1206_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1207_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1208_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1209_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst121_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1210_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1211_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1212_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1213_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1214_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1215_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1216_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1217_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1218_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1219_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst122_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1220_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1221_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1222_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1223_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1224_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1225_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1226_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1227_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1228_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1229_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst123_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1230_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1231_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1232_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1233_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1234_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1235_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1236_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1237_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1238_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1239_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst124_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1240_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1241_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1242_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1243_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1244_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1245_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1246_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1247_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1248_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1249_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst125_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1250_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1251_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1252_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1253_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1254_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1255_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1256_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1257_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1258_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1259_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst126_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1260_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1261_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1262_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1263_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1264_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1265_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1266_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1267_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1268_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1269_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst127_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1270_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1271_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1272_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1273_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1274_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1275_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1276_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1277_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1278_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1279_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst128_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1280_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1281_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1282_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1283_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1284_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1285_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1286_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1287_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1288_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1289_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst129_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1290_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1291_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1292_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1293_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1294_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1295_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1296_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1297_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1298_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1299_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst130_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1300_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1301_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1302_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1303_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1304_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1305_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1306_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1307_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1308_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1309_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst131_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1310_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1311_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1312_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1313_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1314_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1315_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1316_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1317_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1318_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1319_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst132_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1320_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1321_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1322_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1323_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1324_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1325_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1326_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1327_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1328_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1329_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst133_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1330_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1331_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1332_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1333_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1334_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1335_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1336_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1337_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1338_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1339_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst134_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1340_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1341_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1342_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1343_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1344_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1345_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1346_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1347_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1348_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1349_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst135_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1350_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1351_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1352_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1353_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1354_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1355_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1356_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1357_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1358_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1359_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst136_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1360_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1361_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1362_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1363_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1364_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1365_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1366_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1367_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1368_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1369_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst137_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1370_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1371_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1372_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1373_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1374_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1375_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1376_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1377_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1378_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1379_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst138_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1380_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1381_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1382_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1383_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1384_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1385_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1386_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1387_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1388_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1389_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst139_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1390_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1391_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1392_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1393_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1394_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1395_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1396_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1397_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1398_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1399_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst140_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1400_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1401_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1402_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1403_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1404_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1405_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1406_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1407_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1408_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1409_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst141_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1410_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1411_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1412_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1413_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1414_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1415_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1416_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1417_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1418_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1419_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst142_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1420_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1421_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1422_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1423_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1424_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1425_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1426_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1427_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1428_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1429_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst143_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1430_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1431_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1432_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1433_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1434_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1435_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1436_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1437_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1438_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1439_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst144_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1440_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1441_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1442_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1443_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1444_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1445_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1446_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1447_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1448_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1449_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst145_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1450_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1451_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1452_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1453_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1454_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1455_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1456_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1457_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1458_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1459_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst146_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1460_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1461_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1462_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1463_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1464_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1465_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1466_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1467_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1468_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1469_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst147_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1470_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1471_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1472_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1473_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1474_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1475_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1476_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1477_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1478_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1479_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst148_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1480_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1481_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1482_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1483_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1484_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1485_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1486_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1487_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1488_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1489_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst149_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1490_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1491_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1492_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1493_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1494_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1495_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1496_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1497_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1498_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1499_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst150_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1500_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1501_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1502_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1503_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1504_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1505_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1506_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1507_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1508_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1509_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst151_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1510_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1511_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1512_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1513_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1514_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1515_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1516_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1517_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1518_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1519_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst152_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1520_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1521_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1522_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1523_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1524_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1525_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1526_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1527_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1528_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1529_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst153_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1530_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1531_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1532_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1533_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1534_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1535_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1536_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1537_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1538_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1539_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst154_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1540_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1541_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1542_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1543_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1544_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1545_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1546_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1547_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1548_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1549_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst155_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1550_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1551_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1552_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1553_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1554_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1555_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1556_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1557_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1558_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1559_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst156_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1560_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1561_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1562_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1563_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1564_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1565_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1566_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1567_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1568_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1569_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst157_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1570_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1571_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1572_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1573_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1574_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1575_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1576_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1577_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1578_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1579_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst158_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1580_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1581_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1582_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1583_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1584_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1585_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1586_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1587_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1588_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1589_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst159_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1590_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1591_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1592_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1593_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1594_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1595_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1596_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1597_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1598_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1599_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst160_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst161_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst162_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst163_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst164_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst165_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst166_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst167_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst168_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst169_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst170_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst171_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst172_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst173_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst174_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst175_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst176_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst177_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst178_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst179_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst180_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst181_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst182_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst183_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst184_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst185_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst186_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst187_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst188_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst189_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst190_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst191_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst192_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst193_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst194_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst195_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst196_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst197_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst198_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst199_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst200_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst201_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst202_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst203_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst204_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst205_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst206_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst207_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst208_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst209_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst210_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst211_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst212_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst213_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst214_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst215_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst216_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst217_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst218_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst219_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst220_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst221_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst222_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst223_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst224_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst225_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst226_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst227_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst228_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst229_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst230_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst231_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst232_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst233_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst234_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst235_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst236_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst237_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst238_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst239_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst240_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst241_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst242_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst243_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst244_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst245_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst246_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst247_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst248_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst249_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst250_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst251_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst252_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst253_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst254_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst255_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst256_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst257_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst258_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst259_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst260_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst261_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst262_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst263_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst264_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst265_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst266_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst267_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst268_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst269_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst270_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst271_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst272_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst273_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst274_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst275_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst276_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst277_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst278_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst279_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst280_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst281_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst282_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst283_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst284_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst285_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst286_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst287_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst288_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst289_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst290_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst291_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst292_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst293_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst294_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst295_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst296_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst297_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst298_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst299_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst300_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst301_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst302_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst303_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst304_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst305_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst306_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst307_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst308_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst309_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst310_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst311_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst312_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst313_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst314_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst315_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst316_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst317_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst318_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst319_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst32_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst320_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst321_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst322_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst323_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst324_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst325_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst326_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst327_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst328_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst329_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst33_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst330_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst331_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst332_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst333_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst334_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst335_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst336_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst337_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst338_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst339_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst34_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst340_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst341_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst342_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst343_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst344_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst345_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst346_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst347_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst348_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst349_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst35_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst350_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst351_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst352_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst353_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst354_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst355_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst356_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst357_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst358_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst359_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst36_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst360_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst361_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst362_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst363_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst364_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst365_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst366_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst367_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst368_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst369_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst37_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst370_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst371_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst372_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst373_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst374_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst375_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst376_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst377_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst378_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst379_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst38_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst380_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst381_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst382_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst383_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst384_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst385_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst386_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst387_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst388_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst389_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst39_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst390_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst391_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst392_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst393_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst394_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst395_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst396_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst397_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst398_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst399_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst40_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst400_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst401_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst402_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst403_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst404_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst405_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst406_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst407_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst408_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst409_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst41_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst410_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst411_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst412_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst413_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst414_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst415_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst416_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst417_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst418_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst419_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst42_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst420_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst421_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst422_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst423_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst424_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst425_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst426_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst427_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst428_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst429_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst43_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst430_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst431_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst432_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst433_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst434_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst435_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst436_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst437_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst438_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst439_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst44_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst440_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst441_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst442_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst443_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst444_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst445_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst446_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst447_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst448_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst449_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst45_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst450_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst451_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst452_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst453_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst454_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst455_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst456_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst457_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst458_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst459_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst46_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst460_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst461_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst462_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst463_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst464_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst465_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst466_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst467_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst468_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst469_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst47_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst470_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst471_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst472_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst473_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst474_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst475_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst476_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst477_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst478_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst479_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst48_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst480_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst481_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst482_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst483_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst484_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst485_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst486_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst487_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst488_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst489_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst49_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst490_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst491_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst492_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst493_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst494_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst495_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst496_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst497_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst498_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst499_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst50_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst500_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst501_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst502_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst503_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst504_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst505_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst506_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst507_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst508_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst509_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst51_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst510_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst511_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst512_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst513_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst514_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst515_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst516_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst517_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst518_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst519_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst52_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst520_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst521_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst522_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst523_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst524_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst525_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst526_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst527_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst528_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst529_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst53_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst530_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst531_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst532_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst533_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst534_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst535_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst536_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst537_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst538_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst539_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst54_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst540_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst541_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst542_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst543_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst544_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst545_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst546_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst547_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst548_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst549_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst55_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst550_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst551_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst552_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst553_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst554_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst555_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst556_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst557_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst558_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst559_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst56_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst560_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst561_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst562_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst563_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst564_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst565_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst566_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst567_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst568_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst569_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst57_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst570_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst571_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst572_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst573_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst574_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst575_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst576_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst577_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst578_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst579_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst58_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst580_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst581_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst582_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst583_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst584_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst585_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst586_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst587_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst588_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst589_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst59_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst590_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst591_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst592_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst593_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst594_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst595_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst596_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst597_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst598_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst599_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst60_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst600_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst601_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst602_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst603_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst604_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst605_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst606_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst607_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst608_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst609_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst61_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst610_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst611_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst612_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst613_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst614_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst615_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst616_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst617_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst618_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst619_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst62_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst620_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst621_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst622_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst623_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst624_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst625_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst626_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst627_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst628_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst629_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst63_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst630_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst631_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst632_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst633_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst634_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst635_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst636_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst637_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst638_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst639_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst64_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst640_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst641_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst642_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst643_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst644_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst645_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst646_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst647_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst648_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst649_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst65_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst650_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst651_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst652_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst653_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst654_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst655_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst656_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst657_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst658_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst659_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst66_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst660_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst661_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst662_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst663_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst664_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst665_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst666_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst667_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst668_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst669_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst67_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst670_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst671_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst672_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst673_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst674_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst675_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst676_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst677_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst678_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst679_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst68_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst680_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst681_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst682_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst683_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst684_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst685_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst686_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst687_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst688_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst689_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst69_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst690_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst691_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst692_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst693_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst694_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst695_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst696_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst697_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst698_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst699_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst70_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst700_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst701_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst702_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst703_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst704_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst705_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst706_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst707_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst708_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst709_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst71_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst710_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst711_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst712_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst713_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst714_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst715_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst716_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst717_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst718_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst719_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst72_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst720_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst721_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst722_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst723_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst724_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst725_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst726_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst727_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst728_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst729_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst73_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst730_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst731_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst732_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst733_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst734_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst735_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst736_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst737_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst738_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst739_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst74_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst740_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst741_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst742_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst743_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst744_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst745_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst746_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst747_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst748_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst749_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst75_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst750_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst751_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst752_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst753_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst754_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst755_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst756_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst757_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst758_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst759_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst76_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst760_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst761_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst762_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst763_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst764_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst765_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst766_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst767_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst768_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst769_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst77_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst770_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst771_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst772_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst773_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst774_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst775_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst776_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst777_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst778_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst779_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst78_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst780_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst781_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst782_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst783_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst784_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst785_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst786_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst787_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst788_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst789_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst79_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst790_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst791_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst792_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst793_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst794_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst795_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst796_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst797_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst798_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst799_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst80_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst800_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst801_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst802_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst803_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst804_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst805_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst806_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst807_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst808_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst809_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst81_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst810_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst811_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst812_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst813_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst814_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst815_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst816_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst817_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst818_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst819_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst82_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst820_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst821_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst822_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst823_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst824_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst825_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst826_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst827_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst828_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst829_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst83_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst830_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst831_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst832_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst833_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst834_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst835_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst836_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst837_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst838_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst839_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst84_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst840_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst841_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst842_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst843_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst844_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst845_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst846_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst847_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst848_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst849_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst85_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst850_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst851_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst852_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst853_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst854_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst855_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst856_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst857_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst858_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst859_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst86_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst860_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst861_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst862_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst863_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst864_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst865_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst866_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst867_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst868_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst869_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst87_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst870_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst871_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst872_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst873_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst874_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst875_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst876_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst877_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst878_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst879_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst88_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst880_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst881_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst882_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst883_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst884_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst885_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst886_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst887_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst888_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst889_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst89_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst890_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst891_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst892_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst893_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst894_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst895_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst896_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst897_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst898_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst899_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst90_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst900_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst901_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst902_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst903_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst904_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst905_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst906_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst907_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst908_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst909_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst91_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst910_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst911_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst912_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst913_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst914_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst915_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst916_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst917_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst918_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst919_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst92_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst920_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst921_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst922_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst923_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst924_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst925_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst926_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst927_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst928_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst929_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst93_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst930_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst931_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst932_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst933_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst934_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst935_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst936_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst937_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst938_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst939_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst94_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst940_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst941_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst942_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst943_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst944_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst945_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst946_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst947_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst948_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst949_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst95_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst950_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst951_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst952_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst953_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst954_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst955_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst956_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst957_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst958_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst959_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst96_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst960_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst961_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst962_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst963_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst964_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst965_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst966_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst967_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst968_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst969_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst97_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst970_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst971_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst972_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst973_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst974_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst975_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst976_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst977_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst978_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst979_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst98_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst980_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst981_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst982_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst983_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst984_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst985_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst986_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst987_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst988_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst989_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst99_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst990_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst991_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst992_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst993_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst994_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst995_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst996_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst997_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst998_O;
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst999_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1(.CLK(CLK), .I(I[1]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10(.CLK(CLK), .I(I[10]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst100(.CLK(CLK), .I(I[100]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst100_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1000(.CLK(CLK), .I(I[1000]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1000_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1001(.CLK(CLK), .I(I[1001]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1001_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1002(.CLK(CLK), .I(I[1002]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1002_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1003(.CLK(CLK), .I(I[1003]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1003_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1004(.CLK(CLK), .I(I[1004]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1004_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1005(.CLK(CLK), .I(I[1005]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1005_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1006(.CLK(CLK), .I(I[1006]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1006_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1007(.CLK(CLK), .I(I[1007]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1007_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1008(.CLK(CLK), .I(I[1008]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1008_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1009(.CLK(CLK), .I(I[1009]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1009_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst101(.CLK(CLK), .I(I[101]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst101_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1010(.CLK(CLK), .I(I[1010]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1010_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1011(.CLK(CLK), .I(I[1011]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1011_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1012(.CLK(CLK), .I(I[1012]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1012_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1013(.CLK(CLK), .I(I[1013]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1013_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1014(.CLK(CLK), .I(I[1014]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1014_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1015(.CLK(CLK), .I(I[1015]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1015_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1016(.CLK(CLK), .I(I[1016]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1016_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1017(.CLK(CLK), .I(I[1017]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1017_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1018(.CLK(CLK), .I(I[1018]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1018_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1019(.CLK(CLK), .I(I[1019]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1019_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst102(.CLK(CLK), .I(I[102]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst102_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1020(.CLK(CLK), .I(I[1020]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1020_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1021(.CLK(CLK), .I(I[1021]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1021_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1022(.CLK(CLK), .I(I[1022]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1022_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1023(.CLK(CLK), .I(I[1023]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1023_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1024(.CLK(CLK), .I(I[1024]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1024_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1025(.CLK(CLK), .I(I[1025]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1025_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1026(.CLK(CLK), .I(I[1026]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1026_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1027(.CLK(CLK), .I(I[1027]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1027_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1028(.CLK(CLK), .I(I[1028]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1028_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1029(.CLK(CLK), .I(I[1029]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1029_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst103(.CLK(CLK), .I(I[103]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst103_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1030(.CLK(CLK), .I(I[1030]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1030_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1031(.CLK(CLK), .I(I[1031]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1031_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1032(.CLK(CLK), .I(I[1032]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1032_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1033(.CLK(CLK), .I(I[1033]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1033_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1034(.CLK(CLK), .I(I[1034]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1034_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1035(.CLK(CLK), .I(I[1035]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1035_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1036(.CLK(CLK), .I(I[1036]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1036_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1037(.CLK(CLK), .I(I[1037]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1037_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1038(.CLK(CLK), .I(I[1038]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1038_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1039(.CLK(CLK), .I(I[1039]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1039_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst104(.CLK(CLK), .I(I[104]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst104_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1040(.CLK(CLK), .I(I[1040]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1040_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1041(.CLK(CLK), .I(I[1041]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1041_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1042(.CLK(CLK), .I(I[1042]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1042_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1043(.CLK(CLK), .I(I[1043]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1043_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1044(.CLK(CLK), .I(I[1044]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1044_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1045(.CLK(CLK), .I(I[1045]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1045_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1046(.CLK(CLK), .I(I[1046]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1046_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1047(.CLK(CLK), .I(I[1047]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1047_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1048(.CLK(CLK), .I(I[1048]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1048_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1049(.CLK(CLK), .I(I[1049]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1049_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst105(.CLK(CLK), .I(I[105]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst105_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1050(.CLK(CLK), .I(I[1050]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1050_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1051(.CLK(CLK), .I(I[1051]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1051_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1052(.CLK(CLK), .I(I[1052]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1052_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1053(.CLK(CLK), .I(I[1053]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1053_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1054(.CLK(CLK), .I(I[1054]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1054_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1055(.CLK(CLK), .I(I[1055]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1055_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1056(.CLK(CLK), .I(I[1056]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1056_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1057(.CLK(CLK), .I(I[1057]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1057_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1058(.CLK(CLK), .I(I[1058]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1058_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1059(.CLK(CLK), .I(I[1059]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1059_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst106(.CLK(CLK), .I(I[106]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst106_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1060(.CLK(CLK), .I(I[1060]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1060_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1061(.CLK(CLK), .I(I[1061]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1061_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1062(.CLK(CLK), .I(I[1062]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1062_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1063(.CLK(CLK), .I(I[1063]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1063_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1064(.CLK(CLK), .I(I[1064]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1064_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1065(.CLK(CLK), .I(I[1065]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1065_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1066(.CLK(CLK), .I(I[1066]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1066_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1067(.CLK(CLK), .I(I[1067]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1067_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1068(.CLK(CLK), .I(I[1068]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1068_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1069(.CLK(CLK), .I(I[1069]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1069_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst107(.CLK(CLK), .I(I[107]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst107_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1070(.CLK(CLK), .I(I[1070]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1070_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1071(.CLK(CLK), .I(I[1071]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1071_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1072(.CLK(CLK), .I(I[1072]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1072_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1073(.CLK(CLK), .I(I[1073]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1073_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1074(.CLK(CLK), .I(I[1074]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1074_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1075(.CLK(CLK), .I(I[1075]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1075_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1076(.CLK(CLK), .I(I[1076]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1076_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1077(.CLK(CLK), .I(I[1077]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1077_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1078(.CLK(CLK), .I(I[1078]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1078_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1079(.CLK(CLK), .I(I[1079]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1079_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst108(.CLK(CLK), .I(I[108]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst108_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1080(.CLK(CLK), .I(I[1080]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1080_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1081(.CLK(CLK), .I(I[1081]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1081_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1082(.CLK(CLK), .I(I[1082]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1082_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1083(.CLK(CLK), .I(I[1083]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1083_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1084(.CLK(CLK), .I(I[1084]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1084_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1085(.CLK(CLK), .I(I[1085]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1085_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1086(.CLK(CLK), .I(I[1086]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1086_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1087(.CLK(CLK), .I(I[1087]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1087_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1088(.CLK(CLK), .I(I[1088]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1088_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1089(.CLK(CLK), .I(I[1089]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1089_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst109(.CLK(CLK), .I(I[109]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst109_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1090(.CLK(CLK), .I(I[1090]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1090_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1091(.CLK(CLK), .I(I[1091]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1091_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1092(.CLK(CLK), .I(I[1092]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1092_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1093(.CLK(CLK), .I(I[1093]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1093_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1094(.CLK(CLK), .I(I[1094]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1094_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1095(.CLK(CLK), .I(I[1095]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1095_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1096(.CLK(CLK), .I(I[1096]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1096_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1097(.CLK(CLK), .I(I[1097]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1097_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1098(.CLK(CLK), .I(I[1098]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1098_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1099(.CLK(CLK), .I(I[1099]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1099_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11(.CLK(CLK), .I(I[11]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst110(.CLK(CLK), .I(I[110]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst110_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1100(.CLK(CLK), .I(I[1100]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1100_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1101(.CLK(CLK), .I(I[1101]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1101_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1102(.CLK(CLK), .I(I[1102]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1102_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1103(.CLK(CLK), .I(I[1103]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1103_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1104(.CLK(CLK), .I(I[1104]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1104_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1105(.CLK(CLK), .I(I[1105]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1105_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1106(.CLK(CLK), .I(I[1106]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1106_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1107(.CLK(CLK), .I(I[1107]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1107_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1108(.CLK(CLK), .I(I[1108]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1108_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1109(.CLK(CLK), .I(I[1109]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1109_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst111(.CLK(CLK), .I(I[111]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst111_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1110(.CLK(CLK), .I(I[1110]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1110_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1111(.CLK(CLK), .I(I[1111]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1111_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1112(.CLK(CLK), .I(I[1112]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1112_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1113(.CLK(CLK), .I(I[1113]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1113_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1114(.CLK(CLK), .I(I[1114]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1114_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1115(.CLK(CLK), .I(I[1115]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1115_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1116(.CLK(CLK), .I(I[1116]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1116_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1117(.CLK(CLK), .I(I[1117]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1117_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1118(.CLK(CLK), .I(I[1118]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1118_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1119(.CLK(CLK), .I(I[1119]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1119_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst112(.CLK(CLK), .I(I[112]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst112_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1120(.CLK(CLK), .I(I[1120]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1120_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1121(.CLK(CLK), .I(I[1121]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1121_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1122(.CLK(CLK), .I(I[1122]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1122_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1123(.CLK(CLK), .I(I[1123]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1123_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1124(.CLK(CLK), .I(I[1124]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1124_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1125(.CLK(CLK), .I(I[1125]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1125_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1126(.CLK(CLK), .I(I[1126]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1126_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1127(.CLK(CLK), .I(I[1127]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1127_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1128(.CLK(CLK), .I(I[1128]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1128_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1129(.CLK(CLK), .I(I[1129]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1129_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst113(.CLK(CLK), .I(I[113]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst113_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1130(.CLK(CLK), .I(I[1130]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1130_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1131(.CLK(CLK), .I(I[1131]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1131_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1132(.CLK(CLK), .I(I[1132]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1132_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1133(.CLK(CLK), .I(I[1133]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1133_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1134(.CLK(CLK), .I(I[1134]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1134_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1135(.CLK(CLK), .I(I[1135]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1135_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1136(.CLK(CLK), .I(I[1136]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1136_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1137(.CLK(CLK), .I(I[1137]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1137_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1138(.CLK(CLK), .I(I[1138]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1138_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1139(.CLK(CLK), .I(I[1139]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1139_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst114(.CLK(CLK), .I(I[114]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst114_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1140(.CLK(CLK), .I(I[1140]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1140_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1141(.CLK(CLK), .I(I[1141]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1141_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1142(.CLK(CLK), .I(I[1142]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1142_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1143(.CLK(CLK), .I(I[1143]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1143_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1144(.CLK(CLK), .I(I[1144]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1144_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1145(.CLK(CLK), .I(I[1145]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1145_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1146(.CLK(CLK), .I(I[1146]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1146_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1147(.CLK(CLK), .I(I[1147]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1147_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1148(.CLK(CLK), .I(I[1148]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1148_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1149(.CLK(CLK), .I(I[1149]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1149_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst115(.CLK(CLK), .I(I[115]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst115_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1150(.CLK(CLK), .I(I[1150]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1150_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1151(.CLK(CLK), .I(I[1151]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1151_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1152(.CLK(CLK), .I(I[1152]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1152_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1153(.CLK(CLK), .I(I[1153]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1153_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1154(.CLK(CLK), .I(I[1154]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1154_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1155(.CLK(CLK), .I(I[1155]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1155_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1156(.CLK(CLK), .I(I[1156]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1156_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1157(.CLK(CLK), .I(I[1157]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1157_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1158(.CLK(CLK), .I(I[1158]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1158_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1159(.CLK(CLK), .I(I[1159]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1159_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst116(.CLK(CLK), .I(I[116]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst116_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1160(.CLK(CLK), .I(I[1160]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1160_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1161(.CLK(CLK), .I(I[1161]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1161_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1162(.CLK(CLK), .I(I[1162]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1162_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1163(.CLK(CLK), .I(I[1163]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1163_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1164(.CLK(CLK), .I(I[1164]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1164_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1165(.CLK(CLK), .I(I[1165]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1165_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1166(.CLK(CLK), .I(I[1166]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1166_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1167(.CLK(CLK), .I(I[1167]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1167_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1168(.CLK(CLK), .I(I[1168]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1168_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1169(.CLK(CLK), .I(I[1169]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1169_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst117(.CLK(CLK), .I(I[117]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst117_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1170(.CLK(CLK), .I(I[1170]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1170_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1171(.CLK(CLK), .I(I[1171]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1171_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1172(.CLK(CLK), .I(I[1172]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1172_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1173(.CLK(CLK), .I(I[1173]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1173_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1174(.CLK(CLK), .I(I[1174]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1174_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1175(.CLK(CLK), .I(I[1175]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1175_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1176(.CLK(CLK), .I(I[1176]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1176_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1177(.CLK(CLK), .I(I[1177]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1177_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1178(.CLK(CLK), .I(I[1178]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1178_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1179(.CLK(CLK), .I(I[1179]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1179_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst118(.CLK(CLK), .I(I[118]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst118_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1180(.CLK(CLK), .I(I[1180]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1180_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1181(.CLK(CLK), .I(I[1181]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1181_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1182(.CLK(CLK), .I(I[1182]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1182_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1183(.CLK(CLK), .I(I[1183]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1183_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1184(.CLK(CLK), .I(I[1184]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1184_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1185(.CLK(CLK), .I(I[1185]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1185_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1186(.CLK(CLK), .I(I[1186]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1186_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1187(.CLK(CLK), .I(I[1187]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1187_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1188(.CLK(CLK), .I(I[1188]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1188_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1189(.CLK(CLK), .I(I[1189]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1189_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst119(.CLK(CLK), .I(I[119]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst119_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1190(.CLK(CLK), .I(I[1190]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1190_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1191(.CLK(CLK), .I(I[1191]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1191_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1192(.CLK(CLK), .I(I[1192]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1192_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1193(.CLK(CLK), .I(I[1193]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1193_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1194(.CLK(CLK), .I(I[1194]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1194_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1195(.CLK(CLK), .I(I[1195]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1195_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1196(.CLK(CLK), .I(I[1196]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1196_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1197(.CLK(CLK), .I(I[1197]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1197_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1198(.CLK(CLK), .I(I[1198]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1198_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1199(.CLK(CLK), .I(I[1199]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1199_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12(.CLK(CLK), .I(I[12]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst120(.CLK(CLK), .I(I[120]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst120_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1200(.CLK(CLK), .I(I[1200]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1200_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1201(.CLK(CLK), .I(I[1201]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1201_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1202(.CLK(CLK), .I(I[1202]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1202_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1203(.CLK(CLK), .I(I[1203]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1203_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1204(.CLK(CLK), .I(I[1204]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1204_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1205(.CLK(CLK), .I(I[1205]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1205_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1206(.CLK(CLK), .I(I[1206]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1206_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1207(.CLK(CLK), .I(I[1207]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1207_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1208(.CLK(CLK), .I(I[1208]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1208_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1209(.CLK(CLK), .I(I[1209]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1209_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst121(.CLK(CLK), .I(I[121]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst121_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1210(.CLK(CLK), .I(I[1210]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1210_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1211(.CLK(CLK), .I(I[1211]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1211_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1212(.CLK(CLK), .I(I[1212]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1212_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1213(.CLK(CLK), .I(I[1213]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1213_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1214(.CLK(CLK), .I(I[1214]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1214_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1215(.CLK(CLK), .I(I[1215]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1215_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1216(.CLK(CLK), .I(I[1216]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1216_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1217(.CLK(CLK), .I(I[1217]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1217_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1218(.CLK(CLK), .I(I[1218]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1218_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1219(.CLK(CLK), .I(I[1219]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1219_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst122(.CLK(CLK), .I(I[122]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst122_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1220(.CLK(CLK), .I(I[1220]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1220_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1221(.CLK(CLK), .I(I[1221]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1221_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1222(.CLK(CLK), .I(I[1222]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1222_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1223(.CLK(CLK), .I(I[1223]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1223_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1224(.CLK(CLK), .I(I[1224]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1224_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1225(.CLK(CLK), .I(I[1225]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1225_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1226(.CLK(CLK), .I(I[1226]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1226_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1227(.CLK(CLK), .I(I[1227]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1227_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1228(.CLK(CLK), .I(I[1228]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1228_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1229(.CLK(CLK), .I(I[1229]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1229_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst123(.CLK(CLK), .I(I[123]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst123_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1230(.CLK(CLK), .I(I[1230]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1230_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1231(.CLK(CLK), .I(I[1231]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1231_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1232(.CLK(CLK), .I(I[1232]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1232_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1233(.CLK(CLK), .I(I[1233]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1233_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1234(.CLK(CLK), .I(I[1234]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1234_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1235(.CLK(CLK), .I(I[1235]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1235_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1236(.CLK(CLK), .I(I[1236]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1236_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1237(.CLK(CLK), .I(I[1237]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1237_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1238(.CLK(CLK), .I(I[1238]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1238_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1239(.CLK(CLK), .I(I[1239]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1239_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst124(.CLK(CLK), .I(I[124]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst124_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1240(.CLK(CLK), .I(I[1240]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1240_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1241(.CLK(CLK), .I(I[1241]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1241_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1242(.CLK(CLK), .I(I[1242]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1242_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1243(.CLK(CLK), .I(I[1243]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1243_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1244(.CLK(CLK), .I(I[1244]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1244_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1245(.CLK(CLK), .I(I[1245]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1245_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1246(.CLK(CLK), .I(I[1246]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1246_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1247(.CLK(CLK), .I(I[1247]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1247_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1248(.CLK(CLK), .I(I[1248]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1248_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1249(.CLK(CLK), .I(I[1249]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1249_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst125(.CLK(CLK), .I(I[125]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst125_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1250(.CLK(CLK), .I(I[1250]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1250_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1251(.CLK(CLK), .I(I[1251]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1251_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1252(.CLK(CLK), .I(I[1252]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1252_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1253(.CLK(CLK), .I(I[1253]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1253_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1254(.CLK(CLK), .I(I[1254]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1254_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1255(.CLK(CLK), .I(I[1255]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1255_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1256(.CLK(CLK), .I(I[1256]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1256_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1257(.CLK(CLK), .I(I[1257]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1257_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1258(.CLK(CLK), .I(I[1258]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1258_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1259(.CLK(CLK), .I(I[1259]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1259_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst126(.CLK(CLK), .I(I[126]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst126_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1260(.CLK(CLK), .I(I[1260]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1260_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1261(.CLK(CLK), .I(I[1261]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1261_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1262(.CLK(CLK), .I(I[1262]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1262_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1263(.CLK(CLK), .I(I[1263]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1263_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1264(.CLK(CLK), .I(I[1264]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1264_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1265(.CLK(CLK), .I(I[1265]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1265_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1266(.CLK(CLK), .I(I[1266]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1266_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1267(.CLK(CLK), .I(I[1267]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1267_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1268(.CLK(CLK), .I(I[1268]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1268_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1269(.CLK(CLK), .I(I[1269]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1269_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst127(.CLK(CLK), .I(I[127]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst127_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1270(.CLK(CLK), .I(I[1270]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1270_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1271(.CLK(CLK), .I(I[1271]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1271_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1272(.CLK(CLK), .I(I[1272]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1272_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1273(.CLK(CLK), .I(I[1273]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1273_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1274(.CLK(CLK), .I(I[1274]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1274_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1275(.CLK(CLK), .I(I[1275]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1275_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1276(.CLK(CLK), .I(I[1276]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1276_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1277(.CLK(CLK), .I(I[1277]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1277_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1278(.CLK(CLK), .I(I[1278]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1278_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1279(.CLK(CLK), .I(I[1279]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1279_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst128(.CLK(CLK), .I(I[128]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst128_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1280(.CLK(CLK), .I(I[1280]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1280_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1281(.CLK(CLK), .I(I[1281]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1281_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1282(.CLK(CLK), .I(I[1282]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1282_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1283(.CLK(CLK), .I(I[1283]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1283_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1284(.CLK(CLK), .I(I[1284]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1284_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1285(.CLK(CLK), .I(I[1285]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1285_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1286(.CLK(CLK), .I(I[1286]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1286_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1287(.CLK(CLK), .I(I[1287]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1287_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1288(.CLK(CLK), .I(I[1288]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1288_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1289(.CLK(CLK), .I(I[1289]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1289_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst129(.CLK(CLK), .I(I[129]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst129_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1290(.CLK(CLK), .I(I[1290]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1290_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1291(.CLK(CLK), .I(I[1291]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1291_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1292(.CLK(CLK), .I(I[1292]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1292_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1293(.CLK(CLK), .I(I[1293]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1293_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1294(.CLK(CLK), .I(I[1294]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1294_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1295(.CLK(CLK), .I(I[1295]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1295_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1296(.CLK(CLK), .I(I[1296]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1296_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1297(.CLK(CLK), .I(I[1297]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1297_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1298(.CLK(CLK), .I(I[1298]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1298_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1299(.CLK(CLK), .I(I[1299]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1299_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13(.CLK(CLK), .I(I[13]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst130(.CLK(CLK), .I(I[130]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst130_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1300(.CLK(CLK), .I(I[1300]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1300_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1301(.CLK(CLK), .I(I[1301]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1301_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1302(.CLK(CLK), .I(I[1302]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1302_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1303(.CLK(CLK), .I(I[1303]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1303_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1304(.CLK(CLK), .I(I[1304]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1304_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1305(.CLK(CLK), .I(I[1305]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1305_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1306(.CLK(CLK), .I(I[1306]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1306_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1307(.CLK(CLK), .I(I[1307]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1307_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1308(.CLK(CLK), .I(I[1308]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1308_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1309(.CLK(CLK), .I(I[1309]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1309_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst131(.CLK(CLK), .I(I[131]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst131_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1310(.CLK(CLK), .I(I[1310]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1310_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1311(.CLK(CLK), .I(I[1311]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1311_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1312(.CLK(CLK), .I(I[1312]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1312_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1313(.CLK(CLK), .I(I[1313]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1313_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1314(.CLK(CLK), .I(I[1314]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1314_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1315(.CLK(CLK), .I(I[1315]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1315_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1316(.CLK(CLK), .I(I[1316]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1316_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1317(.CLK(CLK), .I(I[1317]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1317_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1318(.CLK(CLK), .I(I[1318]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1318_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1319(.CLK(CLK), .I(I[1319]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1319_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst132(.CLK(CLK), .I(I[132]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst132_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1320(.CLK(CLK), .I(I[1320]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1320_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1321(.CLK(CLK), .I(I[1321]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1321_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1322(.CLK(CLK), .I(I[1322]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1322_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1323(.CLK(CLK), .I(I[1323]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1323_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1324(.CLK(CLK), .I(I[1324]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1324_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1325(.CLK(CLK), .I(I[1325]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1325_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1326(.CLK(CLK), .I(I[1326]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1326_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1327(.CLK(CLK), .I(I[1327]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1327_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1328(.CLK(CLK), .I(I[1328]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1328_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1329(.CLK(CLK), .I(I[1329]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1329_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst133(.CLK(CLK), .I(I[133]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst133_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1330(.CLK(CLK), .I(I[1330]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1330_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1331(.CLK(CLK), .I(I[1331]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1331_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1332(.CLK(CLK), .I(I[1332]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1332_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1333(.CLK(CLK), .I(I[1333]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1333_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1334(.CLK(CLK), .I(I[1334]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1334_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1335(.CLK(CLK), .I(I[1335]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1335_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1336(.CLK(CLK), .I(I[1336]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1336_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1337(.CLK(CLK), .I(I[1337]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1337_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1338(.CLK(CLK), .I(I[1338]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1338_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1339(.CLK(CLK), .I(I[1339]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1339_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst134(.CLK(CLK), .I(I[134]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst134_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1340(.CLK(CLK), .I(I[1340]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1340_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1341(.CLK(CLK), .I(I[1341]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1341_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1342(.CLK(CLK), .I(I[1342]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1342_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1343(.CLK(CLK), .I(I[1343]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1343_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1344(.CLK(CLK), .I(I[1344]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1344_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1345(.CLK(CLK), .I(I[1345]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1345_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1346(.CLK(CLK), .I(I[1346]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1346_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1347(.CLK(CLK), .I(I[1347]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1347_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1348(.CLK(CLK), .I(I[1348]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1348_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1349(.CLK(CLK), .I(I[1349]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1349_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst135(.CLK(CLK), .I(I[135]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst135_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1350(.CLK(CLK), .I(I[1350]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1350_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1351(.CLK(CLK), .I(I[1351]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1351_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1352(.CLK(CLK), .I(I[1352]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1352_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1353(.CLK(CLK), .I(I[1353]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1353_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1354(.CLK(CLK), .I(I[1354]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1354_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1355(.CLK(CLK), .I(I[1355]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1355_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1356(.CLK(CLK), .I(I[1356]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1356_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1357(.CLK(CLK), .I(I[1357]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1357_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1358(.CLK(CLK), .I(I[1358]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1358_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1359(.CLK(CLK), .I(I[1359]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1359_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst136(.CLK(CLK), .I(I[136]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst136_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1360(.CLK(CLK), .I(I[1360]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1360_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1361(.CLK(CLK), .I(I[1361]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1361_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1362(.CLK(CLK), .I(I[1362]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1362_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1363(.CLK(CLK), .I(I[1363]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1363_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1364(.CLK(CLK), .I(I[1364]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1364_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1365(.CLK(CLK), .I(I[1365]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1365_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1366(.CLK(CLK), .I(I[1366]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1366_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1367(.CLK(CLK), .I(I[1367]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1367_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1368(.CLK(CLK), .I(I[1368]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1368_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1369(.CLK(CLK), .I(I[1369]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1369_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst137(.CLK(CLK), .I(I[137]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst137_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1370(.CLK(CLK), .I(I[1370]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1370_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1371(.CLK(CLK), .I(I[1371]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1371_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1372(.CLK(CLK), .I(I[1372]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1372_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1373(.CLK(CLK), .I(I[1373]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1373_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1374(.CLK(CLK), .I(I[1374]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1374_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1375(.CLK(CLK), .I(I[1375]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1375_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1376(.CLK(CLK), .I(I[1376]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1376_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1377(.CLK(CLK), .I(I[1377]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1377_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1378(.CLK(CLK), .I(I[1378]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1378_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1379(.CLK(CLK), .I(I[1379]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1379_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst138(.CLK(CLK), .I(I[138]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst138_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1380(.CLK(CLK), .I(I[1380]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1380_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1381(.CLK(CLK), .I(I[1381]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1381_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1382(.CLK(CLK), .I(I[1382]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1382_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1383(.CLK(CLK), .I(I[1383]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1383_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1384(.CLK(CLK), .I(I[1384]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1384_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1385(.CLK(CLK), .I(I[1385]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1385_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1386(.CLK(CLK), .I(I[1386]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1386_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1387(.CLK(CLK), .I(I[1387]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1387_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1388(.CLK(CLK), .I(I[1388]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1388_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1389(.CLK(CLK), .I(I[1389]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1389_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst139(.CLK(CLK), .I(I[139]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst139_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1390(.CLK(CLK), .I(I[1390]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1390_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1391(.CLK(CLK), .I(I[1391]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1391_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1392(.CLK(CLK), .I(I[1392]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1392_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1393(.CLK(CLK), .I(I[1393]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1393_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1394(.CLK(CLK), .I(I[1394]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1394_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1395(.CLK(CLK), .I(I[1395]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1395_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1396(.CLK(CLK), .I(I[1396]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1396_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1397(.CLK(CLK), .I(I[1397]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1397_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1398(.CLK(CLK), .I(I[1398]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1398_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1399(.CLK(CLK), .I(I[1399]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1399_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14(.CLK(CLK), .I(I[14]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst140(.CLK(CLK), .I(I[140]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst140_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1400(.CLK(CLK), .I(I[1400]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1400_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1401(.CLK(CLK), .I(I[1401]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1401_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1402(.CLK(CLK), .I(I[1402]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1402_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1403(.CLK(CLK), .I(I[1403]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1403_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1404(.CLK(CLK), .I(I[1404]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1404_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1405(.CLK(CLK), .I(I[1405]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1405_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1406(.CLK(CLK), .I(I[1406]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1406_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1407(.CLK(CLK), .I(I[1407]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1407_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1408(.CLK(CLK), .I(I[1408]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1408_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1409(.CLK(CLK), .I(I[1409]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1409_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst141(.CLK(CLK), .I(I[141]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst141_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1410(.CLK(CLK), .I(I[1410]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1410_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1411(.CLK(CLK), .I(I[1411]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1411_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1412(.CLK(CLK), .I(I[1412]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1412_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1413(.CLK(CLK), .I(I[1413]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1413_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1414(.CLK(CLK), .I(I[1414]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1414_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1415(.CLK(CLK), .I(I[1415]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1415_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1416(.CLK(CLK), .I(I[1416]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1416_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1417(.CLK(CLK), .I(I[1417]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1417_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1418(.CLK(CLK), .I(I[1418]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1418_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1419(.CLK(CLK), .I(I[1419]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1419_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst142(.CLK(CLK), .I(I[142]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst142_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1420(.CLK(CLK), .I(I[1420]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1420_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1421(.CLK(CLK), .I(I[1421]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1421_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1422(.CLK(CLK), .I(I[1422]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1422_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1423(.CLK(CLK), .I(I[1423]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1423_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1424(.CLK(CLK), .I(I[1424]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1424_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1425(.CLK(CLK), .I(I[1425]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1425_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1426(.CLK(CLK), .I(I[1426]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1426_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1427(.CLK(CLK), .I(I[1427]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1427_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1428(.CLK(CLK), .I(I[1428]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1428_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1429(.CLK(CLK), .I(I[1429]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1429_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst143(.CLK(CLK), .I(I[143]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst143_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1430(.CLK(CLK), .I(I[1430]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1430_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1431(.CLK(CLK), .I(I[1431]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1431_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1432(.CLK(CLK), .I(I[1432]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1432_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1433(.CLK(CLK), .I(I[1433]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1433_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1434(.CLK(CLK), .I(I[1434]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1434_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1435(.CLK(CLK), .I(I[1435]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1435_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1436(.CLK(CLK), .I(I[1436]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1436_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1437(.CLK(CLK), .I(I[1437]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1437_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1438(.CLK(CLK), .I(I[1438]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1438_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1439(.CLK(CLK), .I(I[1439]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1439_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst144(.CLK(CLK), .I(I[144]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst144_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1440(.CLK(CLK), .I(I[1440]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1440_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1441(.CLK(CLK), .I(I[1441]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1441_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1442(.CLK(CLK), .I(I[1442]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1442_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1443(.CLK(CLK), .I(I[1443]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1443_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1444(.CLK(CLK), .I(I[1444]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1444_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1445(.CLK(CLK), .I(I[1445]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1445_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1446(.CLK(CLK), .I(I[1446]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1446_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1447(.CLK(CLK), .I(I[1447]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1447_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1448(.CLK(CLK), .I(I[1448]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1448_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1449(.CLK(CLK), .I(I[1449]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1449_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst145(.CLK(CLK), .I(I[145]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst145_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1450(.CLK(CLK), .I(I[1450]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1450_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1451(.CLK(CLK), .I(I[1451]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1451_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1452(.CLK(CLK), .I(I[1452]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1452_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1453(.CLK(CLK), .I(I[1453]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1453_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1454(.CLK(CLK), .I(I[1454]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1454_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1455(.CLK(CLK), .I(I[1455]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1455_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1456(.CLK(CLK), .I(I[1456]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1456_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1457(.CLK(CLK), .I(I[1457]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1457_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1458(.CLK(CLK), .I(I[1458]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1458_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1459(.CLK(CLK), .I(I[1459]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1459_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst146(.CLK(CLK), .I(I[146]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst146_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1460(.CLK(CLK), .I(I[1460]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1460_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1461(.CLK(CLK), .I(I[1461]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1461_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1462(.CLK(CLK), .I(I[1462]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1462_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1463(.CLK(CLK), .I(I[1463]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1463_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1464(.CLK(CLK), .I(I[1464]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1464_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1465(.CLK(CLK), .I(I[1465]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1465_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1466(.CLK(CLK), .I(I[1466]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1466_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1467(.CLK(CLK), .I(I[1467]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1467_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1468(.CLK(CLK), .I(I[1468]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1468_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1469(.CLK(CLK), .I(I[1469]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1469_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst147(.CLK(CLK), .I(I[147]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst147_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1470(.CLK(CLK), .I(I[1470]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1470_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1471(.CLK(CLK), .I(I[1471]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1471_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1472(.CLK(CLK), .I(I[1472]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1472_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1473(.CLK(CLK), .I(I[1473]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1473_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1474(.CLK(CLK), .I(I[1474]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1474_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1475(.CLK(CLK), .I(I[1475]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1475_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1476(.CLK(CLK), .I(I[1476]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1476_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1477(.CLK(CLK), .I(I[1477]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1477_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1478(.CLK(CLK), .I(I[1478]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1478_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1479(.CLK(CLK), .I(I[1479]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1479_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst148(.CLK(CLK), .I(I[148]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst148_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1480(.CLK(CLK), .I(I[1480]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1480_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1481(.CLK(CLK), .I(I[1481]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1481_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1482(.CLK(CLK), .I(I[1482]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1482_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1483(.CLK(CLK), .I(I[1483]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1483_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1484(.CLK(CLK), .I(I[1484]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1484_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1485(.CLK(CLK), .I(I[1485]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1485_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1486(.CLK(CLK), .I(I[1486]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1486_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1487(.CLK(CLK), .I(I[1487]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1487_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1488(.CLK(CLK), .I(I[1488]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1488_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1489(.CLK(CLK), .I(I[1489]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1489_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst149(.CLK(CLK), .I(I[149]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst149_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1490(.CLK(CLK), .I(I[1490]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1490_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1491(.CLK(CLK), .I(I[1491]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1491_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1492(.CLK(CLK), .I(I[1492]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1492_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1493(.CLK(CLK), .I(I[1493]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1493_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1494(.CLK(CLK), .I(I[1494]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1494_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1495(.CLK(CLK), .I(I[1495]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1495_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1496(.CLK(CLK), .I(I[1496]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1496_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1497(.CLK(CLK), .I(I[1497]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1497_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1498(.CLK(CLK), .I(I[1498]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1498_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1499(.CLK(CLK), .I(I[1499]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1499_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15(.CLK(CLK), .I(I[15]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst150(.CLK(CLK), .I(I[150]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst150_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1500(.CLK(CLK), .I(I[1500]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1500_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1501(.CLK(CLK), .I(I[1501]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1501_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1502(.CLK(CLK), .I(I[1502]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1502_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1503(.CLK(CLK), .I(I[1503]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1503_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1504(.CLK(CLK), .I(I[1504]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1504_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1505(.CLK(CLK), .I(I[1505]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1505_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1506(.CLK(CLK), .I(I[1506]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1506_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1507(.CLK(CLK), .I(I[1507]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1507_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1508(.CLK(CLK), .I(I[1508]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1508_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1509(.CLK(CLK), .I(I[1509]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1509_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst151(.CLK(CLK), .I(I[151]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst151_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1510(.CLK(CLK), .I(I[1510]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1510_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1511(.CLK(CLK), .I(I[1511]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1511_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1512(.CLK(CLK), .I(I[1512]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1512_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1513(.CLK(CLK), .I(I[1513]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1513_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1514(.CLK(CLK), .I(I[1514]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1514_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1515(.CLK(CLK), .I(I[1515]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1515_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1516(.CLK(CLK), .I(I[1516]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1516_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1517(.CLK(CLK), .I(I[1517]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1517_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1518(.CLK(CLK), .I(I[1518]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1518_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1519(.CLK(CLK), .I(I[1519]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1519_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst152(.CLK(CLK), .I(I[152]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst152_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1520(.CLK(CLK), .I(I[1520]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1520_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1521(.CLK(CLK), .I(I[1521]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1521_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1522(.CLK(CLK), .I(I[1522]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1522_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1523(.CLK(CLK), .I(I[1523]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1523_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1524(.CLK(CLK), .I(I[1524]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1524_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1525(.CLK(CLK), .I(I[1525]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1525_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1526(.CLK(CLK), .I(I[1526]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1526_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1527(.CLK(CLK), .I(I[1527]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1527_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1528(.CLK(CLK), .I(I[1528]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1528_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1529(.CLK(CLK), .I(I[1529]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1529_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst153(.CLK(CLK), .I(I[153]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst153_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1530(.CLK(CLK), .I(I[1530]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1530_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1531(.CLK(CLK), .I(I[1531]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1531_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1532(.CLK(CLK), .I(I[1532]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1532_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1533(.CLK(CLK), .I(I[1533]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1533_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1534(.CLK(CLK), .I(I[1534]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1534_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1535(.CLK(CLK), .I(I[1535]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1535_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1536(.CLK(CLK), .I(I[1536]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1536_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1537(.CLK(CLK), .I(I[1537]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1537_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1538(.CLK(CLK), .I(I[1538]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1538_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1539(.CLK(CLK), .I(I[1539]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1539_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst154(.CLK(CLK), .I(I[154]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst154_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1540(.CLK(CLK), .I(I[1540]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1540_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1541(.CLK(CLK), .I(I[1541]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1541_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1542(.CLK(CLK), .I(I[1542]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1542_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1543(.CLK(CLK), .I(I[1543]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1543_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1544(.CLK(CLK), .I(I[1544]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1544_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1545(.CLK(CLK), .I(I[1545]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1545_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1546(.CLK(CLK), .I(I[1546]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1546_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1547(.CLK(CLK), .I(I[1547]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1547_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1548(.CLK(CLK), .I(I[1548]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1548_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1549(.CLK(CLK), .I(I[1549]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1549_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst155(.CLK(CLK), .I(I[155]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst155_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1550(.CLK(CLK), .I(I[1550]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1550_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1551(.CLK(CLK), .I(I[1551]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1551_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1552(.CLK(CLK), .I(I[1552]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1552_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1553(.CLK(CLK), .I(I[1553]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1553_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1554(.CLK(CLK), .I(I[1554]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1554_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1555(.CLK(CLK), .I(I[1555]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1555_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1556(.CLK(CLK), .I(I[1556]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1556_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1557(.CLK(CLK), .I(I[1557]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1557_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1558(.CLK(CLK), .I(I[1558]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1558_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1559(.CLK(CLK), .I(I[1559]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1559_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst156(.CLK(CLK), .I(I[156]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst156_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1560(.CLK(CLK), .I(I[1560]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1560_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1561(.CLK(CLK), .I(I[1561]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1561_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1562(.CLK(CLK), .I(I[1562]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1562_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1563(.CLK(CLK), .I(I[1563]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1563_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1564(.CLK(CLK), .I(I[1564]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1564_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1565(.CLK(CLK), .I(I[1565]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1565_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1566(.CLK(CLK), .I(I[1566]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1566_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1567(.CLK(CLK), .I(I[1567]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1567_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1568(.CLK(CLK), .I(I[1568]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1568_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1569(.CLK(CLK), .I(I[1569]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1569_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst157(.CLK(CLK), .I(I[157]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst157_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1570(.CLK(CLK), .I(I[1570]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1570_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1571(.CLK(CLK), .I(I[1571]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1571_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1572(.CLK(CLK), .I(I[1572]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1572_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1573(.CLK(CLK), .I(I[1573]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1573_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1574(.CLK(CLK), .I(I[1574]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1574_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1575(.CLK(CLK), .I(I[1575]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1575_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1576(.CLK(CLK), .I(I[1576]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1576_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1577(.CLK(CLK), .I(I[1577]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1577_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1578(.CLK(CLK), .I(I[1578]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1578_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1579(.CLK(CLK), .I(I[1579]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1579_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst158(.CLK(CLK), .I(I[158]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst158_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1580(.CLK(CLK), .I(I[1580]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1580_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1581(.CLK(CLK), .I(I[1581]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1581_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1582(.CLK(CLK), .I(I[1582]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1582_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1583(.CLK(CLK), .I(I[1583]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1583_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1584(.CLK(CLK), .I(I[1584]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1584_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1585(.CLK(CLK), .I(I[1585]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1585_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1586(.CLK(CLK), .I(I[1586]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1586_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1587(.CLK(CLK), .I(I[1587]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1587_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1588(.CLK(CLK), .I(I[1588]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1588_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1589(.CLK(CLK), .I(I[1589]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1589_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst159(.CLK(CLK), .I(I[159]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst159_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1590(.CLK(CLK), .I(I[1590]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1590_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1591(.CLK(CLK), .I(I[1591]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1591_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1592(.CLK(CLK), .I(I[1592]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1592_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1593(.CLK(CLK), .I(I[1593]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1593_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1594(.CLK(CLK), .I(I[1594]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1594_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1595(.CLK(CLK), .I(I[1595]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1595_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1596(.CLK(CLK), .I(I[1596]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1596_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1597(.CLK(CLK), .I(I[1597]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1597_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1598(.CLK(CLK), .I(I[1598]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1598_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1599(.CLK(CLK), .I(I[1599]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1599_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16(.CLK(CLK), .I(I[16]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst160(.CLK(CLK), .I(I[160]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst160_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst161(.CLK(CLK), .I(I[161]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst161_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst162(.CLK(CLK), .I(I[162]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst162_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst163(.CLK(CLK), .I(I[163]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst163_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst164(.CLK(CLK), .I(I[164]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst164_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst165(.CLK(CLK), .I(I[165]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst165_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst166(.CLK(CLK), .I(I[166]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst166_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst167(.CLK(CLK), .I(I[167]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst167_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst168(.CLK(CLK), .I(I[168]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst168_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst169(.CLK(CLK), .I(I[169]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst169_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17(.CLK(CLK), .I(I[17]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst170(.CLK(CLK), .I(I[170]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst170_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst171(.CLK(CLK), .I(I[171]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst171_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst172(.CLK(CLK), .I(I[172]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst172_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst173(.CLK(CLK), .I(I[173]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst173_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst174(.CLK(CLK), .I(I[174]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst174_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst175(.CLK(CLK), .I(I[175]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst175_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst176(.CLK(CLK), .I(I[176]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst176_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst177(.CLK(CLK), .I(I[177]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst177_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst178(.CLK(CLK), .I(I[178]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst178_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst179(.CLK(CLK), .I(I[179]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst179_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18(.CLK(CLK), .I(I[18]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst180(.CLK(CLK), .I(I[180]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst180_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst181(.CLK(CLK), .I(I[181]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst181_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst182(.CLK(CLK), .I(I[182]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst182_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst183(.CLK(CLK), .I(I[183]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst183_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst184(.CLK(CLK), .I(I[184]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst184_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst185(.CLK(CLK), .I(I[185]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst185_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst186(.CLK(CLK), .I(I[186]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst186_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst187(.CLK(CLK), .I(I[187]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst187_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst188(.CLK(CLK), .I(I[188]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst188_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst189(.CLK(CLK), .I(I[189]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst189_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19(.CLK(CLK), .I(I[19]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst190(.CLK(CLK), .I(I[190]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst190_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst191(.CLK(CLK), .I(I[191]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst191_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst192(.CLK(CLK), .I(I[192]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst192_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst193(.CLK(CLK), .I(I[193]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst193_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst194(.CLK(CLK), .I(I[194]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst194_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst195(.CLK(CLK), .I(I[195]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst195_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst196(.CLK(CLK), .I(I[196]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst196_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst197(.CLK(CLK), .I(I[197]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst197_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst198(.CLK(CLK), .I(I[198]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst198_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst199(.CLK(CLK), .I(I[199]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst199_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2(.CLK(CLK), .I(I[2]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20(.CLK(CLK), .I(I[20]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst200(.CLK(CLK), .I(I[200]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst200_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst201(.CLK(CLK), .I(I[201]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst201_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst202(.CLK(CLK), .I(I[202]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst202_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst203(.CLK(CLK), .I(I[203]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst203_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst204(.CLK(CLK), .I(I[204]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst204_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst205(.CLK(CLK), .I(I[205]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst205_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst206(.CLK(CLK), .I(I[206]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst206_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst207(.CLK(CLK), .I(I[207]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst207_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst208(.CLK(CLK), .I(I[208]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst208_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst209(.CLK(CLK), .I(I[209]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst209_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21(.CLK(CLK), .I(I[21]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst210(.CLK(CLK), .I(I[210]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst210_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst211(.CLK(CLK), .I(I[211]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst211_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst212(.CLK(CLK), .I(I[212]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst212_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst213(.CLK(CLK), .I(I[213]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst213_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst214(.CLK(CLK), .I(I[214]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst214_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst215(.CLK(CLK), .I(I[215]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst215_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst216(.CLK(CLK), .I(I[216]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst216_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst217(.CLK(CLK), .I(I[217]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst217_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst218(.CLK(CLK), .I(I[218]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst218_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst219(.CLK(CLK), .I(I[219]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst219_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22(.CLK(CLK), .I(I[22]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst220(.CLK(CLK), .I(I[220]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst220_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst221(.CLK(CLK), .I(I[221]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst221_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst222(.CLK(CLK), .I(I[222]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst222_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst223(.CLK(CLK), .I(I[223]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst223_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst224(.CLK(CLK), .I(I[224]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst224_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst225(.CLK(CLK), .I(I[225]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst225_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst226(.CLK(CLK), .I(I[226]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst226_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst227(.CLK(CLK), .I(I[227]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst227_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst228(.CLK(CLK), .I(I[228]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst228_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst229(.CLK(CLK), .I(I[229]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst229_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23(.CLK(CLK), .I(I[23]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst230(.CLK(CLK), .I(I[230]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst230_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst231(.CLK(CLK), .I(I[231]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst231_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst232(.CLK(CLK), .I(I[232]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst232_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst233(.CLK(CLK), .I(I[233]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst233_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst234(.CLK(CLK), .I(I[234]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst234_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst235(.CLK(CLK), .I(I[235]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst235_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst236(.CLK(CLK), .I(I[236]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst236_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst237(.CLK(CLK), .I(I[237]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst237_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst238(.CLK(CLK), .I(I[238]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst238_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst239(.CLK(CLK), .I(I[239]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst239_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24(.CLK(CLK), .I(I[24]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst240(.CLK(CLK), .I(I[240]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst240_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst241(.CLK(CLK), .I(I[241]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst241_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst242(.CLK(CLK), .I(I[242]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst242_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst243(.CLK(CLK), .I(I[243]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst243_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst244(.CLK(CLK), .I(I[244]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst244_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst245(.CLK(CLK), .I(I[245]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst245_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst246(.CLK(CLK), .I(I[246]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst246_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst247(.CLK(CLK), .I(I[247]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst247_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst248(.CLK(CLK), .I(I[248]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst248_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst249(.CLK(CLK), .I(I[249]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst249_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25(.CLK(CLK), .I(I[25]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst250(.CLK(CLK), .I(I[250]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst250_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst251(.CLK(CLK), .I(I[251]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst251_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst252(.CLK(CLK), .I(I[252]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst252_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst253(.CLK(CLK), .I(I[253]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst253_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst254(.CLK(CLK), .I(I[254]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst254_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst255(.CLK(CLK), .I(I[255]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst255_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst256(.CLK(CLK), .I(I[256]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst256_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst257(.CLK(CLK), .I(I[257]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst257_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst258(.CLK(CLK), .I(I[258]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst258_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst259(.CLK(CLK), .I(I[259]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst259_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26(.CLK(CLK), .I(I[26]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst260(.CLK(CLK), .I(I[260]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst260_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst261(.CLK(CLK), .I(I[261]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst261_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst262(.CLK(CLK), .I(I[262]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst262_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst263(.CLK(CLK), .I(I[263]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst263_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst264(.CLK(CLK), .I(I[264]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst264_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst265(.CLK(CLK), .I(I[265]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst265_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst266(.CLK(CLK), .I(I[266]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst266_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst267(.CLK(CLK), .I(I[267]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst267_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst268(.CLK(CLK), .I(I[268]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst268_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst269(.CLK(CLK), .I(I[269]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst269_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27(.CLK(CLK), .I(I[27]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst270(.CLK(CLK), .I(I[270]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst270_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst271(.CLK(CLK), .I(I[271]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst271_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst272(.CLK(CLK), .I(I[272]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst272_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst273(.CLK(CLK), .I(I[273]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst273_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst274(.CLK(CLK), .I(I[274]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst274_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst275(.CLK(CLK), .I(I[275]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst275_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst276(.CLK(CLK), .I(I[276]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst276_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst277(.CLK(CLK), .I(I[277]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst277_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst278(.CLK(CLK), .I(I[278]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst278_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst279(.CLK(CLK), .I(I[279]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst279_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28(.CLK(CLK), .I(I[28]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst280(.CLK(CLK), .I(I[280]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst280_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst281(.CLK(CLK), .I(I[281]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst281_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst282(.CLK(CLK), .I(I[282]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst282_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst283(.CLK(CLK), .I(I[283]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst283_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst284(.CLK(CLK), .I(I[284]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst284_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst285(.CLK(CLK), .I(I[285]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst285_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst286(.CLK(CLK), .I(I[286]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst286_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst287(.CLK(CLK), .I(I[287]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst287_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst288(.CLK(CLK), .I(I[288]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst288_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst289(.CLK(CLK), .I(I[289]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst289_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29(.CLK(CLK), .I(I[29]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst290(.CLK(CLK), .I(I[290]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst290_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst291(.CLK(CLK), .I(I[291]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst291_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst292(.CLK(CLK), .I(I[292]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst292_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst293(.CLK(CLK), .I(I[293]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst293_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst294(.CLK(CLK), .I(I[294]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst294_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst295(.CLK(CLK), .I(I[295]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst295_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst296(.CLK(CLK), .I(I[296]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst296_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst297(.CLK(CLK), .I(I[297]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst297_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst298(.CLK(CLK), .I(I[298]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst298_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst299(.CLK(CLK), .I(I[299]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst299_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3(.CLK(CLK), .I(I[3]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30(.CLK(CLK), .I(I[30]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst300(.CLK(CLK), .I(I[300]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst300_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst301(.CLK(CLK), .I(I[301]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst301_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst302(.CLK(CLK), .I(I[302]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst302_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst303(.CLK(CLK), .I(I[303]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst303_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst304(.CLK(CLK), .I(I[304]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst304_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst305(.CLK(CLK), .I(I[305]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst305_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst306(.CLK(CLK), .I(I[306]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst306_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst307(.CLK(CLK), .I(I[307]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst307_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst308(.CLK(CLK), .I(I[308]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst308_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst309(.CLK(CLK), .I(I[309]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst309_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31(.CLK(CLK), .I(I[31]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst310(.CLK(CLK), .I(I[310]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst310_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst311(.CLK(CLK), .I(I[311]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst311_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst312(.CLK(CLK), .I(I[312]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst312_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst313(.CLK(CLK), .I(I[313]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst313_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst314(.CLK(CLK), .I(I[314]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst314_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst315(.CLK(CLK), .I(I[315]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst315_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst316(.CLK(CLK), .I(I[316]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst316_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst317(.CLK(CLK), .I(I[317]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst317_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst318(.CLK(CLK), .I(I[318]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst318_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst319(.CLK(CLK), .I(I[319]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst319_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst32(.CLK(CLK), .I(I[32]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst32_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst320(.CLK(CLK), .I(I[320]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst320_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst321(.CLK(CLK), .I(I[321]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst321_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst322(.CLK(CLK), .I(I[322]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst322_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst323(.CLK(CLK), .I(I[323]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst323_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst324(.CLK(CLK), .I(I[324]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst324_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst325(.CLK(CLK), .I(I[325]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst325_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst326(.CLK(CLK), .I(I[326]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst326_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst327(.CLK(CLK), .I(I[327]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst327_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst328(.CLK(CLK), .I(I[328]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst328_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst329(.CLK(CLK), .I(I[329]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst329_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst33(.CLK(CLK), .I(I[33]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst33_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst330(.CLK(CLK), .I(I[330]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst330_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst331(.CLK(CLK), .I(I[331]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst331_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst332(.CLK(CLK), .I(I[332]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst332_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst333(.CLK(CLK), .I(I[333]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst333_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst334(.CLK(CLK), .I(I[334]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst334_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst335(.CLK(CLK), .I(I[335]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst335_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst336(.CLK(CLK), .I(I[336]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst336_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst337(.CLK(CLK), .I(I[337]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst337_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst338(.CLK(CLK), .I(I[338]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst338_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst339(.CLK(CLK), .I(I[339]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst339_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst34(.CLK(CLK), .I(I[34]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst34_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst340(.CLK(CLK), .I(I[340]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst340_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst341(.CLK(CLK), .I(I[341]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst341_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst342(.CLK(CLK), .I(I[342]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst342_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst343(.CLK(CLK), .I(I[343]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst343_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst344(.CLK(CLK), .I(I[344]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst344_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst345(.CLK(CLK), .I(I[345]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst345_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst346(.CLK(CLK), .I(I[346]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst346_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst347(.CLK(CLK), .I(I[347]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst347_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst348(.CLK(CLK), .I(I[348]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst348_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst349(.CLK(CLK), .I(I[349]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst349_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst35(.CLK(CLK), .I(I[35]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst35_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst350(.CLK(CLK), .I(I[350]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst350_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst351(.CLK(CLK), .I(I[351]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst351_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst352(.CLK(CLK), .I(I[352]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst352_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst353(.CLK(CLK), .I(I[353]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst353_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst354(.CLK(CLK), .I(I[354]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst354_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst355(.CLK(CLK), .I(I[355]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst355_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst356(.CLK(CLK), .I(I[356]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst356_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst357(.CLK(CLK), .I(I[357]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst357_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst358(.CLK(CLK), .I(I[358]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst358_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst359(.CLK(CLK), .I(I[359]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst359_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst36(.CLK(CLK), .I(I[36]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst36_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst360(.CLK(CLK), .I(I[360]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst360_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst361(.CLK(CLK), .I(I[361]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst361_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst362(.CLK(CLK), .I(I[362]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst362_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst363(.CLK(CLK), .I(I[363]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst363_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst364(.CLK(CLK), .I(I[364]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst364_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst365(.CLK(CLK), .I(I[365]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst365_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst366(.CLK(CLK), .I(I[366]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst366_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst367(.CLK(CLK), .I(I[367]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst367_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst368(.CLK(CLK), .I(I[368]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst368_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst369(.CLK(CLK), .I(I[369]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst369_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst37(.CLK(CLK), .I(I[37]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst37_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst370(.CLK(CLK), .I(I[370]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst370_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst371(.CLK(CLK), .I(I[371]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst371_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst372(.CLK(CLK), .I(I[372]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst372_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst373(.CLK(CLK), .I(I[373]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst373_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst374(.CLK(CLK), .I(I[374]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst374_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst375(.CLK(CLK), .I(I[375]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst375_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst376(.CLK(CLK), .I(I[376]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst376_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst377(.CLK(CLK), .I(I[377]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst377_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst378(.CLK(CLK), .I(I[378]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst378_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst379(.CLK(CLK), .I(I[379]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst379_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst38(.CLK(CLK), .I(I[38]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst38_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst380(.CLK(CLK), .I(I[380]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst380_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst381(.CLK(CLK), .I(I[381]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst381_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst382(.CLK(CLK), .I(I[382]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst382_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst383(.CLK(CLK), .I(I[383]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst383_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst384(.CLK(CLK), .I(I[384]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst384_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst385(.CLK(CLK), .I(I[385]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst385_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst386(.CLK(CLK), .I(I[386]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst386_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst387(.CLK(CLK), .I(I[387]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst387_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst388(.CLK(CLK), .I(I[388]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst388_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst389(.CLK(CLK), .I(I[389]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst389_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst39(.CLK(CLK), .I(I[39]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst39_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst390(.CLK(CLK), .I(I[390]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst390_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst391(.CLK(CLK), .I(I[391]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst391_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst392(.CLK(CLK), .I(I[392]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst392_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst393(.CLK(CLK), .I(I[393]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst393_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst394(.CLK(CLK), .I(I[394]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst394_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst395(.CLK(CLK), .I(I[395]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst395_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst396(.CLK(CLK), .I(I[396]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst396_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst397(.CLK(CLK), .I(I[397]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst397_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst398(.CLK(CLK), .I(I[398]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst398_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst399(.CLK(CLK), .I(I[399]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst399_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4(.CLK(CLK), .I(I[4]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst40(.CLK(CLK), .I(I[40]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst40_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst400(.CLK(CLK), .I(I[400]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst400_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst401(.CLK(CLK), .I(I[401]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst401_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst402(.CLK(CLK), .I(I[402]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst402_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst403(.CLK(CLK), .I(I[403]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst403_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst404(.CLK(CLK), .I(I[404]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst404_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst405(.CLK(CLK), .I(I[405]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst405_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst406(.CLK(CLK), .I(I[406]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst406_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst407(.CLK(CLK), .I(I[407]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst407_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst408(.CLK(CLK), .I(I[408]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst408_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst409(.CLK(CLK), .I(I[409]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst409_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst41(.CLK(CLK), .I(I[41]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst41_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst410(.CLK(CLK), .I(I[410]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst410_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst411(.CLK(CLK), .I(I[411]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst411_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst412(.CLK(CLK), .I(I[412]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst412_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst413(.CLK(CLK), .I(I[413]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst413_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst414(.CLK(CLK), .I(I[414]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst414_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst415(.CLK(CLK), .I(I[415]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst415_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst416(.CLK(CLK), .I(I[416]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst416_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst417(.CLK(CLK), .I(I[417]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst417_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst418(.CLK(CLK), .I(I[418]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst418_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst419(.CLK(CLK), .I(I[419]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst419_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst42(.CLK(CLK), .I(I[42]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst42_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst420(.CLK(CLK), .I(I[420]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst420_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst421(.CLK(CLK), .I(I[421]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst421_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst422(.CLK(CLK), .I(I[422]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst422_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst423(.CLK(CLK), .I(I[423]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst423_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst424(.CLK(CLK), .I(I[424]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst424_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst425(.CLK(CLK), .I(I[425]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst425_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst426(.CLK(CLK), .I(I[426]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst426_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst427(.CLK(CLK), .I(I[427]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst427_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst428(.CLK(CLK), .I(I[428]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst428_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst429(.CLK(CLK), .I(I[429]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst429_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst43(.CLK(CLK), .I(I[43]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst43_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst430(.CLK(CLK), .I(I[430]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst430_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst431(.CLK(CLK), .I(I[431]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst431_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst432(.CLK(CLK), .I(I[432]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst432_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst433(.CLK(CLK), .I(I[433]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst433_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst434(.CLK(CLK), .I(I[434]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst434_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst435(.CLK(CLK), .I(I[435]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst435_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst436(.CLK(CLK), .I(I[436]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst436_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst437(.CLK(CLK), .I(I[437]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst437_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst438(.CLK(CLK), .I(I[438]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst438_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst439(.CLK(CLK), .I(I[439]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst439_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst44(.CLK(CLK), .I(I[44]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst44_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst440(.CLK(CLK), .I(I[440]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst440_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst441(.CLK(CLK), .I(I[441]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst441_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst442(.CLK(CLK), .I(I[442]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst442_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst443(.CLK(CLK), .I(I[443]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst443_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst444(.CLK(CLK), .I(I[444]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst444_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst445(.CLK(CLK), .I(I[445]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst445_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst446(.CLK(CLK), .I(I[446]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst446_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst447(.CLK(CLK), .I(I[447]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst447_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst448(.CLK(CLK), .I(I[448]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst448_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst449(.CLK(CLK), .I(I[449]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst449_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst45(.CLK(CLK), .I(I[45]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst45_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst450(.CLK(CLK), .I(I[450]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst450_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst451(.CLK(CLK), .I(I[451]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst451_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst452(.CLK(CLK), .I(I[452]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst452_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst453(.CLK(CLK), .I(I[453]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst453_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst454(.CLK(CLK), .I(I[454]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst454_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst455(.CLK(CLK), .I(I[455]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst455_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst456(.CLK(CLK), .I(I[456]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst456_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst457(.CLK(CLK), .I(I[457]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst457_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst458(.CLK(CLK), .I(I[458]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst458_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst459(.CLK(CLK), .I(I[459]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst459_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst46(.CLK(CLK), .I(I[46]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst46_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst460(.CLK(CLK), .I(I[460]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst460_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst461(.CLK(CLK), .I(I[461]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst461_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst462(.CLK(CLK), .I(I[462]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst462_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst463(.CLK(CLK), .I(I[463]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst463_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst464(.CLK(CLK), .I(I[464]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst464_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst465(.CLK(CLK), .I(I[465]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst465_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst466(.CLK(CLK), .I(I[466]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst466_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst467(.CLK(CLK), .I(I[467]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst467_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst468(.CLK(CLK), .I(I[468]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst468_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst469(.CLK(CLK), .I(I[469]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst469_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst47(.CLK(CLK), .I(I[47]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst47_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst470(.CLK(CLK), .I(I[470]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst470_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst471(.CLK(CLK), .I(I[471]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst471_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst472(.CLK(CLK), .I(I[472]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst472_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst473(.CLK(CLK), .I(I[473]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst473_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst474(.CLK(CLK), .I(I[474]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst474_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst475(.CLK(CLK), .I(I[475]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst475_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst476(.CLK(CLK), .I(I[476]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst476_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst477(.CLK(CLK), .I(I[477]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst477_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst478(.CLK(CLK), .I(I[478]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst478_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst479(.CLK(CLK), .I(I[479]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst479_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst48(.CLK(CLK), .I(I[48]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst48_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst480(.CLK(CLK), .I(I[480]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst480_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst481(.CLK(CLK), .I(I[481]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst481_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst482(.CLK(CLK), .I(I[482]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst482_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst483(.CLK(CLK), .I(I[483]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst483_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst484(.CLK(CLK), .I(I[484]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst484_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst485(.CLK(CLK), .I(I[485]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst485_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst486(.CLK(CLK), .I(I[486]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst486_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst487(.CLK(CLK), .I(I[487]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst487_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst488(.CLK(CLK), .I(I[488]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst488_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst489(.CLK(CLK), .I(I[489]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst489_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst49(.CLK(CLK), .I(I[49]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst49_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst490(.CLK(CLK), .I(I[490]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst490_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst491(.CLK(CLK), .I(I[491]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst491_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst492(.CLK(CLK), .I(I[492]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst492_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst493(.CLK(CLK), .I(I[493]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst493_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst494(.CLK(CLK), .I(I[494]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst494_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst495(.CLK(CLK), .I(I[495]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst495_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst496(.CLK(CLK), .I(I[496]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst496_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst497(.CLK(CLK), .I(I[497]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst497_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst498(.CLK(CLK), .I(I[498]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst498_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst499(.CLK(CLK), .I(I[499]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst499_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5(.CLK(CLK), .I(I[5]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst50(.CLK(CLK), .I(I[50]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst50_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst500(.CLK(CLK), .I(I[500]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst500_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst501(.CLK(CLK), .I(I[501]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst501_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst502(.CLK(CLK), .I(I[502]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst502_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst503(.CLK(CLK), .I(I[503]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst503_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst504(.CLK(CLK), .I(I[504]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst504_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst505(.CLK(CLK), .I(I[505]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst505_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst506(.CLK(CLK), .I(I[506]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst506_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst507(.CLK(CLK), .I(I[507]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst507_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst508(.CLK(CLK), .I(I[508]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst508_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst509(.CLK(CLK), .I(I[509]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst509_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst51(.CLK(CLK), .I(I[51]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst51_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst510(.CLK(CLK), .I(I[510]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst510_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst511(.CLK(CLK), .I(I[511]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst511_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst512(.CLK(CLK), .I(I[512]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst512_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst513(.CLK(CLK), .I(I[513]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst513_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst514(.CLK(CLK), .I(I[514]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst514_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst515(.CLK(CLK), .I(I[515]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst515_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst516(.CLK(CLK), .I(I[516]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst516_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst517(.CLK(CLK), .I(I[517]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst517_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst518(.CLK(CLK), .I(I[518]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst518_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst519(.CLK(CLK), .I(I[519]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst519_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst52(.CLK(CLK), .I(I[52]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst52_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst520(.CLK(CLK), .I(I[520]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst520_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst521(.CLK(CLK), .I(I[521]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst521_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst522(.CLK(CLK), .I(I[522]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst522_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst523(.CLK(CLK), .I(I[523]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst523_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst524(.CLK(CLK), .I(I[524]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst524_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst525(.CLK(CLK), .I(I[525]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst525_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst526(.CLK(CLK), .I(I[526]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst526_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst527(.CLK(CLK), .I(I[527]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst527_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst528(.CLK(CLK), .I(I[528]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst528_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst529(.CLK(CLK), .I(I[529]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst529_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst53(.CLK(CLK), .I(I[53]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst53_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst530(.CLK(CLK), .I(I[530]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst530_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst531(.CLK(CLK), .I(I[531]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst531_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst532(.CLK(CLK), .I(I[532]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst532_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst533(.CLK(CLK), .I(I[533]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst533_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst534(.CLK(CLK), .I(I[534]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst534_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst535(.CLK(CLK), .I(I[535]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst535_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst536(.CLK(CLK), .I(I[536]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst536_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst537(.CLK(CLK), .I(I[537]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst537_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst538(.CLK(CLK), .I(I[538]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst538_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst539(.CLK(CLK), .I(I[539]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst539_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst54(.CLK(CLK), .I(I[54]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst54_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst540(.CLK(CLK), .I(I[540]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst540_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst541(.CLK(CLK), .I(I[541]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst541_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst542(.CLK(CLK), .I(I[542]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst542_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst543(.CLK(CLK), .I(I[543]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst543_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst544(.CLK(CLK), .I(I[544]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst544_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst545(.CLK(CLK), .I(I[545]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst545_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst546(.CLK(CLK), .I(I[546]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst546_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst547(.CLK(CLK), .I(I[547]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst547_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst548(.CLK(CLK), .I(I[548]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst548_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst549(.CLK(CLK), .I(I[549]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst549_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst55(.CLK(CLK), .I(I[55]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst55_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst550(.CLK(CLK), .I(I[550]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst550_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst551(.CLK(CLK), .I(I[551]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst551_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst552(.CLK(CLK), .I(I[552]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst552_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst553(.CLK(CLK), .I(I[553]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst553_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst554(.CLK(CLK), .I(I[554]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst554_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst555(.CLK(CLK), .I(I[555]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst555_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst556(.CLK(CLK), .I(I[556]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst556_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst557(.CLK(CLK), .I(I[557]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst557_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst558(.CLK(CLK), .I(I[558]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst558_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst559(.CLK(CLK), .I(I[559]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst559_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst56(.CLK(CLK), .I(I[56]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst56_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst560(.CLK(CLK), .I(I[560]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst560_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst561(.CLK(CLK), .I(I[561]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst561_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst562(.CLK(CLK), .I(I[562]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst562_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst563(.CLK(CLK), .I(I[563]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst563_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst564(.CLK(CLK), .I(I[564]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst564_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst565(.CLK(CLK), .I(I[565]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst565_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst566(.CLK(CLK), .I(I[566]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst566_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst567(.CLK(CLK), .I(I[567]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst567_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst568(.CLK(CLK), .I(I[568]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst568_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst569(.CLK(CLK), .I(I[569]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst569_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst57(.CLK(CLK), .I(I[57]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst57_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst570(.CLK(CLK), .I(I[570]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst570_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst571(.CLK(CLK), .I(I[571]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst571_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst572(.CLK(CLK), .I(I[572]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst572_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst573(.CLK(CLK), .I(I[573]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst573_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst574(.CLK(CLK), .I(I[574]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst574_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst575(.CLK(CLK), .I(I[575]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst575_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst576(.CLK(CLK), .I(I[576]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst576_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst577(.CLK(CLK), .I(I[577]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst577_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst578(.CLK(CLK), .I(I[578]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst578_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst579(.CLK(CLK), .I(I[579]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst579_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst58(.CLK(CLK), .I(I[58]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst58_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst580(.CLK(CLK), .I(I[580]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst580_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst581(.CLK(CLK), .I(I[581]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst581_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst582(.CLK(CLK), .I(I[582]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst582_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst583(.CLK(CLK), .I(I[583]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst583_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst584(.CLK(CLK), .I(I[584]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst584_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst585(.CLK(CLK), .I(I[585]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst585_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst586(.CLK(CLK), .I(I[586]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst586_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst587(.CLK(CLK), .I(I[587]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst587_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst588(.CLK(CLK), .I(I[588]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst588_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst589(.CLK(CLK), .I(I[589]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst589_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst59(.CLK(CLK), .I(I[59]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst59_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst590(.CLK(CLK), .I(I[590]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst590_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst591(.CLK(CLK), .I(I[591]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst591_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst592(.CLK(CLK), .I(I[592]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst592_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst593(.CLK(CLK), .I(I[593]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst593_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst594(.CLK(CLK), .I(I[594]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst594_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst595(.CLK(CLK), .I(I[595]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst595_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst596(.CLK(CLK), .I(I[596]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst596_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst597(.CLK(CLK), .I(I[597]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst597_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst598(.CLK(CLK), .I(I[598]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst598_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst599(.CLK(CLK), .I(I[599]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst599_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6(.CLK(CLK), .I(I[6]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst60(.CLK(CLK), .I(I[60]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst60_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst600(.CLK(CLK), .I(I[600]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst600_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst601(.CLK(CLK), .I(I[601]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst601_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst602(.CLK(CLK), .I(I[602]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst602_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst603(.CLK(CLK), .I(I[603]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst603_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst604(.CLK(CLK), .I(I[604]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst604_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst605(.CLK(CLK), .I(I[605]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst605_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst606(.CLK(CLK), .I(I[606]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst606_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst607(.CLK(CLK), .I(I[607]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst607_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst608(.CLK(CLK), .I(I[608]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst608_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst609(.CLK(CLK), .I(I[609]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst609_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst61(.CLK(CLK), .I(I[61]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst61_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst610(.CLK(CLK), .I(I[610]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst610_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst611(.CLK(CLK), .I(I[611]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst611_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst612(.CLK(CLK), .I(I[612]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst612_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst613(.CLK(CLK), .I(I[613]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst613_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst614(.CLK(CLK), .I(I[614]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst614_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst615(.CLK(CLK), .I(I[615]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst615_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst616(.CLK(CLK), .I(I[616]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst616_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst617(.CLK(CLK), .I(I[617]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst617_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst618(.CLK(CLK), .I(I[618]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst618_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst619(.CLK(CLK), .I(I[619]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst619_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst62(.CLK(CLK), .I(I[62]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst62_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst620(.CLK(CLK), .I(I[620]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst620_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst621(.CLK(CLK), .I(I[621]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst621_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst622(.CLK(CLK), .I(I[622]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst622_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst623(.CLK(CLK), .I(I[623]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst623_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst624(.CLK(CLK), .I(I[624]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst624_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst625(.CLK(CLK), .I(I[625]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst625_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst626(.CLK(CLK), .I(I[626]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst626_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst627(.CLK(CLK), .I(I[627]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst627_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst628(.CLK(CLK), .I(I[628]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst628_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst629(.CLK(CLK), .I(I[629]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst629_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst63(.CLK(CLK), .I(I[63]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst63_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst630(.CLK(CLK), .I(I[630]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst630_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst631(.CLK(CLK), .I(I[631]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst631_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst632(.CLK(CLK), .I(I[632]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst632_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst633(.CLK(CLK), .I(I[633]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst633_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst634(.CLK(CLK), .I(I[634]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst634_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst635(.CLK(CLK), .I(I[635]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst635_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst636(.CLK(CLK), .I(I[636]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst636_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst637(.CLK(CLK), .I(I[637]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst637_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst638(.CLK(CLK), .I(I[638]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst638_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst639(.CLK(CLK), .I(I[639]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst639_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst64(.CLK(CLK), .I(I[64]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst64_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst640(.CLK(CLK), .I(I[640]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst640_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst641(.CLK(CLK), .I(I[641]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst641_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst642(.CLK(CLK), .I(I[642]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst642_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst643(.CLK(CLK), .I(I[643]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst643_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst644(.CLK(CLK), .I(I[644]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst644_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst645(.CLK(CLK), .I(I[645]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst645_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst646(.CLK(CLK), .I(I[646]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst646_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst647(.CLK(CLK), .I(I[647]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst647_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst648(.CLK(CLK), .I(I[648]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst648_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst649(.CLK(CLK), .I(I[649]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst649_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst65(.CLK(CLK), .I(I[65]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst65_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst650(.CLK(CLK), .I(I[650]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst650_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst651(.CLK(CLK), .I(I[651]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst651_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst652(.CLK(CLK), .I(I[652]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst652_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst653(.CLK(CLK), .I(I[653]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst653_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst654(.CLK(CLK), .I(I[654]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst654_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst655(.CLK(CLK), .I(I[655]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst655_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst656(.CLK(CLK), .I(I[656]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst656_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst657(.CLK(CLK), .I(I[657]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst657_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst658(.CLK(CLK), .I(I[658]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst658_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst659(.CLK(CLK), .I(I[659]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst659_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst66(.CLK(CLK), .I(I[66]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst66_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst660(.CLK(CLK), .I(I[660]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst660_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst661(.CLK(CLK), .I(I[661]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst661_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst662(.CLK(CLK), .I(I[662]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst662_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst663(.CLK(CLK), .I(I[663]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst663_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst664(.CLK(CLK), .I(I[664]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst664_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst665(.CLK(CLK), .I(I[665]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst665_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst666(.CLK(CLK), .I(I[666]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst666_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst667(.CLK(CLK), .I(I[667]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst667_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst668(.CLK(CLK), .I(I[668]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst668_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst669(.CLK(CLK), .I(I[669]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst669_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst67(.CLK(CLK), .I(I[67]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst67_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst670(.CLK(CLK), .I(I[670]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst670_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst671(.CLK(CLK), .I(I[671]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst671_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst672(.CLK(CLK), .I(I[672]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst672_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst673(.CLK(CLK), .I(I[673]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst673_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst674(.CLK(CLK), .I(I[674]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst674_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst675(.CLK(CLK), .I(I[675]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst675_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst676(.CLK(CLK), .I(I[676]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst676_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst677(.CLK(CLK), .I(I[677]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst677_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst678(.CLK(CLK), .I(I[678]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst678_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst679(.CLK(CLK), .I(I[679]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst679_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst68(.CLK(CLK), .I(I[68]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst68_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst680(.CLK(CLK), .I(I[680]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst680_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst681(.CLK(CLK), .I(I[681]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst681_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst682(.CLK(CLK), .I(I[682]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst682_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst683(.CLK(CLK), .I(I[683]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst683_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst684(.CLK(CLK), .I(I[684]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst684_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst685(.CLK(CLK), .I(I[685]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst685_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst686(.CLK(CLK), .I(I[686]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst686_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst687(.CLK(CLK), .I(I[687]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst687_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst688(.CLK(CLK), .I(I[688]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst688_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst689(.CLK(CLK), .I(I[689]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst689_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst69(.CLK(CLK), .I(I[69]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst69_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst690(.CLK(CLK), .I(I[690]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst690_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst691(.CLK(CLK), .I(I[691]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst691_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst692(.CLK(CLK), .I(I[692]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst692_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst693(.CLK(CLK), .I(I[693]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst693_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst694(.CLK(CLK), .I(I[694]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst694_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst695(.CLK(CLK), .I(I[695]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst695_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst696(.CLK(CLK), .I(I[696]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst696_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst697(.CLK(CLK), .I(I[697]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst697_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst698(.CLK(CLK), .I(I[698]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst698_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst699(.CLK(CLK), .I(I[699]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst699_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7(.CLK(CLK), .I(I[7]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst70(.CLK(CLK), .I(I[70]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst70_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst700(.CLK(CLK), .I(I[700]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst700_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst701(.CLK(CLK), .I(I[701]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst701_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst702(.CLK(CLK), .I(I[702]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst702_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst703(.CLK(CLK), .I(I[703]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst703_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst704(.CLK(CLK), .I(I[704]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst704_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst705(.CLK(CLK), .I(I[705]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst705_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst706(.CLK(CLK), .I(I[706]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst706_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst707(.CLK(CLK), .I(I[707]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst707_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst708(.CLK(CLK), .I(I[708]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst708_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst709(.CLK(CLK), .I(I[709]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst709_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst71(.CLK(CLK), .I(I[71]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst71_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst710(.CLK(CLK), .I(I[710]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst710_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst711(.CLK(CLK), .I(I[711]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst711_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst712(.CLK(CLK), .I(I[712]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst712_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst713(.CLK(CLK), .I(I[713]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst713_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst714(.CLK(CLK), .I(I[714]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst714_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst715(.CLK(CLK), .I(I[715]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst715_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst716(.CLK(CLK), .I(I[716]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst716_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst717(.CLK(CLK), .I(I[717]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst717_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst718(.CLK(CLK), .I(I[718]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst718_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst719(.CLK(CLK), .I(I[719]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst719_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst72(.CLK(CLK), .I(I[72]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst72_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst720(.CLK(CLK), .I(I[720]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst720_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst721(.CLK(CLK), .I(I[721]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst721_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst722(.CLK(CLK), .I(I[722]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst722_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst723(.CLK(CLK), .I(I[723]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst723_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst724(.CLK(CLK), .I(I[724]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst724_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst725(.CLK(CLK), .I(I[725]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst725_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst726(.CLK(CLK), .I(I[726]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst726_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst727(.CLK(CLK), .I(I[727]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst727_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst728(.CLK(CLK), .I(I[728]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst728_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst729(.CLK(CLK), .I(I[729]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst729_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst73(.CLK(CLK), .I(I[73]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst73_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst730(.CLK(CLK), .I(I[730]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst730_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst731(.CLK(CLK), .I(I[731]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst731_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst732(.CLK(CLK), .I(I[732]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst732_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst733(.CLK(CLK), .I(I[733]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst733_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst734(.CLK(CLK), .I(I[734]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst734_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst735(.CLK(CLK), .I(I[735]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst735_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst736(.CLK(CLK), .I(I[736]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst736_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst737(.CLK(CLK), .I(I[737]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst737_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst738(.CLK(CLK), .I(I[738]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst738_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst739(.CLK(CLK), .I(I[739]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst739_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst74(.CLK(CLK), .I(I[74]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst74_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst740(.CLK(CLK), .I(I[740]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst740_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst741(.CLK(CLK), .I(I[741]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst741_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst742(.CLK(CLK), .I(I[742]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst742_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst743(.CLK(CLK), .I(I[743]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst743_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst744(.CLK(CLK), .I(I[744]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst744_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst745(.CLK(CLK), .I(I[745]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst745_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst746(.CLK(CLK), .I(I[746]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst746_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst747(.CLK(CLK), .I(I[747]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst747_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst748(.CLK(CLK), .I(I[748]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst748_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst749(.CLK(CLK), .I(I[749]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst749_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst75(.CLK(CLK), .I(I[75]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst75_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst750(.CLK(CLK), .I(I[750]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst750_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst751(.CLK(CLK), .I(I[751]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst751_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst752(.CLK(CLK), .I(I[752]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst752_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst753(.CLK(CLK), .I(I[753]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst753_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst754(.CLK(CLK), .I(I[754]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst754_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst755(.CLK(CLK), .I(I[755]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst755_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst756(.CLK(CLK), .I(I[756]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst756_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst757(.CLK(CLK), .I(I[757]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst757_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst758(.CLK(CLK), .I(I[758]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst758_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst759(.CLK(CLK), .I(I[759]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst759_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst76(.CLK(CLK), .I(I[76]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst76_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst760(.CLK(CLK), .I(I[760]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst760_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst761(.CLK(CLK), .I(I[761]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst761_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst762(.CLK(CLK), .I(I[762]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst762_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst763(.CLK(CLK), .I(I[763]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst763_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst764(.CLK(CLK), .I(I[764]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst764_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst765(.CLK(CLK), .I(I[765]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst765_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst766(.CLK(CLK), .I(I[766]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst766_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst767(.CLK(CLK), .I(I[767]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst767_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst768(.CLK(CLK), .I(I[768]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst768_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst769(.CLK(CLK), .I(I[769]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst769_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst77(.CLK(CLK), .I(I[77]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst77_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst770(.CLK(CLK), .I(I[770]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst770_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst771(.CLK(CLK), .I(I[771]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst771_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst772(.CLK(CLK), .I(I[772]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst772_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst773(.CLK(CLK), .I(I[773]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst773_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst774(.CLK(CLK), .I(I[774]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst774_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst775(.CLK(CLK), .I(I[775]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst775_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst776(.CLK(CLK), .I(I[776]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst776_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst777(.CLK(CLK), .I(I[777]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst777_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst778(.CLK(CLK), .I(I[778]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst778_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst779(.CLK(CLK), .I(I[779]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst779_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst78(.CLK(CLK), .I(I[78]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst78_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst780(.CLK(CLK), .I(I[780]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst780_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst781(.CLK(CLK), .I(I[781]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst781_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst782(.CLK(CLK), .I(I[782]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst782_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst783(.CLK(CLK), .I(I[783]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst783_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst784(.CLK(CLK), .I(I[784]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst784_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst785(.CLK(CLK), .I(I[785]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst785_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst786(.CLK(CLK), .I(I[786]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst786_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst787(.CLK(CLK), .I(I[787]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst787_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst788(.CLK(CLK), .I(I[788]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst788_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst789(.CLK(CLK), .I(I[789]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst789_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst79(.CLK(CLK), .I(I[79]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst79_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst790(.CLK(CLK), .I(I[790]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst790_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst791(.CLK(CLK), .I(I[791]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst791_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst792(.CLK(CLK), .I(I[792]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst792_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst793(.CLK(CLK), .I(I[793]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst793_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst794(.CLK(CLK), .I(I[794]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst794_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst795(.CLK(CLK), .I(I[795]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst795_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst796(.CLK(CLK), .I(I[796]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst796_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst797(.CLK(CLK), .I(I[797]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst797_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst798(.CLK(CLK), .I(I[798]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst798_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst799(.CLK(CLK), .I(I[799]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst799_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8(.CLK(CLK), .I(I[8]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst80(.CLK(CLK), .I(I[80]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst80_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst800(.CLK(CLK), .I(I[800]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst800_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst801(.CLK(CLK), .I(I[801]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst801_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst802(.CLK(CLK), .I(I[802]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst802_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst803(.CLK(CLK), .I(I[803]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst803_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst804(.CLK(CLK), .I(I[804]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst804_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst805(.CLK(CLK), .I(I[805]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst805_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst806(.CLK(CLK), .I(I[806]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst806_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst807(.CLK(CLK), .I(I[807]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst807_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst808(.CLK(CLK), .I(I[808]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst808_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst809(.CLK(CLK), .I(I[809]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst809_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst81(.CLK(CLK), .I(I[81]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst81_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst810(.CLK(CLK), .I(I[810]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst810_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst811(.CLK(CLK), .I(I[811]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst811_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst812(.CLK(CLK), .I(I[812]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst812_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst813(.CLK(CLK), .I(I[813]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst813_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst814(.CLK(CLK), .I(I[814]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst814_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst815(.CLK(CLK), .I(I[815]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst815_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst816(.CLK(CLK), .I(I[816]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst816_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst817(.CLK(CLK), .I(I[817]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst817_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst818(.CLK(CLK), .I(I[818]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst818_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst819(.CLK(CLK), .I(I[819]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst819_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst82(.CLK(CLK), .I(I[82]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst82_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst820(.CLK(CLK), .I(I[820]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst820_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst821(.CLK(CLK), .I(I[821]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst821_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst822(.CLK(CLK), .I(I[822]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst822_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst823(.CLK(CLK), .I(I[823]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst823_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst824(.CLK(CLK), .I(I[824]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst824_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst825(.CLK(CLK), .I(I[825]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst825_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst826(.CLK(CLK), .I(I[826]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst826_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst827(.CLK(CLK), .I(I[827]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst827_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst828(.CLK(CLK), .I(I[828]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst828_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst829(.CLK(CLK), .I(I[829]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst829_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst83(.CLK(CLK), .I(I[83]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst83_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst830(.CLK(CLK), .I(I[830]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst830_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst831(.CLK(CLK), .I(I[831]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst831_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst832(.CLK(CLK), .I(I[832]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst832_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst833(.CLK(CLK), .I(I[833]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst833_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst834(.CLK(CLK), .I(I[834]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst834_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst835(.CLK(CLK), .I(I[835]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst835_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst836(.CLK(CLK), .I(I[836]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst836_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst837(.CLK(CLK), .I(I[837]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst837_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst838(.CLK(CLK), .I(I[838]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst838_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst839(.CLK(CLK), .I(I[839]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst839_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst84(.CLK(CLK), .I(I[84]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst84_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst840(.CLK(CLK), .I(I[840]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst840_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst841(.CLK(CLK), .I(I[841]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst841_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst842(.CLK(CLK), .I(I[842]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst842_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst843(.CLK(CLK), .I(I[843]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst843_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst844(.CLK(CLK), .I(I[844]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst844_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst845(.CLK(CLK), .I(I[845]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst845_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst846(.CLK(CLK), .I(I[846]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst846_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst847(.CLK(CLK), .I(I[847]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst847_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst848(.CLK(CLK), .I(I[848]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst848_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst849(.CLK(CLK), .I(I[849]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst849_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst85(.CLK(CLK), .I(I[85]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst85_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst850(.CLK(CLK), .I(I[850]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst850_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst851(.CLK(CLK), .I(I[851]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst851_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst852(.CLK(CLK), .I(I[852]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst852_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst853(.CLK(CLK), .I(I[853]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst853_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst854(.CLK(CLK), .I(I[854]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst854_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst855(.CLK(CLK), .I(I[855]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst855_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst856(.CLK(CLK), .I(I[856]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst856_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst857(.CLK(CLK), .I(I[857]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst857_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst858(.CLK(CLK), .I(I[858]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst858_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst859(.CLK(CLK), .I(I[859]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst859_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst86(.CLK(CLK), .I(I[86]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst86_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst860(.CLK(CLK), .I(I[860]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst860_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst861(.CLK(CLK), .I(I[861]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst861_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst862(.CLK(CLK), .I(I[862]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst862_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst863(.CLK(CLK), .I(I[863]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst863_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst864(.CLK(CLK), .I(I[864]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst864_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst865(.CLK(CLK), .I(I[865]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst865_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst866(.CLK(CLK), .I(I[866]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst866_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst867(.CLK(CLK), .I(I[867]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst867_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst868(.CLK(CLK), .I(I[868]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst868_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst869(.CLK(CLK), .I(I[869]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst869_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst87(.CLK(CLK), .I(I[87]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst87_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst870(.CLK(CLK), .I(I[870]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst870_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst871(.CLK(CLK), .I(I[871]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst871_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst872(.CLK(CLK), .I(I[872]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst872_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst873(.CLK(CLK), .I(I[873]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst873_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst874(.CLK(CLK), .I(I[874]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst874_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst875(.CLK(CLK), .I(I[875]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst875_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst876(.CLK(CLK), .I(I[876]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst876_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst877(.CLK(CLK), .I(I[877]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst877_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst878(.CLK(CLK), .I(I[878]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst878_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst879(.CLK(CLK), .I(I[879]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst879_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst88(.CLK(CLK), .I(I[88]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst88_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst880(.CLK(CLK), .I(I[880]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst880_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst881(.CLK(CLK), .I(I[881]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst881_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst882(.CLK(CLK), .I(I[882]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst882_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst883(.CLK(CLK), .I(I[883]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst883_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst884(.CLK(CLK), .I(I[884]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst884_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst885(.CLK(CLK), .I(I[885]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst885_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst886(.CLK(CLK), .I(I[886]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst886_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst887(.CLK(CLK), .I(I[887]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst887_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst888(.CLK(CLK), .I(I[888]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst888_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst889(.CLK(CLK), .I(I[889]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst889_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst89(.CLK(CLK), .I(I[89]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst89_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst890(.CLK(CLK), .I(I[890]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst890_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst891(.CLK(CLK), .I(I[891]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst891_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst892(.CLK(CLK), .I(I[892]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst892_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst893(.CLK(CLK), .I(I[893]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst893_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst894(.CLK(CLK), .I(I[894]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst894_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst895(.CLK(CLK), .I(I[895]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst895_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst896(.CLK(CLK), .I(I[896]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst896_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst897(.CLK(CLK), .I(I[897]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst897_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst898(.CLK(CLK), .I(I[898]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst898_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst899(.CLK(CLK), .I(I[899]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst899_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9(.CLK(CLK), .I(I[9]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst90(.CLK(CLK), .I(I[90]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst90_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst900(.CLK(CLK), .I(I[900]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst900_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst901(.CLK(CLK), .I(I[901]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst901_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst902(.CLK(CLK), .I(I[902]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst902_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst903(.CLK(CLK), .I(I[903]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst903_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst904(.CLK(CLK), .I(I[904]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst904_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst905(.CLK(CLK), .I(I[905]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst905_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst906(.CLK(CLK), .I(I[906]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst906_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst907(.CLK(CLK), .I(I[907]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst907_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst908(.CLK(CLK), .I(I[908]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst908_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst909(.CLK(CLK), .I(I[909]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst909_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst91(.CLK(CLK), .I(I[91]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst91_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst910(.CLK(CLK), .I(I[910]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst910_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst911(.CLK(CLK), .I(I[911]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst911_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst912(.CLK(CLK), .I(I[912]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst912_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst913(.CLK(CLK), .I(I[913]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst913_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst914(.CLK(CLK), .I(I[914]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst914_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst915(.CLK(CLK), .I(I[915]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst915_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst916(.CLK(CLK), .I(I[916]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst916_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst917(.CLK(CLK), .I(I[917]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst917_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst918(.CLK(CLK), .I(I[918]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst918_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst919(.CLK(CLK), .I(I[919]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst919_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst92(.CLK(CLK), .I(I[92]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst92_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst920(.CLK(CLK), .I(I[920]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst920_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst921(.CLK(CLK), .I(I[921]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst921_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst922(.CLK(CLK), .I(I[922]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst922_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst923(.CLK(CLK), .I(I[923]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst923_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst924(.CLK(CLK), .I(I[924]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst924_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst925(.CLK(CLK), .I(I[925]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst925_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst926(.CLK(CLK), .I(I[926]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst926_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst927(.CLK(CLK), .I(I[927]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst927_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst928(.CLK(CLK), .I(I[928]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst928_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst929(.CLK(CLK), .I(I[929]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst929_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst93(.CLK(CLK), .I(I[93]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst93_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst930(.CLK(CLK), .I(I[930]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst930_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst931(.CLK(CLK), .I(I[931]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst931_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst932(.CLK(CLK), .I(I[932]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst932_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst933(.CLK(CLK), .I(I[933]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst933_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst934(.CLK(CLK), .I(I[934]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst934_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst935(.CLK(CLK), .I(I[935]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst935_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst936(.CLK(CLK), .I(I[936]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst936_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst937(.CLK(CLK), .I(I[937]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst937_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst938(.CLK(CLK), .I(I[938]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst938_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst939(.CLK(CLK), .I(I[939]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst939_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst94(.CLK(CLK), .I(I[94]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst94_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst940(.CLK(CLK), .I(I[940]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst940_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst941(.CLK(CLK), .I(I[941]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst941_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst942(.CLK(CLK), .I(I[942]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst942_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst943(.CLK(CLK), .I(I[943]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst943_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst944(.CLK(CLK), .I(I[944]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst944_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst945(.CLK(CLK), .I(I[945]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst945_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst946(.CLK(CLK), .I(I[946]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst946_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst947(.CLK(CLK), .I(I[947]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst947_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst948(.CLK(CLK), .I(I[948]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst948_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst949(.CLK(CLK), .I(I[949]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst949_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst95(.CLK(CLK), .I(I[95]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst95_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst950(.CLK(CLK), .I(I[950]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst950_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst951(.CLK(CLK), .I(I[951]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst951_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst952(.CLK(CLK), .I(I[952]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst952_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst953(.CLK(CLK), .I(I[953]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst953_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst954(.CLK(CLK), .I(I[954]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst954_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst955(.CLK(CLK), .I(I[955]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst955_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst956(.CLK(CLK), .I(I[956]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst956_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst957(.CLK(CLK), .I(I[957]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst957_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst958(.CLK(CLK), .I(I[958]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst958_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst959(.CLK(CLK), .I(I[959]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst959_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst96(.CLK(CLK), .I(I[96]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst96_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst960(.CLK(CLK), .I(I[960]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst960_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst961(.CLK(CLK), .I(I[961]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst961_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst962(.CLK(CLK), .I(I[962]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst962_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst963(.CLK(CLK), .I(I[963]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst963_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst964(.CLK(CLK), .I(I[964]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst964_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst965(.CLK(CLK), .I(I[965]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst965_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst966(.CLK(CLK), .I(I[966]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst966_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst967(.CLK(CLK), .I(I[967]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst967_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst968(.CLK(CLK), .I(I[968]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst968_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst969(.CLK(CLK), .I(I[969]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst969_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst97(.CLK(CLK), .I(I[97]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst97_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst970(.CLK(CLK), .I(I[970]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst970_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst971(.CLK(CLK), .I(I[971]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst971_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst972(.CLK(CLK), .I(I[972]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst972_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst973(.CLK(CLK), .I(I[973]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst973_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst974(.CLK(CLK), .I(I[974]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst974_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst975(.CLK(CLK), .I(I[975]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst975_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst976(.CLK(CLK), .I(I[976]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst976_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst977(.CLK(CLK), .I(I[977]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst977_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst978(.CLK(CLK), .I(I[978]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst978_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst979(.CLK(CLK), .I(I[979]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst979_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst98(.CLK(CLK), .I(I[98]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst98_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst980(.CLK(CLK), .I(I[980]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst980_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst981(.CLK(CLK), .I(I[981]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst981_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst982(.CLK(CLK), .I(I[982]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst982_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst983(.CLK(CLK), .I(I[983]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst983_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst984(.CLK(CLK), .I(I[984]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst984_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst985(.CLK(CLK), .I(I[985]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst985_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst986(.CLK(CLK), .I(I[986]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst986_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst987(.CLK(CLK), .I(I[987]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst987_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst988(.CLK(CLK), .I(I[988]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst988_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst989(.CLK(CLK), .I(I[989]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst989_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst99(.CLK(CLK), .I(I[99]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst99_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst990(.CLK(CLK), .I(I[990]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst990_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst991(.CLK(CLK), .I(I[991]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst991_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst992(.CLK(CLK), .I(I[992]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst992_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst993(.CLK(CLK), .I(I[993]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst993_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst994(.CLK(CLK), .I(I[994]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst994_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst995(.CLK(CLK), .I(I[995]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst995_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst996(.CLK(CLK), .I(I[996]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst996_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst997(.CLK(CLK), .I(I[997]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst997_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst998(.CLK(CLK), .I(I[998]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst998_O));
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst999(.CLK(CLK), .I(I[999]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst999_O));
assign O = {DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1599_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1598_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1597_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1596_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1595_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1594_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1593_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1592_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1591_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1590_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1589_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1588_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1587_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1586_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1585_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1584_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1583_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1582_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1581_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1580_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1579_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1578_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1577_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1576_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1575_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1574_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1573_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1572_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1571_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1570_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1569_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1568_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1567_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1566_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1565_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1564_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1563_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1562_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1561_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1560_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1559_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1558_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1557_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1556_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1555_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1554_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1553_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1552_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1551_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1550_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1549_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1548_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1547_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1546_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1545_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1544_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1543_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1542_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1541_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1540_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1539_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1538_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1537_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1536_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1535_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1534_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1533_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1532_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1531_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1530_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1529_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1528_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1527_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1526_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1525_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1524_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1523_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1522_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1521_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1520_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1519_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1518_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1517_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1516_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1515_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1514_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1513_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1512_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1511_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1510_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1509_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1508_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1507_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1506_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1505_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1504_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1503_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1502_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1501_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1500_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1499_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1498_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1497_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1496_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1495_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1494_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1493_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1492_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1491_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1490_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1489_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1488_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1487_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1486_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1485_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1484_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1483_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1482_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1481_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1480_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1479_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1478_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1477_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1476_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1475_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1474_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1473_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1472_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1471_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1470_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1469_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1468_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1467_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1466_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1465_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1464_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1463_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1462_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1461_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1460_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1459_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1458_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1457_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1456_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1455_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1454_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1453_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1452_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1451_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1450_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1449_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1448_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1447_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1446_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1445_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1444_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1443_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1442_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1441_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1440_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1439_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1438_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1437_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1436_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1435_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1434_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1433_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1432_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1431_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1430_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1429_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1428_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1427_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1426_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1425_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1424_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1423_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1422_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1421_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1420_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1419_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1418_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1417_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1416_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1415_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1414_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1413_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1412_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1411_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1410_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1409_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1408_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1407_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1406_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1405_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1404_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1403_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1402_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1401_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1400_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1399_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1398_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1397_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1396_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1395_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1394_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1393_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1392_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1391_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1390_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1389_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1388_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1387_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1386_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1385_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1384_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1383_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1382_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1381_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1380_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1379_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1378_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1377_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1376_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1375_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1374_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1373_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1372_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1371_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1370_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1369_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1368_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1367_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1366_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1365_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1364_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1363_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1362_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1361_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1360_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1359_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1358_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1357_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1356_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1355_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1354_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1353_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1352_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1351_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1350_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1349_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1348_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1347_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1346_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1345_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1344_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1343_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1342_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1341_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1340_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1339_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1338_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1337_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1336_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1335_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1334_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1333_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1332_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1331_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1330_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1329_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1328_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1327_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1326_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1325_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1324_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1323_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1322_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1321_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1320_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1319_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1318_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1317_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1316_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1315_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1314_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1313_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1312_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1311_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1310_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1309_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1308_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1307_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1306_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1305_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1304_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1303_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1302_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1301_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1300_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1299_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1298_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1297_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1296_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1295_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1294_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1293_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1292_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1291_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1290_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1289_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1288_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1287_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1286_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1285_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1284_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1283_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1282_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1281_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1280_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1279_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1278_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1277_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1276_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1275_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1274_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1273_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1272_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1271_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1270_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1269_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1268_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1267_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1266_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1265_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1264_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1263_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1262_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1261_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1260_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1259_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1258_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1257_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1256_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1255_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1254_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1253_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1252_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1251_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1250_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1249_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1248_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1247_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1246_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1245_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1244_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1243_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1242_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1241_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1240_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1239_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1238_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1237_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1236_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1235_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1234_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1233_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1232_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1231_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1230_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1229_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1228_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1227_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1226_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1225_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1224_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1223_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1222_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1221_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1220_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1219_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1218_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1217_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1216_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1215_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1214_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1213_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1212_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1211_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1210_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1209_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1208_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1207_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1206_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1205_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1204_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1203_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1202_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1201_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1200_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1199_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1198_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1197_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1196_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1195_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1194_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1193_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1192_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1191_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1190_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1189_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1188_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1187_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1186_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1185_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1184_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1183_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1182_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1181_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1180_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1179_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1178_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1177_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1176_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1175_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1174_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1173_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1172_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1171_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1170_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1169_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1168_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1167_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1166_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1165_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1164_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1163_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1162_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1161_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1160_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1159_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1158_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1157_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1156_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1155_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1154_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1153_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1152_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1151_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1150_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1149_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1148_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1147_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1146_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1145_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1144_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1143_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1142_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1141_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1140_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1139_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1138_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1137_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1136_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1135_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1134_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1133_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1132_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1131_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1130_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1129_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1128_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1127_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1126_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1125_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1124_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1123_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1122_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1121_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1120_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1119_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1118_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1117_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1116_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1115_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1114_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1113_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1112_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1111_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1110_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1109_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1108_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1107_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1106_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1105_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1104_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1103_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1102_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1101_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1100_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1099_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1098_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1097_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1096_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1095_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1094_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1093_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1092_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1091_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1090_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1089_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1088_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1087_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1086_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1085_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1084_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1083_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1082_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1081_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1080_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1079_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1078_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1077_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1076_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1075_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1074_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1073_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1072_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1071_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1070_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1069_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1068_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1067_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1066_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1065_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1064_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1063_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1062_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1061_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1060_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1059_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1058_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1057_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1056_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1055_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1054_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1053_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1052_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1051_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1050_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1049_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1048_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1047_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1046_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1045_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1044_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1043_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1042_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1041_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1040_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1039_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1038_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1037_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1036_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1035_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1034_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1033_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1032_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1031_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1030_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1029_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1028_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1027_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1026_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1025_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1024_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1023_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1022_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1021_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1020_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1019_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1018_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1017_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1016_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1015_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1014_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1013_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1012_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1011_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1010_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1009_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1008_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1007_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1006_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1005_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1004_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1003_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1002_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1001_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1000_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst999_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst998_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst997_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst996_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst995_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst994_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst993_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst992_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst991_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst990_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst989_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst988_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst987_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst986_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst985_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst984_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst983_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst982_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst981_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst980_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst979_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst978_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst977_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst976_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst975_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst974_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst973_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst972_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst971_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst970_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst969_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst968_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst967_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst966_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst965_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst964_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst963_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst962_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst961_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst960_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst959_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst958_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst957_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst956_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst955_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst954_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst953_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst952_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst951_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst950_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst949_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst948_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst947_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst946_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst945_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst944_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst943_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst942_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst941_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst940_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst939_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst938_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst937_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst936_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst935_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst934_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst933_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst932_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst931_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst930_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst929_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst928_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst927_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst926_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst925_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst924_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst923_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst922_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst921_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst920_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst919_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst918_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst917_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst916_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst915_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst914_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst913_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst912_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst911_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst910_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst909_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst908_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst907_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst906_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst905_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst904_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst903_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst902_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst901_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst900_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst899_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst898_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst897_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst896_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst895_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst894_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst893_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst892_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst891_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst890_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst889_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst888_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst887_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst886_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst885_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst884_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst883_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst882_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst881_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst880_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst879_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst878_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst877_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst876_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst875_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst874_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst873_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst872_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst871_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst870_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst869_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst868_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst867_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst866_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst865_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst864_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst863_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst862_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst861_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst860_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst859_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst858_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst857_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst856_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst855_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst854_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst853_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst852_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst851_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst850_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst849_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst848_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst847_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst846_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst845_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst844_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst843_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst842_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst841_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst840_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst839_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst838_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst837_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst836_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst835_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst834_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst833_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst832_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst831_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst830_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst829_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst828_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst827_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst826_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst825_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst824_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst823_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst822_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst821_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst820_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst819_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst818_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst817_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst816_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst815_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst814_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst813_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst812_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst811_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst810_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst809_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst808_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst807_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst806_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst805_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst804_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst803_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst802_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst801_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst800_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst799_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst798_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst797_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst796_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst795_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst794_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst793_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst792_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst791_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst790_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst789_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst788_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst787_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst786_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst785_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst784_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst783_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst782_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst781_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst780_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst779_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst778_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst777_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst776_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst775_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst774_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst773_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst772_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst771_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst770_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst769_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst768_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst767_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst766_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst765_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst764_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst763_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst762_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst761_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst760_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst759_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst758_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst757_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst756_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst755_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst754_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst753_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst752_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst751_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst750_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst749_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst748_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst747_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst746_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst745_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst744_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst743_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst742_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst741_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst740_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst739_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst738_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst737_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst736_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst735_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst734_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst733_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst732_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst731_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst730_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst729_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst728_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst727_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst726_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst725_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst724_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst723_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst722_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst721_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst720_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst719_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst718_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst717_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst716_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst715_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst714_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst713_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst712_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst711_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst710_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst709_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst708_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst707_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst706_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst705_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst704_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst703_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst702_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst701_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst700_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst699_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst698_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst697_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst696_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst695_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst694_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst693_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst692_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst691_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst690_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst689_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst688_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst687_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst686_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst685_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst684_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst683_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst682_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst681_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst680_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst679_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst678_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst677_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst676_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst675_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst674_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst673_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst672_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst671_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst670_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst669_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst668_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst667_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst666_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst665_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst664_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst663_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst662_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst661_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst660_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst659_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst658_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst657_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst656_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst655_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst654_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst653_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst652_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst651_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst650_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst649_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst648_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst647_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst646_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst645_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst644_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst643_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst642_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst641_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst640_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst639_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst638_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst637_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst636_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst635_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst634_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst633_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst632_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst631_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst630_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst629_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst628_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst627_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst626_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst625_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst624_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst623_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst622_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst621_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst620_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst619_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst618_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst617_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst616_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst615_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst614_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst613_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst612_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst611_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst610_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst609_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst608_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst607_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst606_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst605_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst604_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst603_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst602_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst601_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst600_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst599_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst598_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst597_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst596_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst595_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst594_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst593_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst592_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst591_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst590_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst589_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst588_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst587_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst586_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst585_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst584_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst583_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst582_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst581_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst580_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst579_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst578_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst577_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst576_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst575_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst574_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst573_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst572_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst571_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst570_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst569_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst568_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst567_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst566_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst565_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst564_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst563_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst562_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst561_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst560_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst559_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst558_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst557_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst556_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst555_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst554_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst553_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst552_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst551_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst550_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst549_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst548_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst547_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst546_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst545_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst544_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst543_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst542_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst541_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst540_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst539_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst538_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst537_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst536_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst535_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst534_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst533_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst532_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst531_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst530_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst529_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst528_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst527_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst526_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst525_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst524_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst523_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst522_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst521_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst520_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst519_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst518_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst517_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst516_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst515_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst514_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst513_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst512_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst511_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst510_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst509_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst508_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst507_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst506_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst505_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst504_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst503_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst502_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst501_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst500_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst499_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst498_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst497_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst496_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst495_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst494_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst493_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst492_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst491_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst490_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst489_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst488_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst487_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst486_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst485_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst484_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst483_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst482_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst481_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst480_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst479_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst478_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst477_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst476_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst475_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst474_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst473_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst472_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst471_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst470_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst469_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst468_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst467_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst466_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst465_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst464_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst463_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst462_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst461_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst460_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst459_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst458_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst457_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst456_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst455_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst454_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst453_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst452_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst451_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst450_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst449_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst448_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst447_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst446_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst445_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst444_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst443_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst442_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst441_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst440_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst439_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst438_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst437_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst436_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst435_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst434_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst433_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst432_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst431_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst430_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst429_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst428_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst427_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst426_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst425_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst424_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst423_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst422_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst421_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst420_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst419_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst418_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst417_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst416_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst415_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst414_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst413_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst412_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst411_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst410_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst409_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst408_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst407_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst406_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst405_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst404_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst403_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst402_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst401_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst400_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst399_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst398_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst397_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst396_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst395_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst394_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst393_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst392_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst391_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst390_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst389_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst388_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst387_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst386_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst385_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst384_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst383_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst382_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst381_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst380_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst379_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst378_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst377_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst376_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst375_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst374_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst373_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst372_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst371_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst370_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst369_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst368_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst367_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst366_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst365_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst364_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst363_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst362_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst361_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst360_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst359_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst358_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst357_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst356_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst355_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst354_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst353_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst352_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst351_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst350_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst349_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst348_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst347_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst346_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst345_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst344_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst343_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst342_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst341_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst340_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst339_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst338_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst337_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst336_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst335_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst334_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst333_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst332_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst331_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst330_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst329_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst328_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst327_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst326_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst325_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst324_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst323_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst322_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst321_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst320_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst319_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst318_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst317_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst316_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst315_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst314_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst313_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst312_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst311_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst310_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst309_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst308_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst307_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst306_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst305_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst304_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst303_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst302_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst301_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst300_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst299_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst298_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst297_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst296_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst295_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst294_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst293_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst292_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst291_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst290_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst289_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst288_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst287_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst286_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst285_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst284_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst283_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst282_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst281_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst280_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst279_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst278_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst277_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst276_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst275_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst274_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst273_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst272_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst271_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst270_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst269_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst268_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst267_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst266_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst265_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst264_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst263_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst262_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst261_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst260_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst259_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst258_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst257_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst256_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst255_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst254_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst253_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst252_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst251_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst250_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst249_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst248_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst247_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst246_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst245_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst244_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst243_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst242_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst241_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst240_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst239_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst238_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst237_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst236_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst235_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst234_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst233_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst232_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst231_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst230_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst229_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst228_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst227_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst226_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst225_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst224_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst223_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst222_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst221_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst220_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst219_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst218_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst217_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst216_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst215_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst214_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst213_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst212_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst211_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst210_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst209_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst208_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst207_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst206_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst205_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst204_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst203_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst202_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst201_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst200_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst199_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst198_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst197_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst196_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst195_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst194_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst193_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst192_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst191_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst190_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst189_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst188_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst187_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst186_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst185_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst184_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst183_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst182_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst181_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst180_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst179_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst178_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst177_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst176_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst175_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst174_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst173_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst172_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst171_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst170_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst169_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst168_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst167_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst166_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst165_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst164_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst163_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst162_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst161_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst160_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst159_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst158_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst157_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst156_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst155_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst154_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst153_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst152_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst151_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst150_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst149_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst148_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst147_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst146_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst145_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst144_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst143_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst142_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst141_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst140_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst139_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst138_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst137_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst136_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst135_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst134_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst133_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst132_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst131_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst130_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst129_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst128_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst127_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst126_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst125_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst124_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst123_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst122_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst121_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst120_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst119_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst118_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst117_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst116_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst115_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst114_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst113_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst112_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst111_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst110_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst109_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst108_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst107_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst106_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst105_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst104_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst103_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst102_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst101_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst100_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst99_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst98_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst97_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst96_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst95_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst94_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst93_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst92_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst91_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst90_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst89_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst88_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst87_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst86_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst85_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst84_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst83_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst82_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst81_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst80_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst79_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst78_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst77_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst76_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst75_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst74_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst73_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst72_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst71_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst70_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst69_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst68_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst67_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst66_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst65_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst64_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst63_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst62_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst61_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst60_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst59_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst58_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst57_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst56_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst55_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst54_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst53_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst52_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst51_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst50_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst49_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst48_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst47_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst46_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst45_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst44_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst43_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst42_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst41_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst40_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst39_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst38_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst37_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst36_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst35_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst34_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst33_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst32_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst31_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst30_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst29_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst28_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst27_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst26_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst25_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst24_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst23_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst22_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst21_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst20_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst19_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst18_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst17_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst16_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst15_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst14_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst13_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst12_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst11_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst10_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst9_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst8_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst7_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst6_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst5_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst4_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst3_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst2_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst1_O,DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O};
endmodule

module Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_100/*verilator public*/, input [7:0] I_101/*verilator public*/, input [7:0] I_102/*verilator public*/, input [7:0] I_103/*verilator public*/, input [7:0] I_104/*verilator public*/, input [7:0] I_105/*verilator public*/, input [7:0] I_106/*verilator public*/, input [7:0] I_107/*verilator public*/, input [7:0] I_108/*verilator public*/, input [7:0] I_109/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_110/*verilator public*/, input [7:0] I_111/*verilator public*/, input [7:0] I_112/*verilator public*/, input [7:0] I_113/*verilator public*/, input [7:0] I_114/*verilator public*/, input [7:0] I_115/*verilator public*/, input [7:0] I_116/*verilator public*/, input [7:0] I_117/*verilator public*/, input [7:0] I_118/*verilator public*/, input [7:0] I_119/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_120/*verilator public*/, input [7:0] I_121/*verilator public*/, input [7:0] I_122/*verilator public*/, input [7:0] I_123/*verilator public*/, input [7:0] I_124/*verilator public*/, input [7:0] I_125/*verilator public*/, input [7:0] I_126/*verilator public*/, input [7:0] I_127/*verilator public*/, input [7:0] I_128/*verilator public*/, input [7:0] I_129/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_130/*verilator public*/, input [7:0] I_131/*verilator public*/, input [7:0] I_132/*verilator public*/, input [7:0] I_133/*verilator public*/, input [7:0] I_134/*verilator public*/, input [7:0] I_135/*verilator public*/, input [7:0] I_136/*verilator public*/, input [7:0] I_137/*verilator public*/, input [7:0] I_138/*verilator public*/, input [7:0] I_139/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_140/*verilator public*/, input [7:0] I_141/*verilator public*/, input [7:0] I_142/*verilator public*/, input [7:0] I_143/*verilator public*/, input [7:0] I_144/*verilator public*/, input [7:0] I_145/*verilator public*/, input [7:0] I_146/*verilator public*/, input [7:0] I_147/*verilator public*/, input [7:0] I_148/*verilator public*/, input [7:0] I_149/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_150/*verilator public*/, input [7:0] I_151/*verilator public*/, input [7:0] I_152/*verilator public*/, input [7:0] I_153/*verilator public*/, input [7:0] I_154/*verilator public*/, input [7:0] I_155/*verilator public*/, input [7:0] I_156/*verilator public*/, input [7:0] I_157/*verilator public*/, input [7:0] I_158/*verilator public*/, input [7:0] I_159/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_160/*verilator public*/, input [7:0] I_161/*verilator public*/, input [7:0] I_162/*verilator public*/, input [7:0] I_163/*verilator public*/, input [7:0] I_164/*verilator public*/, input [7:0] I_165/*verilator public*/, input [7:0] I_166/*verilator public*/, input [7:0] I_167/*verilator public*/, input [7:0] I_168/*verilator public*/, input [7:0] I_169/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_170/*verilator public*/, input [7:0] I_171/*verilator public*/, input [7:0] I_172/*verilator public*/, input [7:0] I_173/*verilator public*/, input [7:0] I_174/*verilator public*/, input [7:0] I_175/*verilator public*/, input [7:0] I_176/*verilator public*/, input [7:0] I_177/*verilator public*/, input [7:0] I_178/*verilator public*/, input [7:0] I_179/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_180/*verilator public*/, input [7:0] I_181/*verilator public*/, input [7:0] I_182/*verilator public*/, input [7:0] I_183/*verilator public*/, input [7:0] I_184/*verilator public*/, input [7:0] I_185/*verilator public*/, input [7:0] I_186/*verilator public*/, input [7:0] I_187/*verilator public*/, input [7:0] I_188/*verilator public*/, input [7:0] I_189/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_190/*verilator public*/, input [7:0] I_191/*verilator public*/, input [7:0] I_192/*verilator public*/, input [7:0] I_193/*verilator public*/, input [7:0] I_194/*verilator public*/, input [7:0] I_195/*verilator public*/, input [7:0] I_196/*verilator public*/, input [7:0] I_197/*verilator public*/, input [7:0] I_198/*verilator public*/, input [7:0] I_199/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_40/*verilator public*/, input [7:0] I_41/*verilator public*/, input [7:0] I_42/*verilator public*/, input [7:0] I_43/*verilator public*/, input [7:0] I_44/*verilator public*/, input [7:0] I_45/*verilator public*/, input [7:0] I_46/*verilator public*/, input [7:0] I_47/*verilator public*/, input [7:0] I_48/*verilator public*/, input [7:0] I_49/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_50/*verilator public*/, input [7:0] I_51/*verilator public*/, input [7:0] I_52/*verilator public*/, input [7:0] I_53/*verilator public*/, input [7:0] I_54/*verilator public*/, input [7:0] I_55/*verilator public*/, input [7:0] I_56/*verilator public*/, input [7:0] I_57/*verilator public*/, input [7:0] I_58/*verilator public*/, input [7:0] I_59/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_60/*verilator public*/, input [7:0] I_61/*verilator public*/, input [7:0] I_62/*verilator public*/, input [7:0] I_63/*verilator public*/, input [7:0] I_64/*verilator public*/, input [7:0] I_65/*verilator public*/, input [7:0] I_66/*verilator public*/, input [7:0] I_67/*verilator public*/, input [7:0] I_68/*verilator public*/, input [7:0] I_69/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_70/*verilator public*/, input [7:0] I_71/*verilator public*/, input [7:0] I_72/*verilator public*/, input [7:0] I_73/*verilator public*/, input [7:0] I_74/*verilator public*/, input [7:0] I_75/*verilator public*/, input [7:0] I_76/*verilator public*/, input [7:0] I_77/*verilator public*/, input [7:0] I_78/*verilator public*/, input [7:0] I_79/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_80/*verilator public*/, input [7:0] I_81/*verilator public*/, input [7:0] I_82/*verilator public*/, input [7:0] I_83/*verilator public*/, input [7:0] I_84/*verilator public*/, input [7:0] I_85/*verilator public*/, input [7:0] I_86/*verilator public*/, input [7:0] I_87/*verilator public*/, input [7:0] I_88/*verilator public*/, input [7:0] I_89/*verilator public*/, input [7:0] I_9/*verilator public*/, input [7:0] I_90/*verilator public*/, input [7:0] I_91/*verilator public*/, input [7:0] I_92/*verilator public*/, input [7:0] I_93/*verilator public*/, input [7:0] I_94/*verilator public*/, input [7:0] I_95/*verilator public*/, input [7:0] I_96/*verilator public*/, input [7:0] I_97/*verilator public*/, input [7:0] I_98/*verilator public*/, input [7:0] I_99/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_100/*verilator public*/, output [7:0] O_101/*verilator public*/, output [7:0] O_102/*verilator public*/, output [7:0] O_103/*verilator public*/, output [7:0] O_104/*verilator public*/, output [7:0] O_105/*verilator public*/, output [7:0] O_106/*verilator public*/, output [7:0] O_107/*verilator public*/, output [7:0] O_108/*verilator public*/, output [7:0] O_109/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_110/*verilator public*/, output [7:0] O_111/*verilator public*/, output [7:0] O_112/*verilator public*/, output [7:0] O_113/*verilator public*/, output [7:0] O_114/*verilator public*/, output [7:0] O_115/*verilator public*/, output [7:0] O_116/*verilator public*/, output [7:0] O_117/*verilator public*/, output [7:0] O_118/*verilator public*/, output [7:0] O_119/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_120/*verilator public*/, output [7:0] O_121/*verilator public*/, output [7:0] O_122/*verilator public*/, output [7:0] O_123/*verilator public*/, output [7:0] O_124/*verilator public*/, output [7:0] O_125/*verilator public*/, output [7:0] O_126/*verilator public*/, output [7:0] O_127/*verilator public*/, output [7:0] O_128/*verilator public*/, output [7:0] O_129/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_130/*verilator public*/, output [7:0] O_131/*verilator public*/, output [7:0] O_132/*verilator public*/, output [7:0] O_133/*verilator public*/, output [7:0] O_134/*verilator public*/, output [7:0] O_135/*verilator public*/, output [7:0] O_136/*verilator public*/, output [7:0] O_137/*verilator public*/, output [7:0] O_138/*verilator public*/, output [7:0] O_139/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_140/*verilator public*/, output [7:0] O_141/*verilator public*/, output [7:0] O_142/*verilator public*/, output [7:0] O_143/*verilator public*/, output [7:0] O_144/*verilator public*/, output [7:0] O_145/*verilator public*/, output [7:0] O_146/*verilator public*/, output [7:0] O_147/*verilator public*/, output [7:0] O_148/*verilator public*/, output [7:0] O_149/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_150/*verilator public*/, output [7:0] O_151/*verilator public*/, output [7:0] O_152/*verilator public*/, output [7:0] O_153/*verilator public*/, output [7:0] O_154/*verilator public*/, output [7:0] O_155/*verilator public*/, output [7:0] O_156/*verilator public*/, output [7:0] O_157/*verilator public*/, output [7:0] O_158/*verilator public*/, output [7:0] O_159/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_160/*verilator public*/, output [7:0] O_161/*verilator public*/, output [7:0] O_162/*verilator public*/, output [7:0] O_163/*verilator public*/, output [7:0] O_164/*verilator public*/, output [7:0] O_165/*verilator public*/, output [7:0] O_166/*verilator public*/, output [7:0] O_167/*verilator public*/, output [7:0] O_168/*verilator public*/, output [7:0] O_169/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_170/*verilator public*/, output [7:0] O_171/*verilator public*/, output [7:0] O_172/*verilator public*/, output [7:0] O_173/*verilator public*/, output [7:0] O_174/*verilator public*/, output [7:0] O_175/*verilator public*/, output [7:0] O_176/*verilator public*/, output [7:0] O_177/*verilator public*/, output [7:0] O_178/*verilator public*/, output [7:0] O_179/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_180/*verilator public*/, output [7:0] O_181/*verilator public*/, output [7:0] O_182/*verilator public*/, output [7:0] O_183/*verilator public*/, output [7:0] O_184/*verilator public*/, output [7:0] O_185/*verilator public*/, output [7:0] O_186/*verilator public*/, output [7:0] O_187/*verilator public*/, output [7:0] O_188/*verilator public*/, output [7:0] O_189/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_190/*verilator public*/, output [7:0] O_191/*verilator public*/, output [7:0] O_192/*verilator public*/, output [7:0] O_193/*verilator public*/, output [7:0] O_194/*verilator public*/, output [7:0] O_195/*verilator public*/, output [7:0] O_196/*verilator public*/, output [7:0] O_197/*verilator public*/, output [7:0] O_198/*verilator public*/, output [7:0] O_199/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_40/*verilator public*/, output [7:0] O_41/*verilator public*/, output [7:0] O_42/*verilator public*/, output [7:0] O_43/*verilator public*/, output [7:0] O_44/*verilator public*/, output [7:0] O_45/*verilator public*/, output [7:0] O_46/*verilator public*/, output [7:0] O_47/*verilator public*/, output [7:0] O_48/*verilator public*/, output [7:0] O_49/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_50/*verilator public*/, output [7:0] O_51/*verilator public*/, output [7:0] O_52/*verilator public*/, output [7:0] O_53/*verilator public*/, output [7:0] O_54/*verilator public*/, output [7:0] O_55/*verilator public*/, output [7:0] O_56/*verilator public*/, output [7:0] O_57/*verilator public*/, output [7:0] O_58/*verilator public*/, output [7:0] O_59/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_60/*verilator public*/, output [7:0] O_61/*verilator public*/, output [7:0] O_62/*verilator public*/, output [7:0] O_63/*verilator public*/, output [7:0] O_64/*verilator public*/, output [7:0] O_65/*verilator public*/, output [7:0] O_66/*verilator public*/, output [7:0] O_67/*verilator public*/, output [7:0] O_68/*verilator public*/, output [7:0] O_69/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_70/*verilator public*/, output [7:0] O_71/*verilator public*/, output [7:0] O_72/*verilator public*/, output [7:0] O_73/*verilator public*/, output [7:0] O_74/*verilator public*/, output [7:0] O_75/*verilator public*/, output [7:0] O_76/*verilator public*/, output [7:0] O_77/*verilator public*/, output [7:0] O_78/*verilator public*/, output [7:0] O_79/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_80/*verilator public*/, output [7:0] O_81/*verilator public*/, output [7:0] O_82/*verilator public*/, output [7:0] O_83/*verilator public*/, output [7:0] O_84/*verilator public*/, output [7:0] O_85/*verilator public*/, output [7:0] O_86/*verilator public*/, output [7:0] O_87/*verilator public*/, output [7:0] O_88/*verilator public*/, output [7:0] O_89/*verilator public*/, output [7:0] O_9/*verilator public*/, output [7:0] O_90/*verilator public*/, output [7:0] O_91/*verilator public*/, output [7:0] O_92/*verilator public*/, output [7:0] O_93/*verilator public*/, output [7:0] O_94/*verilator public*/, output [7:0] O_95/*verilator public*/, output [7:0] O_96/*verilator public*/, output [7:0] O_97/*verilator public*/, output [7:0] O_98/*verilator public*/, output [7:0] O_99/*verilator public*/);
wire [1599:0] Register1600_inst0_O;
wire [1599:0] dehydrate_tArray_200_Array_8_Bit___inst0_out;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_0;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_1;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_10;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_100;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_101;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_102;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_103;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_104;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_105;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_106;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_107;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_108;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_109;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_11;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_110;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_111;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_112;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_113;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_114;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_115;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_116;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_117;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_118;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_119;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_12;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_120;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_121;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_122;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_123;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_124;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_125;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_126;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_127;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_128;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_129;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_13;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_130;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_131;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_132;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_133;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_134;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_135;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_136;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_137;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_138;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_139;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_14;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_140;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_141;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_142;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_143;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_144;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_145;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_146;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_147;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_148;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_149;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_15;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_150;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_151;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_152;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_153;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_154;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_155;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_156;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_157;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_158;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_159;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_16;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_160;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_161;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_162;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_163;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_164;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_165;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_166;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_167;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_168;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_169;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_17;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_170;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_171;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_172;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_173;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_174;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_175;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_176;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_177;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_178;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_179;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_18;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_180;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_181;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_182;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_183;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_184;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_185;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_186;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_187;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_188;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_189;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_19;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_190;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_191;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_192;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_193;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_194;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_195;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_196;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_197;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_198;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_199;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_2;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_20;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_21;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_22;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_23;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_24;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_25;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_26;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_27;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_28;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_29;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_3;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_30;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_31;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_32;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_33;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_34;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_35;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_36;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_37;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_38;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_39;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_4;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_40;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_41;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_42;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_43;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_44;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_45;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_46;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_47;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_48;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_49;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_5;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_50;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_51;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_52;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_53;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_54;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_55;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_56;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_57;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_58;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_59;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_6;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_60;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_61;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_62;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_63;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_64;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_65;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_66;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_67;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_68;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_69;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_7;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_70;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_71;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_72;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_73;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_74;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_75;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_76;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_77;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_78;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_79;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_8;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_80;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_81;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_82;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_83;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_84;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_85;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_86;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_87;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_88;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_89;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_9;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_90;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_91;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_92;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_93;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_94;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_95;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_96;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_97;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_98;
wire [7:0] hydrate_tArray_200_Array_8_Bit___inst0_out_99;
Register1600 Register1600_inst0(.CLK(CLK), .I(dehydrate_tArray_200_Array_8_Bit___inst0_out), .O(Register1600_inst0_O));
\aetherlinglib_dehydrate__hydratedTypeBit8200 dehydrate_tArray_200_Array_8_Bit___inst0(.in_0(I_0), .in_1(I_1), .in_10(I_10), .in_100(I_100), .in_101(I_101), .in_102(I_102), .in_103(I_103), .in_104(I_104), .in_105(I_105), .in_106(I_106), .in_107(I_107), .in_108(I_108), .in_109(I_109), .in_11(I_11), .in_110(I_110), .in_111(I_111), .in_112(I_112), .in_113(I_113), .in_114(I_114), .in_115(I_115), .in_116(I_116), .in_117(I_117), .in_118(I_118), .in_119(I_119), .in_12(I_12), .in_120(I_120), .in_121(I_121), .in_122(I_122), .in_123(I_123), .in_124(I_124), .in_125(I_125), .in_126(I_126), .in_127(I_127), .in_128(I_128), .in_129(I_129), .in_13(I_13), .in_130(I_130), .in_131(I_131), .in_132(I_132), .in_133(I_133), .in_134(I_134), .in_135(I_135), .in_136(I_136), .in_137(I_137), .in_138(I_138), .in_139(I_139), .in_14(I_14), .in_140(I_140), .in_141(I_141), .in_142(I_142), .in_143(I_143), .in_144(I_144), .in_145(I_145), .in_146(I_146), .in_147(I_147), .in_148(I_148), .in_149(I_149), .in_15(I_15), .in_150(I_150), .in_151(I_151), .in_152(I_152), .in_153(I_153), .in_154(I_154), .in_155(I_155), .in_156(I_156), .in_157(I_157), .in_158(I_158), .in_159(I_159), .in_16(I_16), .in_160(I_160), .in_161(I_161), .in_162(I_162), .in_163(I_163), .in_164(I_164), .in_165(I_165), .in_166(I_166), .in_167(I_167), .in_168(I_168), .in_169(I_169), .in_17(I_17), .in_170(I_170), .in_171(I_171), .in_172(I_172), .in_173(I_173), .in_174(I_174), .in_175(I_175), .in_176(I_176), .in_177(I_177), .in_178(I_178), .in_179(I_179), .in_18(I_18), .in_180(I_180), .in_181(I_181), .in_182(I_182), .in_183(I_183), .in_184(I_184), .in_185(I_185), .in_186(I_186), .in_187(I_187), .in_188(I_188), .in_189(I_189), .in_19(I_19), .in_190(I_190), .in_191(I_191), .in_192(I_192), .in_193(I_193), .in_194(I_194), .in_195(I_195), .in_196(I_196), .in_197(I_197), .in_198(I_198), .in_199(I_199), .in_2(I_2), .in_20(I_20), .in_21(I_21), .in_22(I_22), .in_23(I_23), .in_24(I_24), .in_25(I_25), .in_26(I_26), .in_27(I_27), .in_28(I_28), .in_29(I_29), .in_3(I_3), .in_30(I_30), .in_31(I_31), .in_32(I_32), .in_33(I_33), .in_34(I_34), .in_35(I_35), .in_36(I_36), .in_37(I_37), .in_38(I_38), .in_39(I_39), .in_4(I_4), .in_40(I_40), .in_41(I_41), .in_42(I_42), .in_43(I_43), .in_44(I_44), .in_45(I_45), .in_46(I_46), .in_47(I_47), .in_48(I_48), .in_49(I_49), .in_5(I_5), .in_50(I_50), .in_51(I_51), .in_52(I_52), .in_53(I_53), .in_54(I_54), .in_55(I_55), .in_56(I_56), .in_57(I_57), .in_58(I_58), .in_59(I_59), .in_6(I_6), .in_60(I_60), .in_61(I_61), .in_62(I_62), .in_63(I_63), .in_64(I_64), .in_65(I_65), .in_66(I_66), .in_67(I_67), .in_68(I_68), .in_69(I_69), .in_7(I_7), .in_70(I_70), .in_71(I_71), .in_72(I_72), .in_73(I_73), .in_74(I_74), .in_75(I_75), .in_76(I_76), .in_77(I_77), .in_78(I_78), .in_79(I_79), .in_8(I_8), .in_80(I_80), .in_81(I_81), .in_82(I_82), .in_83(I_83), .in_84(I_84), .in_85(I_85), .in_86(I_86), .in_87(I_87), .in_88(I_88), .in_89(I_89), .in_9(I_9), .in_90(I_90), .in_91(I_91), .in_92(I_92), .in_93(I_93), .in_94(I_94), .in_95(I_95), .in_96(I_96), .in_97(I_97), .in_98(I_98), .in_99(I_99), .out(dehydrate_tArray_200_Array_8_Bit___inst0_out));
\aetherlinglib_hydrate__hydratedTypeBit8200 hydrate_tArray_200_Array_8_Bit___inst0(.in(Register1600_inst0_O), .out_0(hydrate_tArray_200_Array_8_Bit___inst0_out_0), .out_1(hydrate_tArray_200_Array_8_Bit___inst0_out_1), .out_10(hydrate_tArray_200_Array_8_Bit___inst0_out_10), .out_100(hydrate_tArray_200_Array_8_Bit___inst0_out_100), .out_101(hydrate_tArray_200_Array_8_Bit___inst0_out_101), .out_102(hydrate_tArray_200_Array_8_Bit___inst0_out_102), .out_103(hydrate_tArray_200_Array_8_Bit___inst0_out_103), .out_104(hydrate_tArray_200_Array_8_Bit___inst0_out_104), .out_105(hydrate_tArray_200_Array_8_Bit___inst0_out_105), .out_106(hydrate_tArray_200_Array_8_Bit___inst0_out_106), .out_107(hydrate_tArray_200_Array_8_Bit___inst0_out_107), .out_108(hydrate_tArray_200_Array_8_Bit___inst0_out_108), .out_109(hydrate_tArray_200_Array_8_Bit___inst0_out_109), .out_11(hydrate_tArray_200_Array_8_Bit___inst0_out_11), .out_110(hydrate_tArray_200_Array_8_Bit___inst0_out_110), .out_111(hydrate_tArray_200_Array_8_Bit___inst0_out_111), .out_112(hydrate_tArray_200_Array_8_Bit___inst0_out_112), .out_113(hydrate_tArray_200_Array_8_Bit___inst0_out_113), .out_114(hydrate_tArray_200_Array_8_Bit___inst0_out_114), .out_115(hydrate_tArray_200_Array_8_Bit___inst0_out_115), .out_116(hydrate_tArray_200_Array_8_Bit___inst0_out_116), .out_117(hydrate_tArray_200_Array_8_Bit___inst0_out_117), .out_118(hydrate_tArray_200_Array_8_Bit___inst0_out_118), .out_119(hydrate_tArray_200_Array_8_Bit___inst0_out_119), .out_12(hydrate_tArray_200_Array_8_Bit___inst0_out_12), .out_120(hydrate_tArray_200_Array_8_Bit___inst0_out_120), .out_121(hydrate_tArray_200_Array_8_Bit___inst0_out_121), .out_122(hydrate_tArray_200_Array_8_Bit___inst0_out_122), .out_123(hydrate_tArray_200_Array_8_Bit___inst0_out_123), .out_124(hydrate_tArray_200_Array_8_Bit___inst0_out_124), .out_125(hydrate_tArray_200_Array_8_Bit___inst0_out_125), .out_126(hydrate_tArray_200_Array_8_Bit___inst0_out_126), .out_127(hydrate_tArray_200_Array_8_Bit___inst0_out_127), .out_128(hydrate_tArray_200_Array_8_Bit___inst0_out_128), .out_129(hydrate_tArray_200_Array_8_Bit___inst0_out_129), .out_13(hydrate_tArray_200_Array_8_Bit___inst0_out_13), .out_130(hydrate_tArray_200_Array_8_Bit___inst0_out_130), .out_131(hydrate_tArray_200_Array_8_Bit___inst0_out_131), .out_132(hydrate_tArray_200_Array_8_Bit___inst0_out_132), .out_133(hydrate_tArray_200_Array_8_Bit___inst0_out_133), .out_134(hydrate_tArray_200_Array_8_Bit___inst0_out_134), .out_135(hydrate_tArray_200_Array_8_Bit___inst0_out_135), .out_136(hydrate_tArray_200_Array_8_Bit___inst0_out_136), .out_137(hydrate_tArray_200_Array_8_Bit___inst0_out_137), .out_138(hydrate_tArray_200_Array_8_Bit___inst0_out_138), .out_139(hydrate_tArray_200_Array_8_Bit___inst0_out_139), .out_14(hydrate_tArray_200_Array_8_Bit___inst0_out_14), .out_140(hydrate_tArray_200_Array_8_Bit___inst0_out_140), .out_141(hydrate_tArray_200_Array_8_Bit___inst0_out_141), .out_142(hydrate_tArray_200_Array_8_Bit___inst0_out_142), .out_143(hydrate_tArray_200_Array_8_Bit___inst0_out_143), .out_144(hydrate_tArray_200_Array_8_Bit___inst0_out_144), .out_145(hydrate_tArray_200_Array_8_Bit___inst0_out_145), .out_146(hydrate_tArray_200_Array_8_Bit___inst0_out_146), .out_147(hydrate_tArray_200_Array_8_Bit___inst0_out_147), .out_148(hydrate_tArray_200_Array_8_Bit___inst0_out_148), .out_149(hydrate_tArray_200_Array_8_Bit___inst0_out_149), .out_15(hydrate_tArray_200_Array_8_Bit___inst0_out_15), .out_150(hydrate_tArray_200_Array_8_Bit___inst0_out_150), .out_151(hydrate_tArray_200_Array_8_Bit___inst0_out_151), .out_152(hydrate_tArray_200_Array_8_Bit___inst0_out_152), .out_153(hydrate_tArray_200_Array_8_Bit___inst0_out_153), .out_154(hydrate_tArray_200_Array_8_Bit___inst0_out_154), .out_155(hydrate_tArray_200_Array_8_Bit___inst0_out_155), .out_156(hydrate_tArray_200_Array_8_Bit___inst0_out_156), .out_157(hydrate_tArray_200_Array_8_Bit___inst0_out_157), .out_158(hydrate_tArray_200_Array_8_Bit___inst0_out_158), .out_159(hydrate_tArray_200_Array_8_Bit___inst0_out_159), .out_16(hydrate_tArray_200_Array_8_Bit___inst0_out_16), .out_160(hydrate_tArray_200_Array_8_Bit___inst0_out_160), .out_161(hydrate_tArray_200_Array_8_Bit___inst0_out_161), .out_162(hydrate_tArray_200_Array_8_Bit___inst0_out_162), .out_163(hydrate_tArray_200_Array_8_Bit___inst0_out_163), .out_164(hydrate_tArray_200_Array_8_Bit___inst0_out_164), .out_165(hydrate_tArray_200_Array_8_Bit___inst0_out_165), .out_166(hydrate_tArray_200_Array_8_Bit___inst0_out_166), .out_167(hydrate_tArray_200_Array_8_Bit___inst0_out_167), .out_168(hydrate_tArray_200_Array_8_Bit___inst0_out_168), .out_169(hydrate_tArray_200_Array_8_Bit___inst0_out_169), .out_17(hydrate_tArray_200_Array_8_Bit___inst0_out_17), .out_170(hydrate_tArray_200_Array_8_Bit___inst0_out_170), .out_171(hydrate_tArray_200_Array_8_Bit___inst0_out_171), .out_172(hydrate_tArray_200_Array_8_Bit___inst0_out_172), .out_173(hydrate_tArray_200_Array_8_Bit___inst0_out_173), .out_174(hydrate_tArray_200_Array_8_Bit___inst0_out_174), .out_175(hydrate_tArray_200_Array_8_Bit___inst0_out_175), .out_176(hydrate_tArray_200_Array_8_Bit___inst0_out_176), .out_177(hydrate_tArray_200_Array_8_Bit___inst0_out_177), .out_178(hydrate_tArray_200_Array_8_Bit___inst0_out_178), .out_179(hydrate_tArray_200_Array_8_Bit___inst0_out_179), .out_18(hydrate_tArray_200_Array_8_Bit___inst0_out_18), .out_180(hydrate_tArray_200_Array_8_Bit___inst0_out_180), .out_181(hydrate_tArray_200_Array_8_Bit___inst0_out_181), .out_182(hydrate_tArray_200_Array_8_Bit___inst0_out_182), .out_183(hydrate_tArray_200_Array_8_Bit___inst0_out_183), .out_184(hydrate_tArray_200_Array_8_Bit___inst0_out_184), .out_185(hydrate_tArray_200_Array_8_Bit___inst0_out_185), .out_186(hydrate_tArray_200_Array_8_Bit___inst0_out_186), .out_187(hydrate_tArray_200_Array_8_Bit___inst0_out_187), .out_188(hydrate_tArray_200_Array_8_Bit___inst0_out_188), .out_189(hydrate_tArray_200_Array_8_Bit___inst0_out_189), .out_19(hydrate_tArray_200_Array_8_Bit___inst0_out_19), .out_190(hydrate_tArray_200_Array_8_Bit___inst0_out_190), .out_191(hydrate_tArray_200_Array_8_Bit___inst0_out_191), .out_192(hydrate_tArray_200_Array_8_Bit___inst0_out_192), .out_193(hydrate_tArray_200_Array_8_Bit___inst0_out_193), .out_194(hydrate_tArray_200_Array_8_Bit___inst0_out_194), .out_195(hydrate_tArray_200_Array_8_Bit___inst0_out_195), .out_196(hydrate_tArray_200_Array_8_Bit___inst0_out_196), .out_197(hydrate_tArray_200_Array_8_Bit___inst0_out_197), .out_198(hydrate_tArray_200_Array_8_Bit___inst0_out_198), .out_199(hydrate_tArray_200_Array_8_Bit___inst0_out_199), .out_2(hydrate_tArray_200_Array_8_Bit___inst0_out_2), .out_20(hydrate_tArray_200_Array_8_Bit___inst0_out_20), .out_21(hydrate_tArray_200_Array_8_Bit___inst0_out_21), .out_22(hydrate_tArray_200_Array_8_Bit___inst0_out_22), .out_23(hydrate_tArray_200_Array_8_Bit___inst0_out_23), .out_24(hydrate_tArray_200_Array_8_Bit___inst0_out_24), .out_25(hydrate_tArray_200_Array_8_Bit___inst0_out_25), .out_26(hydrate_tArray_200_Array_8_Bit___inst0_out_26), .out_27(hydrate_tArray_200_Array_8_Bit___inst0_out_27), .out_28(hydrate_tArray_200_Array_8_Bit___inst0_out_28), .out_29(hydrate_tArray_200_Array_8_Bit___inst0_out_29), .out_3(hydrate_tArray_200_Array_8_Bit___inst0_out_3), .out_30(hydrate_tArray_200_Array_8_Bit___inst0_out_30), .out_31(hydrate_tArray_200_Array_8_Bit___inst0_out_31), .out_32(hydrate_tArray_200_Array_8_Bit___inst0_out_32), .out_33(hydrate_tArray_200_Array_8_Bit___inst0_out_33), .out_34(hydrate_tArray_200_Array_8_Bit___inst0_out_34), .out_35(hydrate_tArray_200_Array_8_Bit___inst0_out_35), .out_36(hydrate_tArray_200_Array_8_Bit___inst0_out_36), .out_37(hydrate_tArray_200_Array_8_Bit___inst0_out_37), .out_38(hydrate_tArray_200_Array_8_Bit___inst0_out_38), .out_39(hydrate_tArray_200_Array_8_Bit___inst0_out_39), .out_4(hydrate_tArray_200_Array_8_Bit___inst0_out_4), .out_40(hydrate_tArray_200_Array_8_Bit___inst0_out_40), .out_41(hydrate_tArray_200_Array_8_Bit___inst0_out_41), .out_42(hydrate_tArray_200_Array_8_Bit___inst0_out_42), .out_43(hydrate_tArray_200_Array_8_Bit___inst0_out_43), .out_44(hydrate_tArray_200_Array_8_Bit___inst0_out_44), .out_45(hydrate_tArray_200_Array_8_Bit___inst0_out_45), .out_46(hydrate_tArray_200_Array_8_Bit___inst0_out_46), .out_47(hydrate_tArray_200_Array_8_Bit___inst0_out_47), .out_48(hydrate_tArray_200_Array_8_Bit___inst0_out_48), .out_49(hydrate_tArray_200_Array_8_Bit___inst0_out_49), .out_5(hydrate_tArray_200_Array_8_Bit___inst0_out_5), .out_50(hydrate_tArray_200_Array_8_Bit___inst0_out_50), .out_51(hydrate_tArray_200_Array_8_Bit___inst0_out_51), .out_52(hydrate_tArray_200_Array_8_Bit___inst0_out_52), .out_53(hydrate_tArray_200_Array_8_Bit___inst0_out_53), .out_54(hydrate_tArray_200_Array_8_Bit___inst0_out_54), .out_55(hydrate_tArray_200_Array_8_Bit___inst0_out_55), .out_56(hydrate_tArray_200_Array_8_Bit___inst0_out_56), .out_57(hydrate_tArray_200_Array_8_Bit___inst0_out_57), .out_58(hydrate_tArray_200_Array_8_Bit___inst0_out_58), .out_59(hydrate_tArray_200_Array_8_Bit___inst0_out_59), .out_6(hydrate_tArray_200_Array_8_Bit___inst0_out_6), .out_60(hydrate_tArray_200_Array_8_Bit___inst0_out_60), .out_61(hydrate_tArray_200_Array_8_Bit___inst0_out_61), .out_62(hydrate_tArray_200_Array_8_Bit___inst0_out_62), .out_63(hydrate_tArray_200_Array_8_Bit___inst0_out_63), .out_64(hydrate_tArray_200_Array_8_Bit___inst0_out_64), .out_65(hydrate_tArray_200_Array_8_Bit___inst0_out_65), .out_66(hydrate_tArray_200_Array_8_Bit___inst0_out_66), .out_67(hydrate_tArray_200_Array_8_Bit___inst0_out_67), .out_68(hydrate_tArray_200_Array_8_Bit___inst0_out_68), .out_69(hydrate_tArray_200_Array_8_Bit___inst0_out_69), .out_7(hydrate_tArray_200_Array_8_Bit___inst0_out_7), .out_70(hydrate_tArray_200_Array_8_Bit___inst0_out_70), .out_71(hydrate_tArray_200_Array_8_Bit___inst0_out_71), .out_72(hydrate_tArray_200_Array_8_Bit___inst0_out_72), .out_73(hydrate_tArray_200_Array_8_Bit___inst0_out_73), .out_74(hydrate_tArray_200_Array_8_Bit___inst0_out_74), .out_75(hydrate_tArray_200_Array_8_Bit___inst0_out_75), .out_76(hydrate_tArray_200_Array_8_Bit___inst0_out_76), .out_77(hydrate_tArray_200_Array_8_Bit___inst0_out_77), .out_78(hydrate_tArray_200_Array_8_Bit___inst0_out_78), .out_79(hydrate_tArray_200_Array_8_Bit___inst0_out_79), .out_8(hydrate_tArray_200_Array_8_Bit___inst0_out_8), .out_80(hydrate_tArray_200_Array_8_Bit___inst0_out_80), .out_81(hydrate_tArray_200_Array_8_Bit___inst0_out_81), .out_82(hydrate_tArray_200_Array_8_Bit___inst0_out_82), .out_83(hydrate_tArray_200_Array_8_Bit___inst0_out_83), .out_84(hydrate_tArray_200_Array_8_Bit___inst0_out_84), .out_85(hydrate_tArray_200_Array_8_Bit___inst0_out_85), .out_86(hydrate_tArray_200_Array_8_Bit___inst0_out_86), .out_87(hydrate_tArray_200_Array_8_Bit___inst0_out_87), .out_88(hydrate_tArray_200_Array_8_Bit___inst0_out_88), .out_89(hydrate_tArray_200_Array_8_Bit___inst0_out_89), .out_9(hydrate_tArray_200_Array_8_Bit___inst0_out_9), .out_90(hydrate_tArray_200_Array_8_Bit___inst0_out_90), .out_91(hydrate_tArray_200_Array_8_Bit___inst0_out_91), .out_92(hydrate_tArray_200_Array_8_Bit___inst0_out_92), .out_93(hydrate_tArray_200_Array_8_Bit___inst0_out_93), .out_94(hydrate_tArray_200_Array_8_Bit___inst0_out_94), .out_95(hydrate_tArray_200_Array_8_Bit___inst0_out_95), .out_96(hydrate_tArray_200_Array_8_Bit___inst0_out_96), .out_97(hydrate_tArray_200_Array_8_Bit___inst0_out_97), .out_98(hydrate_tArray_200_Array_8_Bit___inst0_out_98), .out_99(hydrate_tArray_200_Array_8_Bit___inst0_out_99));
assign O_0 = hydrate_tArray_200_Array_8_Bit___inst0_out_0;
assign O_1 = hydrate_tArray_200_Array_8_Bit___inst0_out_1;
assign O_10 = hydrate_tArray_200_Array_8_Bit___inst0_out_10;
assign O_100 = hydrate_tArray_200_Array_8_Bit___inst0_out_100;
assign O_101 = hydrate_tArray_200_Array_8_Bit___inst0_out_101;
assign O_102 = hydrate_tArray_200_Array_8_Bit___inst0_out_102;
assign O_103 = hydrate_tArray_200_Array_8_Bit___inst0_out_103;
assign O_104 = hydrate_tArray_200_Array_8_Bit___inst0_out_104;
assign O_105 = hydrate_tArray_200_Array_8_Bit___inst0_out_105;
assign O_106 = hydrate_tArray_200_Array_8_Bit___inst0_out_106;
assign O_107 = hydrate_tArray_200_Array_8_Bit___inst0_out_107;
assign O_108 = hydrate_tArray_200_Array_8_Bit___inst0_out_108;
assign O_109 = hydrate_tArray_200_Array_8_Bit___inst0_out_109;
assign O_11 = hydrate_tArray_200_Array_8_Bit___inst0_out_11;
assign O_110 = hydrate_tArray_200_Array_8_Bit___inst0_out_110;
assign O_111 = hydrate_tArray_200_Array_8_Bit___inst0_out_111;
assign O_112 = hydrate_tArray_200_Array_8_Bit___inst0_out_112;
assign O_113 = hydrate_tArray_200_Array_8_Bit___inst0_out_113;
assign O_114 = hydrate_tArray_200_Array_8_Bit___inst0_out_114;
assign O_115 = hydrate_tArray_200_Array_8_Bit___inst0_out_115;
assign O_116 = hydrate_tArray_200_Array_8_Bit___inst0_out_116;
assign O_117 = hydrate_tArray_200_Array_8_Bit___inst0_out_117;
assign O_118 = hydrate_tArray_200_Array_8_Bit___inst0_out_118;
assign O_119 = hydrate_tArray_200_Array_8_Bit___inst0_out_119;
assign O_12 = hydrate_tArray_200_Array_8_Bit___inst0_out_12;
assign O_120 = hydrate_tArray_200_Array_8_Bit___inst0_out_120;
assign O_121 = hydrate_tArray_200_Array_8_Bit___inst0_out_121;
assign O_122 = hydrate_tArray_200_Array_8_Bit___inst0_out_122;
assign O_123 = hydrate_tArray_200_Array_8_Bit___inst0_out_123;
assign O_124 = hydrate_tArray_200_Array_8_Bit___inst0_out_124;
assign O_125 = hydrate_tArray_200_Array_8_Bit___inst0_out_125;
assign O_126 = hydrate_tArray_200_Array_8_Bit___inst0_out_126;
assign O_127 = hydrate_tArray_200_Array_8_Bit___inst0_out_127;
assign O_128 = hydrate_tArray_200_Array_8_Bit___inst0_out_128;
assign O_129 = hydrate_tArray_200_Array_8_Bit___inst0_out_129;
assign O_13 = hydrate_tArray_200_Array_8_Bit___inst0_out_13;
assign O_130 = hydrate_tArray_200_Array_8_Bit___inst0_out_130;
assign O_131 = hydrate_tArray_200_Array_8_Bit___inst0_out_131;
assign O_132 = hydrate_tArray_200_Array_8_Bit___inst0_out_132;
assign O_133 = hydrate_tArray_200_Array_8_Bit___inst0_out_133;
assign O_134 = hydrate_tArray_200_Array_8_Bit___inst0_out_134;
assign O_135 = hydrate_tArray_200_Array_8_Bit___inst0_out_135;
assign O_136 = hydrate_tArray_200_Array_8_Bit___inst0_out_136;
assign O_137 = hydrate_tArray_200_Array_8_Bit___inst0_out_137;
assign O_138 = hydrate_tArray_200_Array_8_Bit___inst0_out_138;
assign O_139 = hydrate_tArray_200_Array_8_Bit___inst0_out_139;
assign O_14 = hydrate_tArray_200_Array_8_Bit___inst0_out_14;
assign O_140 = hydrate_tArray_200_Array_8_Bit___inst0_out_140;
assign O_141 = hydrate_tArray_200_Array_8_Bit___inst0_out_141;
assign O_142 = hydrate_tArray_200_Array_8_Bit___inst0_out_142;
assign O_143 = hydrate_tArray_200_Array_8_Bit___inst0_out_143;
assign O_144 = hydrate_tArray_200_Array_8_Bit___inst0_out_144;
assign O_145 = hydrate_tArray_200_Array_8_Bit___inst0_out_145;
assign O_146 = hydrate_tArray_200_Array_8_Bit___inst0_out_146;
assign O_147 = hydrate_tArray_200_Array_8_Bit___inst0_out_147;
assign O_148 = hydrate_tArray_200_Array_8_Bit___inst0_out_148;
assign O_149 = hydrate_tArray_200_Array_8_Bit___inst0_out_149;
assign O_15 = hydrate_tArray_200_Array_8_Bit___inst0_out_15;
assign O_150 = hydrate_tArray_200_Array_8_Bit___inst0_out_150;
assign O_151 = hydrate_tArray_200_Array_8_Bit___inst0_out_151;
assign O_152 = hydrate_tArray_200_Array_8_Bit___inst0_out_152;
assign O_153 = hydrate_tArray_200_Array_8_Bit___inst0_out_153;
assign O_154 = hydrate_tArray_200_Array_8_Bit___inst0_out_154;
assign O_155 = hydrate_tArray_200_Array_8_Bit___inst0_out_155;
assign O_156 = hydrate_tArray_200_Array_8_Bit___inst0_out_156;
assign O_157 = hydrate_tArray_200_Array_8_Bit___inst0_out_157;
assign O_158 = hydrate_tArray_200_Array_8_Bit___inst0_out_158;
assign O_159 = hydrate_tArray_200_Array_8_Bit___inst0_out_159;
assign O_16 = hydrate_tArray_200_Array_8_Bit___inst0_out_16;
assign O_160 = hydrate_tArray_200_Array_8_Bit___inst0_out_160;
assign O_161 = hydrate_tArray_200_Array_8_Bit___inst0_out_161;
assign O_162 = hydrate_tArray_200_Array_8_Bit___inst0_out_162;
assign O_163 = hydrate_tArray_200_Array_8_Bit___inst0_out_163;
assign O_164 = hydrate_tArray_200_Array_8_Bit___inst0_out_164;
assign O_165 = hydrate_tArray_200_Array_8_Bit___inst0_out_165;
assign O_166 = hydrate_tArray_200_Array_8_Bit___inst0_out_166;
assign O_167 = hydrate_tArray_200_Array_8_Bit___inst0_out_167;
assign O_168 = hydrate_tArray_200_Array_8_Bit___inst0_out_168;
assign O_169 = hydrate_tArray_200_Array_8_Bit___inst0_out_169;
assign O_17 = hydrate_tArray_200_Array_8_Bit___inst0_out_17;
assign O_170 = hydrate_tArray_200_Array_8_Bit___inst0_out_170;
assign O_171 = hydrate_tArray_200_Array_8_Bit___inst0_out_171;
assign O_172 = hydrate_tArray_200_Array_8_Bit___inst0_out_172;
assign O_173 = hydrate_tArray_200_Array_8_Bit___inst0_out_173;
assign O_174 = hydrate_tArray_200_Array_8_Bit___inst0_out_174;
assign O_175 = hydrate_tArray_200_Array_8_Bit___inst0_out_175;
assign O_176 = hydrate_tArray_200_Array_8_Bit___inst0_out_176;
assign O_177 = hydrate_tArray_200_Array_8_Bit___inst0_out_177;
assign O_178 = hydrate_tArray_200_Array_8_Bit___inst0_out_178;
assign O_179 = hydrate_tArray_200_Array_8_Bit___inst0_out_179;
assign O_18 = hydrate_tArray_200_Array_8_Bit___inst0_out_18;
assign O_180 = hydrate_tArray_200_Array_8_Bit___inst0_out_180;
assign O_181 = hydrate_tArray_200_Array_8_Bit___inst0_out_181;
assign O_182 = hydrate_tArray_200_Array_8_Bit___inst0_out_182;
assign O_183 = hydrate_tArray_200_Array_8_Bit___inst0_out_183;
assign O_184 = hydrate_tArray_200_Array_8_Bit___inst0_out_184;
assign O_185 = hydrate_tArray_200_Array_8_Bit___inst0_out_185;
assign O_186 = hydrate_tArray_200_Array_8_Bit___inst0_out_186;
assign O_187 = hydrate_tArray_200_Array_8_Bit___inst0_out_187;
assign O_188 = hydrate_tArray_200_Array_8_Bit___inst0_out_188;
assign O_189 = hydrate_tArray_200_Array_8_Bit___inst0_out_189;
assign O_19 = hydrate_tArray_200_Array_8_Bit___inst0_out_19;
assign O_190 = hydrate_tArray_200_Array_8_Bit___inst0_out_190;
assign O_191 = hydrate_tArray_200_Array_8_Bit___inst0_out_191;
assign O_192 = hydrate_tArray_200_Array_8_Bit___inst0_out_192;
assign O_193 = hydrate_tArray_200_Array_8_Bit___inst0_out_193;
assign O_194 = hydrate_tArray_200_Array_8_Bit___inst0_out_194;
assign O_195 = hydrate_tArray_200_Array_8_Bit___inst0_out_195;
assign O_196 = hydrate_tArray_200_Array_8_Bit___inst0_out_196;
assign O_197 = hydrate_tArray_200_Array_8_Bit___inst0_out_197;
assign O_198 = hydrate_tArray_200_Array_8_Bit___inst0_out_198;
assign O_199 = hydrate_tArray_200_Array_8_Bit___inst0_out_199;
assign O_2 = hydrate_tArray_200_Array_8_Bit___inst0_out_2;
assign O_20 = hydrate_tArray_200_Array_8_Bit___inst0_out_20;
assign O_21 = hydrate_tArray_200_Array_8_Bit___inst0_out_21;
assign O_22 = hydrate_tArray_200_Array_8_Bit___inst0_out_22;
assign O_23 = hydrate_tArray_200_Array_8_Bit___inst0_out_23;
assign O_24 = hydrate_tArray_200_Array_8_Bit___inst0_out_24;
assign O_25 = hydrate_tArray_200_Array_8_Bit___inst0_out_25;
assign O_26 = hydrate_tArray_200_Array_8_Bit___inst0_out_26;
assign O_27 = hydrate_tArray_200_Array_8_Bit___inst0_out_27;
assign O_28 = hydrate_tArray_200_Array_8_Bit___inst0_out_28;
assign O_29 = hydrate_tArray_200_Array_8_Bit___inst0_out_29;
assign O_3 = hydrate_tArray_200_Array_8_Bit___inst0_out_3;
assign O_30 = hydrate_tArray_200_Array_8_Bit___inst0_out_30;
assign O_31 = hydrate_tArray_200_Array_8_Bit___inst0_out_31;
assign O_32 = hydrate_tArray_200_Array_8_Bit___inst0_out_32;
assign O_33 = hydrate_tArray_200_Array_8_Bit___inst0_out_33;
assign O_34 = hydrate_tArray_200_Array_8_Bit___inst0_out_34;
assign O_35 = hydrate_tArray_200_Array_8_Bit___inst0_out_35;
assign O_36 = hydrate_tArray_200_Array_8_Bit___inst0_out_36;
assign O_37 = hydrate_tArray_200_Array_8_Bit___inst0_out_37;
assign O_38 = hydrate_tArray_200_Array_8_Bit___inst0_out_38;
assign O_39 = hydrate_tArray_200_Array_8_Bit___inst0_out_39;
assign O_4 = hydrate_tArray_200_Array_8_Bit___inst0_out_4;
assign O_40 = hydrate_tArray_200_Array_8_Bit___inst0_out_40;
assign O_41 = hydrate_tArray_200_Array_8_Bit___inst0_out_41;
assign O_42 = hydrate_tArray_200_Array_8_Bit___inst0_out_42;
assign O_43 = hydrate_tArray_200_Array_8_Bit___inst0_out_43;
assign O_44 = hydrate_tArray_200_Array_8_Bit___inst0_out_44;
assign O_45 = hydrate_tArray_200_Array_8_Bit___inst0_out_45;
assign O_46 = hydrate_tArray_200_Array_8_Bit___inst0_out_46;
assign O_47 = hydrate_tArray_200_Array_8_Bit___inst0_out_47;
assign O_48 = hydrate_tArray_200_Array_8_Bit___inst0_out_48;
assign O_49 = hydrate_tArray_200_Array_8_Bit___inst0_out_49;
assign O_5 = hydrate_tArray_200_Array_8_Bit___inst0_out_5;
assign O_50 = hydrate_tArray_200_Array_8_Bit___inst0_out_50;
assign O_51 = hydrate_tArray_200_Array_8_Bit___inst0_out_51;
assign O_52 = hydrate_tArray_200_Array_8_Bit___inst0_out_52;
assign O_53 = hydrate_tArray_200_Array_8_Bit___inst0_out_53;
assign O_54 = hydrate_tArray_200_Array_8_Bit___inst0_out_54;
assign O_55 = hydrate_tArray_200_Array_8_Bit___inst0_out_55;
assign O_56 = hydrate_tArray_200_Array_8_Bit___inst0_out_56;
assign O_57 = hydrate_tArray_200_Array_8_Bit___inst0_out_57;
assign O_58 = hydrate_tArray_200_Array_8_Bit___inst0_out_58;
assign O_59 = hydrate_tArray_200_Array_8_Bit___inst0_out_59;
assign O_6 = hydrate_tArray_200_Array_8_Bit___inst0_out_6;
assign O_60 = hydrate_tArray_200_Array_8_Bit___inst0_out_60;
assign O_61 = hydrate_tArray_200_Array_8_Bit___inst0_out_61;
assign O_62 = hydrate_tArray_200_Array_8_Bit___inst0_out_62;
assign O_63 = hydrate_tArray_200_Array_8_Bit___inst0_out_63;
assign O_64 = hydrate_tArray_200_Array_8_Bit___inst0_out_64;
assign O_65 = hydrate_tArray_200_Array_8_Bit___inst0_out_65;
assign O_66 = hydrate_tArray_200_Array_8_Bit___inst0_out_66;
assign O_67 = hydrate_tArray_200_Array_8_Bit___inst0_out_67;
assign O_68 = hydrate_tArray_200_Array_8_Bit___inst0_out_68;
assign O_69 = hydrate_tArray_200_Array_8_Bit___inst0_out_69;
assign O_7 = hydrate_tArray_200_Array_8_Bit___inst0_out_7;
assign O_70 = hydrate_tArray_200_Array_8_Bit___inst0_out_70;
assign O_71 = hydrate_tArray_200_Array_8_Bit___inst0_out_71;
assign O_72 = hydrate_tArray_200_Array_8_Bit___inst0_out_72;
assign O_73 = hydrate_tArray_200_Array_8_Bit___inst0_out_73;
assign O_74 = hydrate_tArray_200_Array_8_Bit___inst0_out_74;
assign O_75 = hydrate_tArray_200_Array_8_Bit___inst0_out_75;
assign O_76 = hydrate_tArray_200_Array_8_Bit___inst0_out_76;
assign O_77 = hydrate_tArray_200_Array_8_Bit___inst0_out_77;
assign O_78 = hydrate_tArray_200_Array_8_Bit___inst0_out_78;
assign O_79 = hydrate_tArray_200_Array_8_Bit___inst0_out_79;
assign O_8 = hydrate_tArray_200_Array_8_Bit___inst0_out_8;
assign O_80 = hydrate_tArray_200_Array_8_Bit___inst0_out_80;
assign O_81 = hydrate_tArray_200_Array_8_Bit___inst0_out_81;
assign O_82 = hydrate_tArray_200_Array_8_Bit___inst0_out_82;
assign O_83 = hydrate_tArray_200_Array_8_Bit___inst0_out_83;
assign O_84 = hydrate_tArray_200_Array_8_Bit___inst0_out_84;
assign O_85 = hydrate_tArray_200_Array_8_Bit___inst0_out_85;
assign O_86 = hydrate_tArray_200_Array_8_Bit___inst0_out_86;
assign O_87 = hydrate_tArray_200_Array_8_Bit___inst0_out_87;
assign O_88 = hydrate_tArray_200_Array_8_Bit___inst0_out_88;
assign O_89 = hydrate_tArray_200_Array_8_Bit___inst0_out_89;
assign O_9 = hydrate_tArray_200_Array_8_Bit___inst0_out_9;
assign O_90 = hydrate_tArray_200_Array_8_Bit___inst0_out_90;
assign O_91 = hydrate_tArray_200_Array_8_Bit___inst0_out_91;
assign O_92 = hydrate_tArray_200_Array_8_Bit___inst0_out_92;
assign O_93 = hydrate_tArray_200_Array_8_Bit___inst0_out_93;
assign O_94 = hydrate_tArray_200_Array_8_Bit___inst0_out_94;
assign O_95 = hydrate_tArray_200_Array_8_Bit___inst0_out_95;
assign O_96 = hydrate_tArray_200_Array_8_Bit___inst0_out_96;
assign O_97 = hydrate_tArray_200_Array_8_Bit___inst0_out_97;
assign O_98 = hydrate_tArray_200_Array_8_Bit___inst0_out_98;
assign O_99 = hydrate_tArray_200_Array_8_Bit___inst0_out_99;
endmodule

module Register1 (input CLK/*verilator public*/, input [0:0] I/*verilator public*/, output [0:0] O/*verilator public*/);
wire DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0(.CLK(CLK), .I(I[0]), .O(DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O));
assign O = DFF_init0_has_ceFalse_has_resetFalse_has_async_resetFalse_inst0_O;
endmodule

module Register_Bitt_0init_FalseCE_FalseRESET (input CLK/*verilator public*/, input I/*verilator public*/, output O/*verilator public*/);
wire [0:0] Register1_inst0_O;
wire [0:0] dehydrate_tBit_inst0_out;
wire hydrate_tBit_inst0_out;
Register1 Register1_inst0(.CLK(CLK), .I(dehydrate_tBit_inst0_out), .O(Register1_inst0_O));
\aetherlinglib_dehydrate__hydratedTypeBit dehydrate_tBit_inst0(.in(I), .out(dehydrate_tBit_inst0_out));
\aetherlinglib_hydrate__hydratedTypeBit hydrate_tBit_inst0(.in(Register1_inst0_O), .out(hydrate_tBit_inst0_out));
assign O = hydrate_tBit_inst0_out;
endmodule

module FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_100/*verilator public*/, input [7:0] I_101/*verilator public*/, input [7:0] I_102/*verilator public*/, input [7:0] I_103/*verilator public*/, input [7:0] I_104/*verilator public*/, input [7:0] I_105/*verilator public*/, input [7:0] I_106/*verilator public*/, input [7:0] I_107/*verilator public*/, input [7:0] I_108/*verilator public*/, input [7:0] I_109/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_110/*verilator public*/, input [7:0] I_111/*verilator public*/, input [7:0] I_112/*verilator public*/, input [7:0] I_113/*verilator public*/, input [7:0] I_114/*verilator public*/, input [7:0] I_115/*verilator public*/, input [7:0] I_116/*verilator public*/, input [7:0] I_117/*verilator public*/, input [7:0] I_118/*verilator public*/, input [7:0] I_119/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_120/*verilator public*/, input [7:0] I_121/*verilator public*/, input [7:0] I_122/*verilator public*/, input [7:0] I_123/*verilator public*/, input [7:0] I_124/*verilator public*/, input [7:0] I_125/*verilator public*/, input [7:0] I_126/*verilator public*/, input [7:0] I_127/*verilator public*/, input [7:0] I_128/*verilator public*/, input [7:0] I_129/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_130/*verilator public*/, input [7:0] I_131/*verilator public*/, input [7:0] I_132/*verilator public*/, input [7:0] I_133/*verilator public*/, input [7:0] I_134/*verilator public*/, input [7:0] I_135/*verilator public*/, input [7:0] I_136/*verilator public*/, input [7:0] I_137/*verilator public*/, input [7:0] I_138/*verilator public*/, input [7:0] I_139/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_140/*verilator public*/, input [7:0] I_141/*verilator public*/, input [7:0] I_142/*verilator public*/, input [7:0] I_143/*verilator public*/, input [7:0] I_144/*verilator public*/, input [7:0] I_145/*verilator public*/, input [7:0] I_146/*verilator public*/, input [7:0] I_147/*verilator public*/, input [7:0] I_148/*verilator public*/, input [7:0] I_149/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_150/*verilator public*/, input [7:0] I_151/*verilator public*/, input [7:0] I_152/*verilator public*/, input [7:0] I_153/*verilator public*/, input [7:0] I_154/*verilator public*/, input [7:0] I_155/*verilator public*/, input [7:0] I_156/*verilator public*/, input [7:0] I_157/*verilator public*/, input [7:0] I_158/*verilator public*/, input [7:0] I_159/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_160/*verilator public*/, input [7:0] I_161/*verilator public*/, input [7:0] I_162/*verilator public*/, input [7:0] I_163/*verilator public*/, input [7:0] I_164/*verilator public*/, input [7:0] I_165/*verilator public*/, input [7:0] I_166/*verilator public*/, input [7:0] I_167/*verilator public*/, input [7:0] I_168/*verilator public*/, input [7:0] I_169/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_170/*verilator public*/, input [7:0] I_171/*verilator public*/, input [7:0] I_172/*verilator public*/, input [7:0] I_173/*verilator public*/, input [7:0] I_174/*verilator public*/, input [7:0] I_175/*verilator public*/, input [7:0] I_176/*verilator public*/, input [7:0] I_177/*verilator public*/, input [7:0] I_178/*verilator public*/, input [7:0] I_179/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_180/*verilator public*/, input [7:0] I_181/*verilator public*/, input [7:0] I_182/*verilator public*/, input [7:0] I_183/*verilator public*/, input [7:0] I_184/*verilator public*/, input [7:0] I_185/*verilator public*/, input [7:0] I_186/*verilator public*/, input [7:0] I_187/*verilator public*/, input [7:0] I_188/*verilator public*/, input [7:0] I_189/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_190/*verilator public*/, input [7:0] I_191/*verilator public*/, input [7:0] I_192/*verilator public*/, input [7:0] I_193/*verilator public*/, input [7:0] I_194/*verilator public*/, input [7:0] I_195/*verilator public*/, input [7:0] I_196/*verilator public*/, input [7:0] I_197/*verilator public*/, input [7:0] I_198/*verilator public*/, input [7:0] I_199/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_40/*verilator public*/, input [7:0] I_41/*verilator public*/, input [7:0] I_42/*verilator public*/, input [7:0] I_43/*verilator public*/, input [7:0] I_44/*verilator public*/, input [7:0] I_45/*verilator public*/, input [7:0] I_46/*verilator public*/, input [7:0] I_47/*verilator public*/, input [7:0] I_48/*verilator public*/, input [7:0] I_49/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_50/*verilator public*/, input [7:0] I_51/*verilator public*/, input [7:0] I_52/*verilator public*/, input [7:0] I_53/*verilator public*/, input [7:0] I_54/*verilator public*/, input [7:0] I_55/*verilator public*/, input [7:0] I_56/*verilator public*/, input [7:0] I_57/*verilator public*/, input [7:0] I_58/*verilator public*/, input [7:0] I_59/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_60/*verilator public*/, input [7:0] I_61/*verilator public*/, input [7:0] I_62/*verilator public*/, input [7:0] I_63/*verilator public*/, input [7:0] I_64/*verilator public*/, input [7:0] I_65/*verilator public*/, input [7:0] I_66/*verilator public*/, input [7:0] I_67/*verilator public*/, input [7:0] I_68/*verilator public*/, input [7:0] I_69/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_70/*verilator public*/, input [7:0] I_71/*verilator public*/, input [7:0] I_72/*verilator public*/, input [7:0] I_73/*verilator public*/, input [7:0] I_74/*verilator public*/, input [7:0] I_75/*verilator public*/, input [7:0] I_76/*verilator public*/, input [7:0] I_77/*verilator public*/, input [7:0] I_78/*verilator public*/, input [7:0] I_79/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_80/*verilator public*/, input [7:0] I_81/*verilator public*/, input [7:0] I_82/*verilator public*/, input [7:0] I_83/*verilator public*/, input [7:0] I_84/*verilator public*/, input [7:0] I_85/*verilator public*/, input [7:0] I_86/*verilator public*/, input [7:0] I_87/*verilator public*/, input [7:0] I_88/*verilator public*/, input [7:0] I_89/*verilator public*/, input [7:0] I_9/*verilator public*/, input [7:0] I_90/*verilator public*/, input [7:0] I_91/*verilator public*/, input [7:0] I_92/*verilator public*/, input [7:0] I_93/*verilator public*/, input [7:0] I_94/*verilator public*/, input [7:0] I_95/*verilator public*/, input [7:0] I_96/*verilator public*/, input [7:0] I_97/*verilator public*/, input [7:0] I_98/*verilator public*/, input [7:0] I_99/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_100/*verilator public*/, output [7:0] O_101/*verilator public*/, output [7:0] O_102/*verilator public*/, output [7:0] O_103/*verilator public*/, output [7:0] O_104/*verilator public*/, output [7:0] O_105/*verilator public*/, output [7:0] O_106/*verilator public*/, output [7:0] O_107/*verilator public*/, output [7:0] O_108/*verilator public*/, output [7:0] O_109/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_110/*verilator public*/, output [7:0] O_111/*verilator public*/, output [7:0] O_112/*verilator public*/, output [7:0] O_113/*verilator public*/, output [7:0] O_114/*verilator public*/, output [7:0] O_115/*verilator public*/, output [7:0] O_116/*verilator public*/, output [7:0] O_117/*verilator public*/, output [7:0] O_118/*verilator public*/, output [7:0] O_119/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_120/*verilator public*/, output [7:0] O_121/*verilator public*/, output [7:0] O_122/*verilator public*/, output [7:0] O_123/*verilator public*/, output [7:0] O_124/*verilator public*/, output [7:0] O_125/*verilator public*/, output [7:0] O_126/*verilator public*/, output [7:0] O_127/*verilator public*/, output [7:0] O_128/*verilator public*/, output [7:0] O_129/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_130/*verilator public*/, output [7:0] O_131/*verilator public*/, output [7:0] O_132/*verilator public*/, output [7:0] O_133/*verilator public*/, output [7:0] O_134/*verilator public*/, output [7:0] O_135/*verilator public*/, output [7:0] O_136/*verilator public*/, output [7:0] O_137/*verilator public*/, output [7:0] O_138/*verilator public*/, output [7:0] O_139/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_140/*verilator public*/, output [7:0] O_141/*verilator public*/, output [7:0] O_142/*verilator public*/, output [7:0] O_143/*verilator public*/, output [7:0] O_144/*verilator public*/, output [7:0] O_145/*verilator public*/, output [7:0] O_146/*verilator public*/, output [7:0] O_147/*verilator public*/, output [7:0] O_148/*verilator public*/, output [7:0] O_149/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_150/*verilator public*/, output [7:0] O_151/*verilator public*/, output [7:0] O_152/*verilator public*/, output [7:0] O_153/*verilator public*/, output [7:0] O_154/*verilator public*/, output [7:0] O_155/*verilator public*/, output [7:0] O_156/*verilator public*/, output [7:0] O_157/*verilator public*/, output [7:0] O_158/*verilator public*/, output [7:0] O_159/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_160/*verilator public*/, output [7:0] O_161/*verilator public*/, output [7:0] O_162/*verilator public*/, output [7:0] O_163/*verilator public*/, output [7:0] O_164/*verilator public*/, output [7:0] O_165/*verilator public*/, output [7:0] O_166/*verilator public*/, output [7:0] O_167/*verilator public*/, output [7:0] O_168/*verilator public*/, output [7:0] O_169/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_170/*verilator public*/, output [7:0] O_171/*verilator public*/, output [7:0] O_172/*verilator public*/, output [7:0] O_173/*verilator public*/, output [7:0] O_174/*verilator public*/, output [7:0] O_175/*verilator public*/, output [7:0] O_176/*verilator public*/, output [7:0] O_177/*verilator public*/, output [7:0] O_178/*verilator public*/, output [7:0] O_179/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_180/*verilator public*/, output [7:0] O_181/*verilator public*/, output [7:0] O_182/*verilator public*/, output [7:0] O_183/*verilator public*/, output [7:0] O_184/*verilator public*/, output [7:0] O_185/*verilator public*/, output [7:0] O_186/*verilator public*/, output [7:0] O_187/*verilator public*/, output [7:0] O_188/*verilator public*/, output [7:0] O_189/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_190/*verilator public*/, output [7:0] O_191/*verilator public*/, output [7:0] O_192/*verilator public*/, output [7:0] O_193/*verilator public*/, output [7:0] O_194/*verilator public*/, output [7:0] O_195/*verilator public*/, output [7:0] O_196/*verilator public*/, output [7:0] O_197/*verilator public*/, output [7:0] O_198/*verilator public*/, output [7:0] O_199/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_40/*verilator public*/, output [7:0] O_41/*verilator public*/, output [7:0] O_42/*verilator public*/, output [7:0] O_43/*verilator public*/, output [7:0] O_44/*verilator public*/, output [7:0] O_45/*verilator public*/, output [7:0] O_46/*verilator public*/, output [7:0] O_47/*verilator public*/, output [7:0] O_48/*verilator public*/, output [7:0] O_49/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_50/*verilator public*/, output [7:0] O_51/*verilator public*/, output [7:0] O_52/*verilator public*/, output [7:0] O_53/*verilator public*/, output [7:0] O_54/*verilator public*/, output [7:0] O_55/*verilator public*/, output [7:0] O_56/*verilator public*/, output [7:0] O_57/*verilator public*/, output [7:0] O_58/*verilator public*/, output [7:0] O_59/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_60/*verilator public*/, output [7:0] O_61/*verilator public*/, output [7:0] O_62/*verilator public*/, output [7:0] O_63/*verilator public*/, output [7:0] O_64/*verilator public*/, output [7:0] O_65/*verilator public*/, output [7:0] O_66/*verilator public*/, output [7:0] O_67/*verilator public*/, output [7:0] O_68/*verilator public*/, output [7:0] O_69/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_70/*verilator public*/, output [7:0] O_71/*verilator public*/, output [7:0] O_72/*verilator public*/, output [7:0] O_73/*verilator public*/, output [7:0] O_74/*verilator public*/, output [7:0] O_75/*verilator public*/, output [7:0] O_76/*verilator public*/, output [7:0] O_77/*verilator public*/, output [7:0] O_78/*verilator public*/, output [7:0] O_79/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_80/*verilator public*/, output [7:0] O_81/*verilator public*/, output [7:0] O_82/*verilator public*/, output [7:0] O_83/*verilator public*/, output [7:0] O_84/*verilator public*/, output [7:0] O_85/*verilator public*/, output [7:0] O_86/*verilator public*/, output [7:0] O_87/*verilator public*/, output [7:0] O_88/*verilator public*/, output [7:0] O_89/*verilator public*/, output [7:0] O_9/*verilator public*/, output [7:0] O_90/*verilator public*/, output [7:0] O_91/*verilator public*/, output [7:0] O_92/*verilator public*/, output [7:0] O_93/*verilator public*/, output [7:0] O_94/*verilator public*/, output [7:0] O_95/*verilator public*/, output [7:0] O_96/*verilator public*/, output [7:0] O_97/*verilator public*/, output [7:0] O_98/*verilator public*/, output [7:0] O_99/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_100;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_101;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_102;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_103;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_104;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_105;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_106;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_107;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_108;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_109;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_110;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_111;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_112;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_113;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_114;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_115;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_116;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_117;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_118;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_119;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_120;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_121;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_122;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_123;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_124;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_125;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_126;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_127;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_128;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_129;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_130;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_131;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_132;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_133;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_134;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_135;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_136;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_137;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_138;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_139;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_140;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_141;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_142;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_143;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_144;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_145;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_146;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_147;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_148;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_149;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_150;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_151;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_152;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_153;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_154;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_155;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_156;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_157;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_158;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_159;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_160;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_161;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_162;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_163;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_164;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_165;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_166;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_167;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_168;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_169;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_170;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_171;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_172;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_173;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_174;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_175;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_176;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_177;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_178;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_179;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_180;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_181;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_182;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_183;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_184;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_185;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_186;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_187;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_188;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_189;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_190;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_191;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_192;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_193;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_194;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_195;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_196;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_197;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_198;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_199;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_40;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_41;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_42;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_43;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_44;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_45;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_46;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_47;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_48;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_49;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_50;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_51;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_52;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_53;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_54;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_55;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_56;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_57;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_58;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_59;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_60;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_61;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_62;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_63;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_64;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_65;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_66;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_67;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_68;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_69;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_70;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_71;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_72;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_73;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_74;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_75;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_76;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_77;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_78;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_79;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_80;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_81;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_82;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_83;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_84;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_85;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_86;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_87;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_88;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_89;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_90;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_91;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_92;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_93;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_94;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_95;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_96;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_97;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_98;
wire [7:0] Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_99;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I_0(I_0), .I_1(I_1), .I_10(I_10), .I_100(I_100), .I_101(I_101), .I_102(I_102), .I_103(I_103), .I_104(I_104), .I_105(I_105), .I_106(I_106), .I_107(I_107), .I_108(I_108), .I_109(I_109), .I_11(I_11), .I_110(I_110), .I_111(I_111), .I_112(I_112), .I_113(I_113), .I_114(I_114), .I_115(I_115), .I_116(I_116), .I_117(I_117), .I_118(I_118), .I_119(I_119), .I_12(I_12), .I_120(I_120), .I_121(I_121), .I_122(I_122), .I_123(I_123), .I_124(I_124), .I_125(I_125), .I_126(I_126), .I_127(I_127), .I_128(I_128), .I_129(I_129), .I_13(I_13), .I_130(I_130), .I_131(I_131), .I_132(I_132), .I_133(I_133), .I_134(I_134), .I_135(I_135), .I_136(I_136), .I_137(I_137), .I_138(I_138), .I_139(I_139), .I_14(I_14), .I_140(I_140), .I_141(I_141), .I_142(I_142), .I_143(I_143), .I_144(I_144), .I_145(I_145), .I_146(I_146), .I_147(I_147), .I_148(I_148), .I_149(I_149), .I_15(I_15), .I_150(I_150), .I_151(I_151), .I_152(I_152), .I_153(I_153), .I_154(I_154), .I_155(I_155), .I_156(I_156), .I_157(I_157), .I_158(I_158), .I_159(I_159), .I_16(I_16), .I_160(I_160), .I_161(I_161), .I_162(I_162), .I_163(I_163), .I_164(I_164), .I_165(I_165), .I_166(I_166), .I_167(I_167), .I_168(I_168), .I_169(I_169), .I_17(I_17), .I_170(I_170), .I_171(I_171), .I_172(I_172), .I_173(I_173), .I_174(I_174), .I_175(I_175), .I_176(I_176), .I_177(I_177), .I_178(I_178), .I_179(I_179), .I_18(I_18), .I_180(I_180), .I_181(I_181), .I_182(I_182), .I_183(I_183), .I_184(I_184), .I_185(I_185), .I_186(I_186), .I_187(I_187), .I_188(I_188), .I_189(I_189), .I_19(I_19), .I_190(I_190), .I_191(I_191), .I_192(I_192), .I_193(I_193), .I_194(I_194), .I_195(I_195), .I_196(I_196), .I_197(I_197), .I_198(I_198), .I_199(I_199), .I_2(I_2), .I_20(I_20), .I_21(I_21), .I_22(I_22), .I_23(I_23), .I_24(I_24), .I_25(I_25), .I_26(I_26), .I_27(I_27), .I_28(I_28), .I_29(I_29), .I_3(I_3), .I_30(I_30), .I_31(I_31), .I_32(I_32), .I_33(I_33), .I_34(I_34), .I_35(I_35), .I_36(I_36), .I_37(I_37), .I_38(I_38), .I_39(I_39), .I_4(I_4), .I_40(I_40), .I_41(I_41), .I_42(I_42), .I_43(I_43), .I_44(I_44), .I_45(I_45), .I_46(I_46), .I_47(I_47), .I_48(I_48), .I_49(I_49), .I_5(I_5), .I_50(I_50), .I_51(I_51), .I_52(I_52), .I_53(I_53), .I_54(I_54), .I_55(I_55), .I_56(I_56), .I_57(I_57), .I_58(I_58), .I_59(I_59), .I_6(I_6), .I_60(I_60), .I_61(I_61), .I_62(I_62), .I_63(I_63), .I_64(I_64), .I_65(I_65), .I_66(I_66), .I_67(I_67), .I_68(I_68), .I_69(I_69), .I_7(I_7), .I_70(I_70), .I_71(I_71), .I_72(I_72), .I_73(I_73), .I_74(I_74), .I_75(I_75), .I_76(I_76), .I_77(I_77), .I_78(I_78), .I_79(I_79), .I_8(I_8), .I_80(I_80), .I_81(I_81), .I_82(I_82), .I_83(I_83), .I_84(I_84), .I_85(I_85), .I_86(I_86), .I_87(I_87), .I_88(I_88), .I_89(I_89), .I_9(I_9), .I_90(I_90), .I_91(I_91), .I_92(I_92), .I_93(I_93), .I_94(I_94), .I_95(I_95), .I_96(I_96), .I_97(I_97), .I_98(I_98), .I_99(I_99), .O_0(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0), .O_1(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1), .O_10(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10), .O_100(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_100), .O_101(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_101), .O_102(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_102), .O_103(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_103), .O_104(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_104), .O_105(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_105), .O_106(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_106), .O_107(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_107), .O_108(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_108), .O_109(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_109), .O_11(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11), .O_110(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_110), .O_111(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_111), .O_112(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_112), .O_113(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_113), .O_114(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_114), .O_115(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_115), .O_116(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_116), .O_117(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_117), .O_118(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_118), .O_119(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_119), .O_12(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12), .O_120(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_120), .O_121(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_121), .O_122(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_122), .O_123(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_123), .O_124(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_124), .O_125(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_125), .O_126(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_126), .O_127(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_127), .O_128(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_128), .O_129(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_129), .O_13(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13), .O_130(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_130), .O_131(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_131), .O_132(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_132), .O_133(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_133), .O_134(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_134), .O_135(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_135), .O_136(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_136), .O_137(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_137), .O_138(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_138), .O_139(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_139), .O_14(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14), .O_140(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_140), .O_141(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_141), .O_142(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_142), .O_143(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_143), .O_144(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_144), .O_145(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_145), .O_146(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_146), .O_147(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_147), .O_148(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_148), .O_149(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_149), .O_15(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15), .O_150(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_150), .O_151(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_151), .O_152(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_152), .O_153(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_153), .O_154(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_154), .O_155(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_155), .O_156(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_156), .O_157(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_157), .O_158(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_158), .O_159(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_159), .O_16(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16), .O_160(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_160), .O_161(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_161), .O_162(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_162), .O_163(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_163), .O_164(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_164), .O_165(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_165), .O_166(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_166), .O_167(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_167), .O_168(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_168), .O_169(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_169), .O_17(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17), .O_170(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_170), .O_171(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_171), .O_172(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_172), .O_173(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_173), .O_174(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_174), .O_175(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_175), .O_176(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_176), .O_177(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_177), .O_178(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_178), .O_179(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_179), .O_18(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18), .O_180(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_180), .O_181(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_181), .O_182(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_182), .O_183(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_183), .O_184(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_184), .O_185(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_185), .O_186(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_186), .O_187(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_187), .O_188(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_188), .O_189(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_189), .O_19(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19), .O_190(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_190), .O_191(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_191), .O_192(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_192), .O_193(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_193), .O_194(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_194), .O_195(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_195), .O_196(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_196), .O_197(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_197), .O_198(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_198), .O_199(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_199), .O_2(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2), .O_20(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20), .O_21(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21), .O_22(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22), .O_23(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23), .O_24(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24), .O_25(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25), .O_26(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26), .O_27(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27), .O_28(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28), .O_29(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29), .O_3(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3), .O_30(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30), .O_31(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31), .O_32(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32), .O_33(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33), .O_34(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34), .O_35(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35), .O_36(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36), .O_37(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37), .O_38(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38), .O_39(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39), .O_4(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4), .O_40(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_40), .O_41(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_41), .O_42(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_42), .O_43(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_43), .O_44(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_44), .O_45(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_45), .O_46(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_46), .O_47(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_47), .O_48(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_48), .O_49(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_49), .O_5(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5), .O_50(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_50), .O_51(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_51), .O_52(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_52), .O_53(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_53), .O_54(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_54), .O_55(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_55), .O_56(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_56), .O_57(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_57), .O_58(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_58), .O_59(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_59), .O_6(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6), .O_60(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_60), .O_61(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_61), .O_62(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_62), .O_63(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_63), .O_64(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_64), .O_65(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_65), .O_66(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_66), .O_67(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_67), .O_68(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_68), .O_69(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_69), .O_7(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7), .O_70(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_70), .O_71(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_71), .O_72(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_72), .O_73(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_73), .O_74(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_74), .O_75(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_75), .O_76(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_76), .O_77(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_77), .O_78(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_78), .O_79(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_79), .O_8(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8), .O_80(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_80), .O_81(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_81), .O_82(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_82), .O_83(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_83), .O_84(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_84), .O_85(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_85), .O_86(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_86), .O_87(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_87), .O_88(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_88), .O_89(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_89), .O_9(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9), .O_90(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_90), .O_91(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_91), .O_92(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_92), .O_93(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_93), .O_94(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_94), .O_95(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_95), .O_96(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_96), .O_97(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_97), .O_98(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_98), .O_99(Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_99));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O_0 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_0;
assign O_1 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_1;
assign O_10 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_10;
assign O_100 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_100;
assign O_101 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_101;
assign O_102 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_102;
assign O_103 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_103;
assign O_104 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_104;
assign O_105 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_105;
assign O_106 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_106;
assign O_107 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_107;
assign O_108 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_108;
assign O_109 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_109;
assign O_11 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_11;
assign O_110 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_110;
assign O_111 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_111;
assign O_112 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_112;
assign O_113 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_113;
assign O_114 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_114;
assign O_115 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_115;
assign O_116 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_116;
assign O_117 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_117;
assign O_118 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_118;
assign O_119 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_119;
assign O_12 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_12;
assign O_120 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_120;
assign O_121 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_121;
assign O_122 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_122;
assign O_123 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_123;
assign O_124 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_124;
assign O_125 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_125;
assign O_126 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_126;
assign O_127 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_127;
assign O_128 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_128;
assign O_129 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_129;
assign O_13 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_13;
assign O_130 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_130;
assign O_131 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_131;
assign O_132 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_132;
assign O_133 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_133;
assign O_134 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_134;
assign O_135 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_135;
assign O_136 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_136;
assign O_137 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_137;
assign O_138 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_138;
assign O_139 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_139;
assign O_14 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_14;
assign O_140 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_140;
assign O_141 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_141;
assign O_142 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_142;
assign O_143 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_143;
assign O_144 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_144;
assign O_145 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_145;
assign O_146 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_146;
assign O_147 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_147;
assign O_148 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_148;
assign O_149 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_149;
assign O_15 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_15;
assign O_150 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_150;
assign O_151 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_151;
assign O_152 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_152;
assign O_153 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_153;
assign O_154 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_154;
assign O_155 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_155;
assign O_156 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_156;
assign O_157 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_157;
assign O_158 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_158;
assign O_159 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_159;
assign O_16 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_16;
assign O_160 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_160;
assign O_161 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_161;
assign O_162 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_162;
assign O_163 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_163;
assign O_164 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_164;
assign O_165 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_165;
assign O_166 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_166;
assign O_167 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_167;
assign O_168 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_168;
assign O_169 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_169;
assign O_17 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_17;
assign O_170 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_170;
assign O_171 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_171;
assign O_172 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_172;
assign O_173 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_173;
assign O_174 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_174;
assign O_175 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_175;
assign O_176 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_176;
assign O_177 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_177;
assign O_178 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_178;
assign O_179 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_179;
assign O_18 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_18;
assign O_180 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_180;
assign O_181 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_181;
assign O_182 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_182;
assign O_183 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_183;
assign O_184 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_184;
assign O_185 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_185;
assign O_186 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_186;
assign O_187 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_187;
assign O_188 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_188;
assign O_189 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_189;
assign O_19 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_19;
assign O_190 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_190;
assign O_191 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_191;
assign O_192 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_192;
assign O_193 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_193;
assign O_194 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_194;
assign O_195 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_195;
assign O_196 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_196;
assign O_197 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_197;
assign O_198 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_198;
assign O_199 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_199;
assign O_2 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_2;
assign O_20 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_20;
assign O_21 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_21;
assign O_22 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_22;
assign O_23 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_23;
assign O_24 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_24;
assign O_25 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_25;
assign O_26 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_26;
assign O_27 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_27;
assign O_28 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_28;
assign O_29 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_29;
assign O_3 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_3;
assign O_30 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_30;
assign O_31 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_31;
assign O_32 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_32;
assign O_33 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_33;
assign O_34 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_34;
assign O_35 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_35;
assign O_36 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_36;
assign O_37 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_37;
assign O_38 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_38;
assign O_39 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_39;
assign O_4 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_4;
assign O_40 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_40;
assign O_41 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_41;
assign O_42 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_42;
assign O_43 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_43;
assign O_44 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_44;
assign O_45 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_45;
assign O_46 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_46;
assign O_47 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_47;
assign O_48 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_48;
assign O_49 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_49;
assign O_5 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_5;
assign O_50 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_50;
assign O_51 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_51;
assign O_52 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_52;
assign O_53 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_53;
assign O_54 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_54;
assign O_55 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_55;
assign O_56 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_56;
assign O_57 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_57;
assign O_58 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_58;
assign O_59 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_59;
assign O_6 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_6;
assign O_60 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_60;
assign O_61 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_61;
assign O_62 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_62;
assign O_63 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_63;
assign O_64 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_64;
assign O_65 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_65;
assign O_66 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_66;
assign O_67 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_67;
assign O_68 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_68;
assign O_69 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_69;
assign O_7 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_7;
assign O_70 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_70;
assign O_71 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_71;
assign O_72 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_72;
assign O_73 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_73;
assign O_74 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_74;
assign O_75 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_75;
assign O_76 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_76;
assign O_77 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_77;
assign O_78 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_78;
assign O_79 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_79;
assign O_8 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_8;
assign O_80 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_80;
assign O_81 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_81;
assign O_82 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_82;
assign O_83 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_83;
assign O_84 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_84;
assign O_85 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_85;
assign O_86 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_86;
assign O_87 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_87;
assign O_88 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_88;
assign O_89 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_89;
assign O_9 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_9;
assign O_90 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_90;
assign O_91 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_91;
assign O_92 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_92;
assign O_93 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_93;
assign O_94 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_94;
assign O_95 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_95;
assign O_96 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_96;
assign O_97 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_97;
assign O_98 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_98;
assign O_99 = Register_Array_200_Array_8_Bit__t_0init_FalseCE_FalseRESET_inst0_O_99;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
wire Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
Register_Array_8_Bit_t_0init_FalseCE_FalseRESET Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(I), .O(Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O));
Register_Bitt_0init_FalseCE_FalseRESET Register_Bitt_0init_FalseCE_FalseRESET_inst0(.CLK(CLK), .I(valid_up), .O(Register_Bitt_0init_FalseCE_FalseRESET_inst0_O));
assign O = Register_Array_8_Bit_t_0init_FalseCE_FalseRESET_inst0_O;
assign valid_down = Register_Bitt_0init_FalseCE_FalseRESET_inst0_O;
endmodule

module Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue (input CLK/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] LUT_Array_8_Bit_t_1n_inst0_data;
wire [0:0] SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O;
wire [0:0] coreir_const11_inst0_out;
LUT_Array_8_Bit_t_1n LUT_Array_8_Bit_t_1n_inst0(.CLK(CLK), .addr(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O), .data(LUT_Array_8_Bit_t_1n_inst0_data));
SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0(.CE(coreir_const11_inst0_out[0]), .CLK(CLK), .O(SizedCounter_1_cinFalse_coutFalse_incr1_hasCETrue_hasResetFalse_inst0_O));
Term_Bitt Term_Bitt_inst0(.I(valid_up));
coreir_const #(.value(1'h1), .width(1)) coreir_const11_inst0(.out(coreir_const11_inst0_out));
assign O = LUT_Array_8_Bit_t_1n_inst0_data;
assign valid_down = coreir_const11_inst0_out[0];
endmodule

module Add_Atom (input [7:0] I__0/*verilator public*/, input [7:0] I__1/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] coreir_add8_inst0_out;
coreir_add #(.width(8)) coreir_add8_inst0(.in0(I__0), .in1(I__1), .out(coreir_add8_inst0_out));
assign O = coreir_add8_inst0_out;
assign valid_down = valid_up;
endmodule

module Module_0 (input CLK/*verilator public*/, input [7:0] I/*verilator public*/, output [7:0] O/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Add_Atom_inst0_O;
wire Add_Atom_inst0_valid_down;
wire [7:0] Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O;
wire Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O;
wire FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire and_inst0_out;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__0;
wire [7:0] atomTupleCreator_t0Int_t1Int_inst0_O__1;
wire atomTupleCreator_t0Int_t1Int_inst0_valid_down;
Add_Atom Add_Atom_inst0(.I__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .I__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .O(Add_Atom_inst0_O), .valid_down(Add_Atom_inst0_valid_down), .valid_up(atomTupleCreator_t0Int_t1Int_inst0_valid_down));
Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .O(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .valid_down(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .O(FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .valid_down(FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(Const_tInt_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
corebit_and and_inst0(.in0(valid_up), .in1(FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .out(and_inst0_out));
atomTupleCreator_t0Int_t1Int atomTupleCreator_t0Int_t1Int_inst0(.I0(I), .I1(FIFO_tInt_delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O), .O__0(atomTupleCreator_t0Int_t1Int_inst0_O__0), .O__1(atomTupleCreator_t0Int_t1Int_inst0_O__1), .valid_down(atomTupleCreator_t0Int_t1Int_inst0_valid_down), .valid_up(and_inst0_out));
assign O = Add_Atom_inst0_O;
assign valid_down = Add_Atom_inst0_valid_down;
endmodule

module NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ (input CLK/*verilator public*/, input [7:0] I_0/*verilator public*/, input [7:0] I_1/*verilator public*/, input [7:0] I_10/*verilator public*/, input [7:0] I_100/*verilator public*/, input [7:0] I_101/*verilator public*/, input [7:0] I_102/*verilator public*/, input [7:0] I_103/*verilator public*/, input [7:0] I_104/*verilator public*/, input [7:0] I_105/*verilator public*/, input [7:0] I_106/*verilator public*/, input [7:0] I_107/*verilator public*/, input [7:0] I_108/*verilator public*/, input [7:0] I_109/*verilator public*/, input [7:0] I_11/*verilator public*/, input [7:0] I_110/*verilator public*/, input [7:0] I_111/*verilator public*/, input [7:0] I_112/*verilator public*/, input [7:0] I_113/*verilator public*/, input [7:0] I_114/*verilator public*/, input [7:0] I_115/*verilator public*/, input [7:0] I_116/*verilator public*/, input [7:0] I_117/*verilator public*/, input [7:0] I_118/*verilator public*/, input [7:0] I_119/*verilator public*/, input [7:0] I_12/*verilator public*/, input [7:0] I_120/*verilator public*/, input [7:0] I_121/*verilator public*/, input [7:0] I_122/*verilator public*/, input [7:0] I_123/*verilator public*/, input [7:0] I_124/*verilator public*/, input [7:0] I_125/*verilator public*/, input [7:0] I_126/*verilator public*/, input [7:0] I_127/*verilator public*/, input [7:0] I_128/*verilator public*/, input [7:0] I_129/*verilator public*/, input [7:0] I_13/*verilator public*/, input [7:0] I_130/*verilator public*/, input [7:0] I_131/*verilator public*/, input [7:0] I_132/*verilator public*/, input [7:0] I_133/*verilator public*/, input [7:0] I_134/*verilator public*/, input [7:0] I_135/*verilator public*/, input [7:0] I_136/*verilator public*/, input [7:0] I_137/*verilator public*/, input [7:0] I_138/*verilator public*/, input [7:0] I_139/*verilator public*/, input [7:0] I_14/*verilator public*/, input [7:0] I_140/*verilator public*/, input [7:0] I_141/*verilator public*/, input [7:0] I_142/*verilator public*/, input [7:0] I_143/*verilator public*/, input [7:0] I_144/*verilator public*/, input [7:0] I_145/*verilator public*/, input [7:0] I_146/*verilator public*/, input [7:0] I_147/*verilator public*/, input [7:0] I_148/*verilator public*/, input [7:0] I_149/*verilator public*/, input [7:0] I_15/*verilator public*/, input [7:0] I_150/*verilator public*/, input [7:0] I_151/*verilator public*/, input [7:0] I_152/*verilator public*/, input [7:0] I_153/*verilator public*/, input [7:0] I_154/*verilator public*/, input [7:0] I_155/*verilator public*/, input [7:0] I_156/*verilator public*/, input [7:0] I_157/*verilator public*/, input [7:0] I_158/*verilator public*/, input [7:0] I_159/*verilator public*/, input [7:0] I_16/*verilator public*/, input [7:0] I_160/*verilator public*/, input [7:0] I_161/*verilator public*/, input [7:0] I_162/*verilator public*/, input [7:0] I_163/*verilator public*/, input [7:0] I_164/*verilator public*/, input [7:0] I_165/*verilator public*/, input [7:0] I_166/*verilator public*/, input [7:0] I_167/*verilator public*/, input [7:0] I_168/*verilator public*/, input [7:0] I_169/*verilator public*/, input [7:0] I_17/*verilator public*/, input [7:0] I_170/*verilator public*/, input [7:0] I_171/*verilator public*/, input [7:0] I_172/*verilator public*/, input [7:0] I_173/*verilator public*/, input [7:0] I_174/*verilator public*/, input [7:0] I_175/*verilator public*/, input [7:0] I_176/*verilator public*/, input [7:0] I_177/*verilator public*/, input [7:0] I_178/*verilator public*/, input [7:0] I_179/*verilator public*/, input [7:0] I_18/*verilator public*/, input [7:0] I_180/*verilator public*/, input [7:0] I_181/*verilator public*/, input [7:0] I_182/*verilator public*/, input [7:0] I_183/*verilator public*/, input [7:0] I_184/*verilator public*/, input [7:0] I_185/*verilator public*/, input [7:0] I_186/*verilator public*/, input [7:0] I_187/*verilator public*/, input [7:0] I_188/*verilator public*/, input [7:0] I_189/*verilator public*/, input [7:0] I_19/*verilator public*/, input [7:0] I_190/*verilator public*/, input [7:0] I_191/*verilator public*/, input [7:0] I_192/*verilator public*/, input [7:0] I_193/*verilator public*/, input [7:0] I_194/*verilator public*/, input [7:0] I_195/*verilator public*/, input [7:0] I_196/*verilator public*/, input [7:0] I_197/*verilator public*/, input [7:0] I_198/*verilator public*/, input [7:0] I_199/*verilator public*/, input [7:0] I_2/*verilator public*/, input [7:0] I_20/*verilator public*/, input [7:0] I_21/*verilator public*/, input [7:0] I_22/*verilator public*/, input [7:0] I_23/*verilator public*/, input [7:0] I_24/*verilator public*/, input [7:0] I_25/*verilator public*/, input [7:0] I_26/*verilator public*/, input [7:0] I_27/*verilator public*/, input [7:0] I_28/*verilator public*/, input [7:0] I_29/*verilator public*/, input [7:0] I_3/*verilator public*/, input [7:0] I_30/*verilator public*/, input [7:0] I_31/*verilator public*/, input [7:0] I_32/*verilator public*/, input [7:0] I_33/*verilator public*/, input [7:0] I_34/*verilator public*/, input [7:0] I_35/*verilator public*/, input [7:0] I_36/*verilator public*/, input [7:0] I_37/*verilator public*/, input [7:0] I_38/*verilator public*/, input [7:0] I_39/*verilator public*/, input [7:0] I_4/*verilator public*/, input [7:0] I_40/*verilator public*/, input [7:0] I_41/*verilator public*/, input [7:0] I_42/*verilator public*/, input [7:0] I_43/*verilator public*/, input [7:0] I_44/*verilator public*/, input [7:0] I_45/*verilator public*/, input [7:0] I_46/*verilator public*/, input [7:0] I_47/*verilator public*/, input [7:0] I_48/*verilator public*/, input [7:0] I_49/*verilator public*/, input [7:0] I_5/*verilator public*/, input [7:0] I_50/*verilator public*/, input [7:0] I_51/*verilator public*/, input [7:0] I_52/*verilator public*/, input [7:0] I_53/*verilator public*/, input [7:0] I_54/*verilator public*/, input [7:0] I_55/*verilator public*/, input [7:0] I_56/*verilator public*/, input [7:0] I_57/*verilator public*/, input [7:0] I_58/*verilator public*/, input [7:0] I_59/*verilator public*/, input [7:0] I_6/*verilator public*/, input [7:0] I_60/*verilator public*/, input [7:0] I_61/*verilator public*/, input [7:0] I_62/*verilator public*/, input [7:0] I_63/*verilator public*/, input [7:0] I_64/*verilator public*/, input [7:0] I_65/*verilator public*/, input [7:0] I_66/*verilator public*/, input [7:0] I_67/*verilator public*/, input [7:0] I_68/*verilator public*/, input [7:0] I_69/*verilator public*/, input [7:0] I_7/*verilator public*/, input [7:0] I_70/*verilator public*/, input [7:0] I_71/*verilator public*/, input [7:0] I_72/*verilator public*/, input [7:0] I_73/*verilator public*/, input [7:0] I_74/*verilator public*/, input [7:0] I_75/*verilator public*/, input [7:0] I_76/*verilator public*/, input [7:0] I_77/*verilator public*/, input [7:0] I_78/*verilator public*/, input [7:0] I_79/*verilator public*/, input [7:0] I_8/*verilator public*/, input [7:0] I_80/*verilator public*/, input [7:0] I_81/*verilator public*/, input [7:0] I_82/*verilator public*/, input [7:0] I_83/*verilator public*/, input [7:0] I_84/*verilator public*/, input [7:0] I_85/*verilator public*/, input [7:0] I_86/*verilator public*/, input [7:0] I_87/*verilator public*/, input [7:0] I_88/*verilator public*/, input [7:0] I_89/*verilator public*/, input [7:0] I_9/*verilator public*/, input [7:0] I_90/*verilator public*/, input [7:0] I_91/*verilator public*/, input [7:0] I_92/*verilator public*/, input [7:0] I_93/*verilator public*/, input [7:0] I_94/*verilator public*/, input [7:0] I_95/*verilator public*/, input [7:0] I_96/*verilator public*/, input [7:0] I_97/*verilator public*/, input [7:0] I_98/*verilator public*/, input [7:0] I_99/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_100/*verilator public*/, output [7:0] O_101/*verilator public*/, output [7:0] O_102/*verilator public*/, output [7:0] O_103/*verilator public*/, output [7:0] O_104/*verilator public*/, output [7:0] O_105/*verilator public*/, output [7:0] O_106/*verilator public*/, output [7:0] O_107/*verilator public*/, output [7:0] O_108/*verilator public*/, output [7:0] O_109/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_110/*verilator public*/, output [7:0] O_111/*verilator public*/, output [7:0] O_112/*verilator public*/, output [7:0] O_113/*verilator public*/, output [7:0] O_114/*verilator public*/, output [7:0] O_115/*verilator public*/, output [7:0] O_116/*verilator public*/, output [7:0] O_117/*verilator public*/, output [7:0] O_118/*verilator public*/, output [7:0] O_119/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_120/*verilator public*/, output [7:0] O_121/*verilator public*/, output [7:0] O_122/*verilator public*/, output [7:0] O_123/*verilator public*/, output [7:0] O_124/*verilator public*/, output [7:0] O_125/*verilator public*/, output [7:0] O_126/*verilator public*/, output [7:0] O_127/*verilator public*/, output [7:0] O_128/*verilator public*/, output [7:0] O_129/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_130/*verilator public*/, output [7:0] O_131/*verilator public*/, output [7:0] O_132/*verilator public*/, output [7:0] O_133/*verilator public*/, output [7:0] O_134/*verilator public*/, output [7:0] O_135/*verilator public*/, output [7:0] O_136/*verilator public*/, output [7:0] O_137/*verilator public*/, output [7:0] O_138/*verilator public*/, output [7:0] O_139/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_140/*verilator public*/, output [7:0] O_141/*verilator public*/, output [7:0] O_142/*verilator public*/, output [7:0] O_143/*verilator public*/, output [7:0] O_144/*verilator public*/, output [7:0] O_145/*verilator public*/, output [7:0] O_146/*verilator public*/, output [7:0] O_147/*verilator public*/, output [7:0] O_148/*verilator public*/, output [7:0] O_149/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_150/*verilator public*/, output [7:0] O_151/*verilator public*/, output [7:0] O_152/*verilator public*/, output [7:0] O_153/*verilator public*/, output [7:0] O_154/*verilator public*/, output [7:0] O_155/*verilator public*/, output [7:0] O_156/*verilator public*/, output [7:0] O_157/*verilator public*/, output [7:0] O_158/*verilator public*/, output [7:0] O_159/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_160/*verilator public*/, output [7:0] O_161/*verilator public*/, output [7:0] O_162/*verilator public*/, output [7:0] O_163/*verilator public*/, output [7:0] O_164/*verilator public*/, output [7:0] O_165/*verilator public*/, output [7:0] O_166/*verilator public*/, output [7:0] O_167/*verilator public*/, output [7:0] O_168/*verilator public*/, output [7:0] O_169/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_170/*verilator public*/, output [7:0] O_171/*verilator public*/, output [7:0] O_172/*verilator public*/, output [7:0] O_173/*verilator public*/, output [7:0] O_174/*verilator public*/, output [7:0] O_175/*verilator public*/, output [7:0] O_176/*verilator public*/, output [7:0] O_177/*verilator public*/, output [7:0] O_178/*verilator public*/, output [7:0] O_179/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_180/*verilator public*/, output [7:0] O_181/*verilator public*/, output [7:0] O_182/*verilator public*/, output [7:0] O_183/*verilator public*/, output [7:0] O_184/*verilator public*/, output [7:0] O_185/*verilator public*/, output [7:0] O_186/*verilator public*/, output [7:0] O_187/*verilator public*/, output [7:0] O_188/*verilator public*/, output [7:0] O_189/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_190/*verilator public*/, output [7:0] O_191/*verilator public*/, output [7:0] O_192/*verilator public*/, output [7:0] O_193/*verilator public*/, output [7:0] O_194/*verilator public*/, output [7:0] O_195/*verilator public*/, output [7:0] O_196/*verilator public*/, output [7:0] O_197/*verilator public*/, output [7:0] O_198/*verilator public*/, output [7:0] O_199/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_40/*verilator public*/, output [7:0] O_41/*verilator public*/, output [7:0] O_42/*verilator public*/, output [7:0] O_43/*verilator public*/, output [7:0] O_44/*verilator public*/, output [7:0] O_45/*verilator public*/, output [7:0] O_46/*verilator public*/, output [7:0] O_47/*verilator public*/, output [7:0] O_48/*verilator public*/, output [7:0] O_49/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_50/*verilator public*/, output [7:0] O_51/*verilator public*/, output [7:0] O_52/*verilator public*/, output [7:0] O_53/*verilator public*/, output [7:0] O_54/*verilator public*/, output [7:0] O_55/*verilator public*/, output [7:0] O_56/*verilator public*/, output [7:0] O_57/*verilator public*/, output [7:0] O_58/*verilator public*/, output [7:0] O_59/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_60/*verilator public*/, output [7:0] O_61/*verilator public*/, output [7:0] O_62/*verilator public*/, output [7:0] O_63/*verilator public*/, output [7:0] O_64/*verilator public*/, output [7:0] O_65/*verilator public*/, output [7:0] O_66/*verilator public*/, output [7:0] O_67/*verilator public*/, output [7:0] O_68/*verilator public*/, output [7:0] O_69/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_70/*verilator public*/, output [7:0] O_71/*verilator public*/, output [7:0] O_72/*verilator public*/, output [7:0] O_73/*verilator public*/, output [7:0] O_74/*verilator public*/, output [7:0] O_75/*verilator public*/, output [7:0] O_76/*verilator public*/, output [7:0] O_77/*verilator public*/, output [7:0] O_78/*verilator public*/, output [7:0] O_79/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_80/*verilator public*/, output [7:0] O_81/*verilator public*/, output [7:0] O_82/*verilator public*/, output [7:0] O_83/*verilator public*/, output [7:0] O_84/*verilator public*/, output [7:0] O_85/*verilator public*/, output [7:0] O_86/*verilator public*/, output [7:0] O_87/*verilator public*/, output [7:0] O_88/*verilator public*/, output [7:0] O_89/*verilator public*/, output [7:0] O_9/*verilator public*/, output [7:0] O_90/*verilator public*/, output [7:0] O_91/*verilator public*/, output [7:0] O_92/*verilator public*/, output [7:0] O_93/*verilator public*/, output [7:0] O_94/*verilator public*/, output [7:0] O_95/*verilator public*/, output [7:0] O_96/*verilator public*/, output [7:0] O_97/*verilator public*/, output [7:0] O_98/*verilator public*/, output [7:0] O_99/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] Module_0_inst0_O;
wire Module_0_inst0_valid_down;
wire [7:0] Module_0_inst1_O;
wire Module_0_inst1_valid_down;
wire [7:0] Module_0_inst10_O;
wire Module_0_inst10_valid_down;
wire [7:0] Module_0_inst100_O;
wire Module_0_inst100_valid_down;
wire [7:0] Module_0_inst101_O;
wire Module_0_inst101_valid_down;
wire [7:0] Module_0_inst102_O;
wire Module_0_inst102_valid_down;
wire [7:0] Module_0_inst103_O;
wire Module_0_inst103_valid_down;
wire [7:0] Module_0_inst104_O;
wire Module_0_inst104_valid_down;
wire [7:0] Module_0_inst105_O;
wire Module_0_inst105_valid_down;
wire [7:0] Module_0_inst106_O;
wire Module_0_inst106_valid_down;
wire [7:0] Module_0_inst107_O;
wire Module_0_inst107_valid_down;
wire [7:0] Module_0_inst108_O;
wire Module_0_inst108_valid_down;
wire [7:0] Module_0_inst109_O;
wire Module_0_inst109_valid_down;
wire [7:0] Module_0_inst11_O;
wire Module_0_inst11_valid_down;
wire [7:0] Module_0_inst110_O;
wire Module_0_inst110_valid_down;
wire [7:0] Module_0_inst111_O;
wire Module_0_inst111_valid_down;
wire [7:0] Module_0_inst112_O;
wire Module_0_inst112_valid_down;
wire [7:0] Module_0_inst113_O;
wire Module_0_inst113_valid_down;
wire [7:0] Module_0_inst114_O;
wire Module_0_inst114_valid_down;
wire [7:0] Module_0_inst115_O;
wire Module_0_inst115_valid_down;
wire [7:0] Module_0_inst116_O;
wire Module_0_inst116_valid_down;
wire [7:0] Module_0_inst117_O;
wire Module_0_inst117_valid_down;
wire [7:0] Module_0_inst118_O;
wire Module_0_inst118_valid_down;
wire [7:0] Module_0_inst119_O;
wire Module_0_inst119_valid_down;
wire [7:0] Module_0_inst12_O;
wire Module_0_inst12_valid_down;
wire [7:0] Module_0_inst120_O;
wire Module_0_inst120_valid_down;
wire [7:0] Module_0_inst121_O;
wire Module_0_inst121_valid_down;
wire [7:0] Module_0_inst122_O;
wire Module_0_inst122_valid_down;
wire [7:0] Module_0_inst123_O;
wire Module_0_inst123_valid_down;
wire [7:0] Module_0_inst124_O;
wire Module_0_inst124_valid_down;
wire [7:0] Module_0_inst125_O;
wire Module_0_inst125_valid_down;
wire [7:0] Module_0_inst126_O;
wire Module_0_inst126_valid_down;
wire [7:0] Module_0_inst127_O;
wire Module_0_inst127_valid_down;
wire [7:0] Module_0_inst128_O;
wire Module_0_inst128_valid_down;
wire [7:0] Module_0_inst129_O;
wire Module_0_inst129_valid_down;
wire [7:0] Module_0_inst13_O;
wire Module_0_inst13_valid_down;
wire [7:0] Module_0_inst130_O;
wire Module_0_inst130_valid_down;
wire [7:0] Module_0_inst131_O;
wire Module_0_inst131_valid_down;
wire [7:0] Module_0_inst132_O;
wire Module_0_inst132_valid_down;
wire [7:0] Module_0_inst133_O;
wire Module_0_inst133_valid_down;
wire [7:0] Module_0_inst134_O;
wire Module_0_inst134_valid_down;
wire [7:0] Module_0_inst135_O;
wire Module_0_inst135_valid_down;
wire [7:0] Module_0_inst136_O;
wire Module_0_inst136_valid_down;
wire [7:0] Module_0_inst137_O;
wire Module_0_inst137_valid_down;
wire [7:0] Module_0_inst138_O;
wire Module_0_inst138_valid_down;
wire [7:0] Module_0_inst139_O;
wire Module_0_inst139_valid_down;
wire [7:0] Module_0_inst14_O;
wire Module_0_inst14_valid_down;
wire [7:0] Module_0_inst140_O;
wire Module_0_inst140_valid_down;
wire [7:0] Module_0_inst141_O;
wire Module_0_inst141_valid_down;
wire [7:0] Module_0_inst142_O;
wire Module_0_inst142_valid_down;
wire [7:0] Module_0_inst143_O;
wire Module_0_inst143_valid_down;
wire [7:0] Module_0_inst144_O;
wire Module_0_inst144_valid_down;
wire [7:0] Module_0_inst145_O;
wire Module_0_inst145_valid_down;
wire [7:0] Module_0_inst146_O;
wire Module_0_inst146_valid_down;
wire [7:0] Module_0_inst147_O;
wire Module_0_inst147_valid_down;
wire [7:0] Module_0_inst148_O;
wire Module_0_inst148_valid_down;
wire [7:0] Module_0_inst149_O;
wire Module_0_inst149_valid_down;
wire [7:0] Module_0_inst15_O;
wire Module_0_inst15_valid_down;
wire [7:0] Module_0_inst150_O;
wire Module_0_inst150_valid_down;
wire [7:0] Module_0_inst151_O;
wire Module_0_inst151_valid_down;
wire [7:0] Module_0_inst152_O;
wire Module_0_inst152_valid_down;
wire [7:0] Module_0_inst153_O;
wire Module_0_inst153_valid_down;
wire [7:0] Module_0_inst154_O;
wire Module_0_inst154_valid_down;
wire [7:0] Module_0_inst155_O;
wire Module_0_inst155_valid_down;
wire [7:0] Module_0_inst156_O;
wire Module_0_inst156_valid_down;
wire [7:0] Module_0_inst157_O;
wire Module_0_inst157_valid_down;
wire [7:0] Module_0_inst158_O;
wire Module_0_inst158_valid_down;
wire [7:0] Module_0_inst159_O;
wire Module_0_inst159_valid_down;
wire [7:0] Module_0_inst16_O;
wire Module_0_inst16_valid_down;
wire [7:0] Module_0_inst160_O;
wire Module_0_inst160_valid_down;
wire [7:0] Module_0_inst161_O;
wire Module_0_inst161_valid_down;
wire [7:0] Module_0_inst162_O;
wire Module_0_inst162_valid_down;
wire [7:0] Module_0_inst163_O;
wire Module_0_inst163_valid_down;
wire [7:0] Module_0_inst164_O;
wire Module_0_inst164_valid_down;
wire [7:0] Module_0_inst165_O;
wire Module_0_inst165_valid_down;
wire [7:0] Module_0_inst166_O;
wire Module_0_inst166_valid_down;
wire [7:0] Module_0_inst167_O;
wire Module_0_inst167_valid_down;
wire [7:0] Module_0_inst168_O;
wire Module_0_inst168_valid_down;
wire [7:0] Module_0_inst169_O;
wire Module_0_inst169_valid_down;
wire [7:0] Module_0_inst17_O;
wire Module_0_inst17_valid_down;
wire [7:0] Module_0_inst170_O;
wire Module_0_inst170_valid_down;
wire [7:0] Module_0_inst171_O;
wire Module_0_inst171_valid_down;
wire [7:0] Module_0_inst172_O;
wire Module_0_inst172_valid_down;
wire [7:0] Module_0_inst173_O;
wire Module_0_inst173_valid_down;
wire [7:0] Module_0_inst174_O;
wire Module_0_inst174_valid_down;
wire [7:0] Module_0_inst175_O;
wire Module_0_inst175_valid_down;
wire [7:0] Module_0_inst176_O;
wire Module_0_inst176_valid_down;
wire [7:0] Module_0_inst177_O;
wire Module_0_inst177_valid_down;
wire [7:0] Module_0_inst178_O;
wire Module_0_inst178_valid_down;
wire [7:0] Module_0_inst179_O;
wire Module_0_inst179_valid_down;
wire [7:0] Module_0_inst18_O;
wire Module_0_inst18_valid_down;
wire [7:0] Module_0_inst180_O;
wire Module_0_inst180_valid_down;
wire [7:0] Module_0_inst181_O;
wire Module_0_inst181_valid_down;
wire [7:0] Module_0_inst182_O;
wire Module_0_inst182_valid_down;
wire [7:0] Module_0_inst183_O;
wire Module_0_inst183_valid_down;
wire [7:0] Module_0_inst184_O;
wire Module_0_inst184_valid_down;
wire [7:0] Module_0_inst185_O;
wire Module_0_inst185_valid_down;
wire [7:0] Module_0_inst186_O;
wire Module_0_inst186_valid_down;
wire [7:0] Module_0_inst187_O;
wire Module_0_inst187_valid_down;
wire [7:0] Module_0_inst188_O;
wire Module_0_inst188_valid_down;
wire [7:0] Module_0_inst189_O;
wire Module_0_inst189_valid_down;
wire [7:0] Module_0_inst19_O;
wire Module_0_inst19_valid_down;
wire [7:0] Module_0_inst190_O;
wire Module_0_inst190_valid_down;
wire [7:0] Module_0_inst191_O;
wire Module_0_inst191_valid_down;
wire [7:0] Module_0_inst192_O;
wire Module_0_inst192_valid_down;
wire [7:0] Module_0_inst193_O;
wire Module_0_inst193_valid_down;
wire [7:0] Module_0_inst194_O;
wire Module_0_inst194_valid_down;
wire [7:0] Module_0_inst195_O;
wire Module_0_inst195_valid_down;
wire [7:0] Module_0_inst196_O;
wire Module_0_inst196_valid_down;
wire [7:0] Module_0_inst197_O;
wire Module_0_inst197_valid_down;
wire [7:0] Module_0_inst198_O;
wire Module_0_inst198_valid_down;
wire [7:0] Module_0_inst199_O;
wire Module_0_inst199_valid_down;
wire [7:0] Module_0_inst2_O;
wire Module_0_inst2_valid_down;
wire [7:0] Module_0_inst20_O;
wire Module_0_inst20_valid_down;
wire [7:0] Module_0_inst21_O;
wire Module_0_inst21_valid_down;
wire [7:0] Module_0_inst22_O;
wire Module_0_inst22_valid_down;
wire [7:0] Module_0_inst23_O;
wire Module_0_inst23_valid_down;
wire [7:0] Module_0_inst24_O;
wire Module_0_inst24_valid_down;
wire [7:0] Module_0_inst25_O;
wire Module_0_inst25_valid_down;
wire [7:0] Module_0_inst26_O;
wire Module_0_inst26_valid_down;
wire [7:0] Module_0_inst27_O;
wire Module_0_inst27_valid_down;
wire [7:0] Module_0_inst28_O;
wire Module_0_inst28_valid_down;
wire [7:0] Module_0_inst29_O;
wire Module_0_inst29_valid_down;
wire [7:0] Module_0_inst3_O;
wire Module_0_inst3_valid_down;
wire [7:0] Module_0_inst30_O;
wire Module_0_inst30_valid_down;
wire [7:0] Module_0_inst31_O;
wire Module_0_inst31_valid_down;
wire [7:0] Module_0_inst32_O;
wire Module_0_inst32_valid_down;
wire [7:0] Module_0_inst33_O;
wire Module_0_inst33_valid_down;
wire [7:0] Module_0_inst34_O;
wire Module_0_inst34_valid_down;
wire [7:0] Module_0_inst35_O;
wire Module_0_inst35_valid_down;
wire [7:0] Module_0_inst36_O;
wire Module_0_inst36_valid_down;
wire [7:0] Module_0_inst37_O;
wire Module_0_inst37_valid_down;
wire [7:0] Module_0_inst38_O;
wire Module_0_inst38_valid_down;
wire [7:0] Module_0_inst39_O;
wire Module_0_inst39_valid_down;
wire [7:0] Module_0_inst4_O;
wire Module_0_inst4_valid_down;
wire [7:0] Module_0_inst40_O;
wire Module_0_inst40_valid_down;
wire [7:0] Module_0_inst41_O;
wire Module_0_inst41_valid_down;
wire [7:0] Module_0_inst42_O;
wire Module_0_inst42_valid_down;
wire [7:0] Module_0_inst43_O;
wire Module_0_inst43_valid_down;
wire [7:0] Module_0_inst44_O;
wire Module_0_inst44_valid_down;
wire [7:0] Module_0_inst45_O;
wire Module_0_inst45_valid_down;
wire [7:0] Module_0_inst46_O;
wire Module_0_inst46_valid_down;
wire [7:0] Module_0_inst47_O;
wire Module_0_inst47_valid_down;
wire [7:0] Module_0_inst48_O;
wire Module_0_inst48_valid_down;
wire [7:0] Module_0_inst49_O;
wire Module_0_inst49_valid_down;
wire [7:0] Module_0_inst5_O;
wire Module_0_inst5_valid_down;
wire [7:0] Module_0_inst50_O;
wire Module_0_inst50_valid_down;
wire [7:0] Module_0_inst51_O;
wire Module_0_inst51_valid_down;
wire [7:0] Module_0_inst52_O;
wire Module_0_inst52_valid_down;
wire [7:0] Module_0_inst53_O;
wire Module_0_inst53_valid_down;
wire [7:0] Module_0_inst54_O;
wire Module_0_inst54_valid_down;
wire [7:0] Module_0_inst55_O;
wire Module_0_inst55_valid_down;
wire [7:0] Module_0_inst56_O;
wire Module_0_inst56_valid_down;
wire [7:0] Module_0_inst57_O;
wire Module_0_inst57_valid_down;
wire [7:0] Module_0_inst58_O;
wire Module_0_inst58_valid_down;
wire [7:0] Module_0_inst59_O;
wire Module_0_inst59_valid_down;
wire [7:0] Module_0_inst6_O;
wire Module_0_inst6_valid_down;
wire [7:0] Module_0_inst60_O;
wire Module_0_inst60_valid_down;
wire [7:0] Module_0_inst61_O;
wire Module_0_inst61_valid_down;
wire [7:0] Module_0_inst62_O;
wire Module_0_inst62_valid_down;
wire [7:0] Module_0_inst63_O;
wire Module_0_inst63_valid_down;
wire [7:0] Module_0_inst64_O;
wire Module_0_inst64_valid_down;
wire [7:0] Module_0_inst65_O;
wire Module_0_inst65_valid_down;
wire [7:0] Module_0_inst66_O;
wire Module_0_inst66_valid_down;
wire [7:0] Module_0_inst67_O;
wire Module_0_inst67_valid_down;
wire [7:0] Module_0_inst68_O;
wire Module_0_inst68_valid_down;
wire [7:0] Module_0_inst69_O;
wire Module_0_inst69_valid_down;
wire [7:0] Module_0_inst7_O;
wire Module_0_inst7_valid_down;
wire [7:0] Module_0_inst70_O;
wire Module_0_inst70_valid_down;
wire [7:0] Module_0_inst71_O;
wire Module_0_inst71_valid_down;
wire [7:0] Module_0_inst72_O;
wire Module_0_inst72_valid_down;
wire [7:0] Module_0_inst73_O;
wire Module_0_inst73_valid_down;
wire [7:0] Module_0_inst74_O;
wire Module_0_inst74_valid_down;
wire [7:0] Module_0_inst75_O;
wire Module_0_inst75_valid_down;
wire [7:0] Module_0_inst76_O;
wire Module_0_inst76_valid_down;
wire [7:0] Module_0_inst77_O;
wire Module_0_inst77_valid_down;
wire [7:0] Module_0_inst78_O;
wire Module_0_inst78_valid_down;
wire [7:0] Module_0_inst79_O;
wire Module_0_inst79_valid_down;
wire [7:0] Module_0_inst8_O;
wire Module_0_inst8_valid_down;
wire [7:0] Module_0_inst80_O;
wire Module_0_inst80_valid_down;
wire [7:0] Module_0_inst81_O;
wire Module_0_inst81_valid_down;
wire [7:0] Module_0_inst82_O;
wire Module_0_inst82_valid_down;
wire [7:0] Module_0_inst83_O;
wire Module_0_inst83_valid_down;
wire [7:0] Module_0_inst84_O;
wire Module_0_inst84_valid_down;
wire [7:0] Module_0_inst85_O;
wire Module_0_inst85_valid_down;
wire [7:0] Module_0_inst86_O;
wire Module_0_inst86_valid_down;
wire [7:0] Module_0_inst87_O;
wire Module_0_inst87_valid_down;
wire [7:0] Module_0_inst88_O;
wire Module_0_inst88_valid_down;
wire [7:0] Module_0_inst89_O;
wire Module_0_inst89_valid_down;
wire [7:0] Module_0_inst9_O;
wire Module_0_inst9_valid_down;
wire [7:0] Module_0_inst90_O;
wire Module_0_inst90_valid_down;
wire [7:0] Module_0_inst91_O;
wire Module_0_inst91_valid_down;
wire [7:0] Module_0_inst92_O;
wire Module_0_inst92_valid_down;
wire [7:0] Module_0_inst93_O;
wire Module_0_inst93_valid_down;
wire [7:0] Module_0_inst94_O;
wire Module_0_inst94_valid_down;
wire [7:0] Module_0_inst95_O;
wire Module_0_inst95_valid_down;
wire [7:0] Module_0_inst96_O;
wire Module_0_inst96_valid_down;
wire [7:0] Module_0_inst97_O;
wire Module_0_inst97_valid_down;
wire [7:0] Module_0_inst98_O;
wire Module_0_inst98_valid_down;
wire [7:0] Module_0_inst99_O;
wire Module_0_inst99_valid_down;
wire and_inst0_out;
wire and_inst1_out;
wire and_inst10_out;
wire and_inst100_out;
wire and_inst101_out;
wire and_inst102_out;
wire and_inst103_out;
wire and_inst104_out;
wire and_inst105_out;
wire and_inst106_out;
wire and_inst107_out;
wire and_inst108_out;
wire and_inst109_out;
wire and_inst11_out;
wire and_inst110_out;
wire and_inst111_out;
wire and_inst112_out;
wire and_inst113_out;
wire and_inst114_out;
wire and_inst115_out;
wire and_inst116_out;
wire and_inst117_out;
wire and_inst118_out;
wire and_inst119_out;
wire and_inst12_out;
wire and_inst120_out;
wire and_inst121_out;
wire and_inst122_out;
wire and_inst123_out;
wire and_inst124_out;
wire and_inst125_out;
wire and_inst126_out;
wire and_inst127_out;
wire and_inst128_out;
wire and_inst129_out;
wire and_inst13_out;
wire and_inst130_out;
wire and_inst131_out;
wire and_inst132_out;
wire and_inst133_out;
wire and_inst134_out;
wire and_inst135_out;
wire and_inst136_out;
wire and_inst137_out;
wire and_inst138_out;
wire and_inst139_out;
wire and_inst14_out;
wire and_inst140_out;
wire and_inst141_out;
wire and_inst142_out;
wire and_inst143_out;
wire and_inst144_out;
wire and_inst145_out;
wire and_inst146_out;
wire and_inst147_out;
wire and_inst148_out;
wire and_inst149_out;
wire and_inst15_out;
wire and_inst150_out;
wire and_inst151_out;
wire and_inst152_out;
wire and_inst153_out;
wire and_inst154_out;
wire and_inst155_out;
wire and_inst156_out;
wire and_inst157_out;
wire and_inst158_out;
wire and_inst159_out;
wire and_inst16_out;
wire and_inst160_out;
wire and_inst161_out;
wire and_inst162_out;
wire and_inst163_out;
wire and_inst164_out;
wire and_inst165_out;
wire and_inst166_out;
wire and_inst167_out;
wire and_inst168_out;
wire and_inst169_out;
wire and_inst17_out;
wire and_inst170_out;
wire and_inst171_out;
wire and_inst172_out;
wire and_inst173_out;
wire and_inst174_out;
wire and_inst175_out;
wire and_inst176_out;
wire and_inst177_out;
wire and_inst178_out;
wire and_inst179_out;
wire and_inst18_out;
wire and_inst180_out;
wire and_inst181_out;
wire and_inst182_out;
wire and_inst183_out;
wire and_inst184_out;
wire and_inst185_out;
wire and_inst186_out;
wire and_inst187_out;
wire and_inst188_out;
wire and_inst189_out;
wire and_inst19_out;
wire and_inst190_out;
wire and_inst191_out;
wire and_inst192_out;
wire and_inst193_out;
wire and_inst194_out;
wire and_inst195_out;
wire and_inst196_out;
wire and_inst197_out;
wire and_inst198_out;
wire and_inst2_out;
wire and_inst20_out;
wire and_inst21_out;
wire and_inst22_out;
wire and_inst23_out;
wire and_inst24_out;
wire and_inst25_out;
wire and_inst26_out;
wire and_inst27_out;
wire and_inst28_out;
wire and_inst29_out;
wire and_inst3_out;
wire and_inst30_out;
wire and_inst31_out;
wire and_inst32_out;
wire and_inst33_out;
wire and_inst34_out;
wire and_inst35_out;
wire and_inst36_out;
wire and_inst37_out;
wire and_inst38_out;
wire and_inst39_out;
wire and_inst4_out;
wire and_inst40_out;
wire and_inst41_out;
wire and_inst42_out;
wire and_inst43_out;
wire and_inst44_out;
wire and_inst45_out;
wire and_inst46_out;
wire and_inst47_out;
wire and_inst48_out;
wire and_inst49_out;
wire and_inst5_out;
wire and_inst50_out;
wire and_inst51_out;
wire and_inst52_out;
wire and_inst53_out;
wire and_inst54_out;
wire and_inst55_out;
wire and_inst56_out;
wire and_inst57_out;
wire and_inst58_out;
wire and_inst59_out;
wire and_inst6_out;
wire and_inst60_out;
wire and_inst61_out;
wire and_inst62_out;
wire and_inst63_out;
wire and_inst64_out;
wire and_inst65_out;
wire and_inst66_out;
wire and_inst67_out;
wire and_inst68_out;
wire and_inst69_out;
wire and_inst7_out;
wire and_inst70_out;
wire and_inst71_out;
wire and_inst72_out;
wire and_inst73_out;
wire and_inst74_out;
wire and_inst75_out;
wire and_inst76_out;
wire and_inst77_out;
wire and_inst78_out;
wire and_inst79_out;
wire and_inst8_out;
wire and_inst80_out;
wire and_inst81_out;
wire and_inst82_out;
wire and_inst83_out;
wire and_inst84_out;
wire and_inst85_out;
wire and_inst86_out;
wire and_inst87_out;
wire and_inst88_out;
wire and_inst89_out;
wire and_inst9_out;
wire and_inst90_out;
wire and_inst91_out;
wire and_inst92_out;
wire and_inst93_out;
wire and_inst94_out;
wire and_inst95_out;
wire and_inst96_out;
wire and_inst97_out;
wire and_inst98_out;
wire and_inst99_out;
Module_0 Module_0_inst0(.CLK(CLK), .I(I_0), .O(Module_0_inst0_O), .valid_down(Module_0_inst0_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst1(.CLK(CLK), .I(I_1), .O(Module_0_inst1_O), .valid_down(Module_0_inst1_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst10(.CLK(CLK), .I(I_10), .O(Module_0_inst10_O), .valid_down(Module_0_inst10_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst100(.CLK(CLK), .I(I_100), .O(Module_0_inst100_O), .valid_down(Module_0_inst100_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst101(.CLK(CLK), .I(I_101), .O(Module_0_inst101_O), .valid_down(Module_0_inst101_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst102(.CLK(CLK), .I(I_102), .O(Module_0_inst102_O), .valid_down(Module_0_inst102_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst103(.CLK(CLK), .I(I_103), .O(Module_0_inst103_O), .valid_down(Module_0_inst103_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst104(.CLK(CLK), .I(I_104), .O(Module_0_inst104_O), .valid_down(Module_0_inst104_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst105(.CLK(CLK), .I(I_105), .O(Module_0_inst105_O), .valid_down(Module_0_inst105_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst106(.CLK(CLK), .I(I_106), .O(Module_0_inst106_O), .valid_down(Module_0_inst106_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst107(.CLK(CLK), .I(I_107), .O(Module_0_inst107_O), .valid_down(Module_0_inst107_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst108(.CLK(CLK), .I(I_108), .O(Module_0_inst108_O), .valid_down(Module_0_inst108_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst109(.CLK(CLK), .I(I_109), .O(Module_0_inst109_O), .valid_down(Module_0_inst109_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst11(.CLK(CLK), .I(I_11), .O(Module_0_inst11_O), .valid_down(Module_0_inst11_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst110(.CLK(CLK), .I(I_110), .O(Module_0_inst110_O), .valid_down(Module_0_inst110_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst111(.CLK(CLK), .I(I_111), .O(Module_0_inst111_O), .valid_down(Module_0_inst111_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst112(.CLK(CLK), .I(I_112), .O(Module_0_inst112_O), .valid_down(Module_0_inst112_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst113(.CLK(CLK), .I(I_113), .O(Module_0_inst113_O), .valid_down(Module_0_inst113_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst114(.CLK(CLK), .I(I_114), .O(Module_0_inst114_O), .valid_down(Module_0_inst114_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst115(.CLK(CLK), .I(I_115), .O(Module_0_inst115_O), .valid_down(Module_0_inst115_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst116(.CLK(CLK), .I(I_116), .O(Module_0_inst116_O), .valid_down(Module_0_inst116_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst117(.CLK(CLK), .I(I_117), .O(Module_0_inst117_O), .valid_down(Module_0_inst117_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst118(.CLK(CLK), .I(I_118), .O(Module_0_inst118_O), .valid_down(Module_0_inst118_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst119(.CLK(CLK), .I(I_119), .O(Module_0_inst119_O), .valid_down(Module_0_inst119_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst12(.CLK(CLK), .I(I_12), .O(Module_0_inst12_O), .valid_down(Module_0_inst12_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst120(.CLK(CLK), .I(I_120), .O(Module_0_inst120_O), .valid_down(Module_0_inst120_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst121(.CLK(CLK), .I(I_121), .O(Module_0_inst121_O), .valid_down(Module_0_inst121_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst122(.CLK(CLK), .I(I_122), .O(Module_0_inst122_O), .valid_down(Module_0_inst122_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst123(.CLK(CLK), .I(I_123), .O(Module_0_inst123_O), .valid_down(Module_0_inst123_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst124(.CLK(CLK), .I(I_124), .O(Module_0_inst124_O), .valid_down(Module_0_inst124_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst125(.CLK(CLK), .I(I_125), .O(Module_0_inst125_O), .valid_down(Module_0_inst125_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst126(.CLK(CLK), .I(I_126), .O(Module_0_inst126_O), .valid_down(Module_0_inst126_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst127(.CLK(CLK), .I(I_127), .O(Module_0_inst127_O), .valid_down(Module_0_inst127_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst128(.CLK(CLK), .I(I_128), .O(Module_0_inst128_O), .valid_down(Module_0_inst128_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst129(.CLK(CLK), .I(I_129), .O(Module_0_inst129_O), .valid_down(Module_0_inst129_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst13(.CLK(CLK), .I(I_13), .O(Module_0_inst13_O), .valid_down(Module_0_inst13_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst130(.CLK(CLK), .I(I_130), .O(Module_0_inst130_O), .valid_down(Module_0_inst130_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst131(.CLK(CLK), .I(I_131), .O(Module_0_inst131_O), .valid_down(Module_0_inst131_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst132(.CLK(CLK), .I(I_132), .O(Module_0_inst132_O), .valid_down(Module_0_inst132_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst133(.CLK(CLK), .I(I_133), .O(Module_0_inst133_O), .valid_down(Module_0_inst133_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst134(.CLK(CLK), .I(I_134), .O(Module_0_inst134_O), .valid_down(Module_0_inst134_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst135(.CLK(CLK), .I(I_135), .O(Module_0_inst135_O), .valid_down(Module_0_inst135_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst136(.CLK(CLK), .I(I_136), .O(Module_0_inst136_O), .valid_down(Module_0_inst136_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst137(.CLK(CLK), .I(I_137), .O(Module_0_inst137_O), .valid_down(Module_0_inst137_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst138(.CLK(CLK), .I(I_138), .O(Module_0_inst138_O), .valid_down(Module_0_inst138_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst139(.CLK(CLK), .I(I_139), .O(Module_0_inst139_O), .valid_down(Module_0_inst139_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst14(.CLK(CLK), .I(I_14), .O(Module_0_inst14_O), .valid_down(Module_0_inst14_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst140(.CLK(CLK), .I(I_140), .O(Module_0_inst140_O), .valid_down(Module_0_inst140_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst141(.CLK(CLK), .I(I_141), .O(Module_0_inst141_O), .valid_down(Module_0_inst141_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst142(.CLK(CLK), .I(I_142), .O(Module_0_inst142_O), .valid_down(Module_0_inst142_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst143(.CLK(CLK), .I(I_143), .O(Module_0_inst143_O), .valid_down(Module_0_inst143_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst144(.CLK(CLK), .I(I_144), .O(Module_0_inst144_O), .valid_down(Module_0_inst144_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst145(.CLK(CLK), .I(I_145), .O(Module_0_inst145_O), .valid_down(Module_0_inst145_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst146(.CLK(CLK), .I(I_146), .O(Module_0_inst146_O), .valid_down(Module_0_inst146_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst147(.CLK(CLK), .I(I_147), .O(Module_0_inst147_O), .valid_down(Module_0_inst147_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst148(.CLK(CLK), .I(I_148), .O(Module_0_inst148_O), .valid_down(Module_0_inst148_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst149(.CLK(CLK), .I(I_149), .O(Module_0_inst149_O), .valid_down(Module_0_inst149_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst15(.CLK(CLK), .I(I_15), .O(Module_0_inst15_O), .valid_down(Module_0_inst15_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst150(.CLK(CLK), .I(I_150), .O(Module_0_inst150_O), .valid_down(Module_0_inst150_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst151(.CLK(CLK), .I(I_151), .O(Module_0_inst151_O), .valid_down(Module_0_inst151_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst152(.CLK(CLK), .I(I_152), .O(Module_0_inst152_O), .valid_down(Module_0_inst152_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst153(.CLK(CLK), .I(I_153), .O(Module_0_inst153_O), .valid_down(Module_0_inst153_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst154(.CLK(CLK), .I(I_154), .O(Module_0_inst154_O), .valid_down(Module_0_inst154_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst155(.CLK(CLK), .I(I_155), .O(Module_0_inst155_O), .valid_down(Module_0_inst155_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst156(.CLK(CLK), .I(I_156), .O(Module_0_inst156_O), .valid_down(Module_0_inst156_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst157(.CLK(CLK), .I(I_157), .O(Module_0_inst157_O), .valid_down(Module_0_inst157_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst158(.CLK(CLK), .I(I_158), .O(Module_0_inst158_O), .valid_down(Module_0_inst158_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst159(.CLK(CLK), .I(I_159), .O(Module_0_inst159_O), .valid_down(Module_0_inst159_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst16(.CLK(CLK), .I(I_16), .O(Module_0_inst16_O), .valid_down(Module_0_inst16_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst160(.CLK(CLK), .I(I_160), .O(Module_0_inst160_O), .valid_down(Module_0_inst160_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst161(.CLK(CLK), .I(I_161), .O(Module_0_inst161_O), .valid_down(Module_0_inst161_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst162(.CLK(CLK), .I(I_162), .O(Module_0_inst162_O), .valid_down(Module_0_inst162_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst163(.CLK(CLK), .I(I_163), .O(Module_0_inst163_O), .valid_down(Module_0_inst163_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst164(.CLK(CLK), .I(I_164), .O(Module_0_inst164_O), .valid_down(Module_0_inst164_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst165(.CLK(CLK), .I(I_165), .O(Module_0_inst165_O), .valid_down(Module_0_inst165_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst166(.CLK(CLK), .I(I_166), .O(Module_0_inst166_O), .valid_down(Module_0_inst166_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst167(.CLK(CLK), .I(I_167), .O(Module_0_inst167_O), .valid_down(Module_0_inst167_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst168(.CLK(CLK), .I(I_168), .O(Module_0_inst168_O), .valid_down(Module_0_inst168_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst169(.CLK(CLK), .I(I_169), .O(Module_0_inst169_O), .valid_down(Module_0_inst169_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst17(.CLK(CLK), .I(I_17), .O(Module_0_inst17_O), .valid_down(Module_0_inst17_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst170(.CLK(CLK), .I(I_170), .O(Module_0_inst170_O), .valid_down(Module_0_inst170_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst171(.CLK(CLK), .I(I_171), .O(Module_0_inst171_O), .valid_down(Module_0_inst171_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst172(.CLK(CLK), .I(I_172), .O(Module_0_inst172_O), .valid_down(Module_0_inst172_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst173(.CLK(CLK), .I(I_173), .O(Module_0_inst173_O), .valid_down(Module_0_inst173_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst174(.CLK(CLK), .I(I_174), .O(Module_0_inst174_O), .valid_down(Module_0_inst174_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst175(.CLK(CLK), .I(I_175), .O(Module_0_inst175_O), .valid_down(Module_0_inst175_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst176(.CLK(CLK), .I(I_176), .O(Module_0_inst176_O), .valid_down(Module_0_inst176_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst177(.CLK(CLK), .I(I_177), .O(Module_0_inst177_O), .valid_down(Module_0_inst177_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst178(.CLK(CLK), .I(I_178), .O(Module_0_inst178_O), .valid_down(Module_0_inst178_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst179(.CLK(CLK), .I(I_179), .O(Module_0_inst179_O), .valid_down(Module_0_inst179_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst18(.CLK(CLK), .I(I_18), .O(Module_0_inst18_O), .valid_down(Module_0_inst18_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst180(.CLK(CLK), .I(I_180), .O(Module_0_inst180_O), .valid_down(Module_0_inst180_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst181(.CLK(CLK), .I(I_181), .O(Module_0_inst181_O), .valid_down(Module_0_inst181_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst182(.CLK(CLK), .I(I_182), .O(Module_0_inst182_O), .valid_down(Module_0_inst182_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst183(.CLK(CLK), .I(I_183), .O(Module_0_inst183_O), .valid_down(Module_0_inst183_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst184(.CLK(CLK), .I(I_184), .O(Module_0_inst184_O), .valid_down(Module_0_inst184_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst185(.CLK(CLK), .I(I_185), .O(Module_0_inst185_O), .valid_down(Module_0_inst185_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst186(.CLK(CLK), .I(I_186), .O(Module_0_inst186_O), .valid_down(Module_0_inst186_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst187(.CLK(CLK), .I(I_187), .O(Module_0_inst187_O), .valid_down(Module_0_inst187_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst188(.CLK(CLK), .I(I_188), .O(Module_0_inst188_O), .valid_down(Module_0_inst188_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst189(.CLK(CLK), .I(I_189), .O(Module_0_inst189_O), .valid_down(Module_0_inst189_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst19(.CLK(CLK), .I(I_19), .O(Module_0_inst19_O), .valid_down(Module_0_inst19_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst190(.CLK(CLK), .I(I_190), .O(Module_0_inst190_O), .valid_down(Module_0_inst190_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst191(.CLK(CLK), .I(I_191), .O(Module_0_inst191_O), .valid_down(Module_0_inst191_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst192(.CLK(CLK), .I(I_192), .O(Module_0_inst192_O), .valid_down(Module_0_inst192_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst193(.CLK(CLK), .I(I_193), .O(Module_0_inst193_O), .valid_down(Module_0_inst193_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst194(.CLK(CLK), .I(I_194), .O(Module_0_inst194_O), .valid_down(Module_0_inst194_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst195(.CLK(CLK), .I(I_195), .O(Module_0_inst195_O), .valid_down(Module_0_inst195_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst196(.CLK(CLK), .I(I_196), .O(Module_0_inst196_O), .valid_down(Module_0_inst196_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst197(.CLK(CLK), .I(I_197), .O(Module_0_inst197_O), .valid_down(Module_0_inst197_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst198(.CLK(CLK), .I(I_198), .O(Module_0_inst198_O), .valid_down(Module_0_inst198_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst199(.CLK(CLK), .I(I_199), .O(Module_0_inst199_O), .valid_down(Module_0_inst199_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst2(.CLK(CLK), .I(I_2), .O(Module_0_inst2_O), .valid_down(Module_0_inst2_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst20(.CLK(CLK), .I(I_20), .O(Module_0_inst20_O), .valid_down(Module_0_inst20_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst21(.CLK(CLK), .I(I_21), .O(Module_0_inst21_O), .valid_down(Module_0_inst21_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst22(.CLK(CLK), .I(I_22), .O(Module_0_inst22_O), .valid_down(Module_0_inst22_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst23(.CLK(CLK), .I(I_23), .O(Module_0_inst23_O), .valid_down(Module_0_inst23_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst24(.CLK(CLK), .I(I_24), .O(Module_0_inst24_O), .valid_down(Module_0_inst24_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst25(.CLK(CLK), .I(I_25), .O(Module_0_inst25_O), .valid_down(Module_0_inst25_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst26(.CLK(CLK), .I(I_26), .O(Module_0_inst26_O), .valid_down(Module_0_inst26_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst27(.CLK(CLK), .I(I_27), .O(Module_0_inst27_O), .valid_down(Module_0_inst27_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst28(.CLK(CLK), .I(I_28), .O(Module_0_inst28_O), .valid_down(Module_0_inst28_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst29(.CLK(CLK), .I(I_29), .O(Module_0_inst29_O), .valid_down(Module_0_inst29_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst3(.CLK(CLK), .I(I_3), .O(Module_0_inst3_O), .valid_down(Module_0_inst3_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst30(.CLK(CLK), .I(I_30), .O(Module_0_inst30_O), .valid_down(Module_0_inst30_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst31(.CLK(CLK), .I(I_31), .O(Module_0_inst31_O), .valid_down(Module_0_inst31_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst32(.CLK(CLK), .I(I_32), .O(Module_0_inst32_O), .valid_down(Module_0_inst32_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst33(.CLK(CLK), .I(I_33), .O(Module_0_inst33_O), .valid_down(Module_0_inst33_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst34(.CLK(CLK), .I(I_34), .O(Module_0_inst34_O), .valid_down(Module_0_inst34_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst35(.CLK(CLK), .I(I_35), .O(Module_0_inst35_O), .valid_down(Module_0_inst35_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst36(.CLK(CLK), .I(I_36), .O(Module_0_inst36_O), .valid_down(Module_0_inst36_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst37(.CLK(CLK), .I(I_37), .O(Module_0_inst37_O), .valid_down(Module_0_inst37_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst38(.CLK(CLK), .I(I_38), .O(Module_0_inst38_O), .valid_down(Module_0_inst38_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst39(.CLK(CLK), .I(I_39), .O(Module_0_inst39_O), .valid_down(Module_0_inst39_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst4(.CLK(CLK), .I(I_4), .O(Module_0_inst4_O), .valid_down(Module_0_inst4_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst40(.CLK(CLK), .I(I_40), .O(Module_0_inst40_O), .valid_down(Module_0_inst40_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst41(.CLK(CLK), .I(I_41), .O(Module_0_inst41_O), .valid_down(Module_0_inst41_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst42(.CLK(CLK), .I(I_42), .O(Module_0_inst42_O), .valid_down(Module_0_inst42_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst43(.CLK(CLK), .I(I_43), .O(Module_0_inst43_O), .valid_down(Module_0_inst43_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst44(.CLK(CLK), .I(I_44), .O(Module_0_inst44_O), .valid_down(Module_0_inst44_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst45(.CLK(CLK), .I(I_45), .O(Module_0_inst45_O), .valid_down(Module_0_inst45_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst46(.CLK(CLK), .I(I_46), .O(Module_0_inst46_O), .valid_down(Module_0_inst46_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst47(.CLK(CLK), .I(I_47), .O(Module_0_inst47_O), .valid_down(Module_0_inst47_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst48(.CLK(CLK), .I(I_48), .O(Module_0_inst48_O), .valid_down(Module_0_inst48_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst49(.CLK(CLK), .I(I_49), .O(Module_0_inst49_O), .valid_down(Module_0_inst49_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst5(.CLK(CLK), .I(I_5), .O(Module_0_inst5_O), .valid_down(Module_0_inst5_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst50(.CLK(CLK), .I(I_50), .O(Module_0_inst50_O), .valid_down(Module_0_inst50_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst51(.CLK(CLK), .I(I_51), .O(Module_0_inst51_O), .valid_down(Module_0_inst51_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst52(.CLK(CLK), .I(I_52), .O(Module_0_inst52_O), .valid_down(Module_0_inst52_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst53(.CLK(CLK), .I(I_53), .O(Module_0_inst53_O), .valid_down(Module_0_inst53_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst54(.CLK(CLK), .I(I_54), .O(Module_0_inst54_O), .valid_down(Module_0_inst54_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst55(.CLK(CLK), .I(I_55), .O(Module_0_inst55_O), .valid_down(Module_0_inst55_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst56(.CLK(CLK), .I(I_56), .O(Module_0_inst56_O), .valid_down(Module_0_inst56_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst57(.CLK(CLK), .I(I_57), .O(Module_0_inst57_O), .valid_down(Module_0_inst57_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst58(.CLK(CLK), .I(I_58), .O(Module_0_inst58_O), .valid_down(Module_0_inst58_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst59(.CLK(CLK), .I(I_59), .O(Module_0_inst59_O), .valid_down(Module_0_inst59_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst6(.CLK(CLK), .I(I_6), .O(Module_0_inst6_O), .valid_down(Module_0_inst6_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst60(.CLK(CLK), .I(I_60), .O(Module_0_inst60_O), .valid_down(Module_0_inst60_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst61(.CLK(CLK), .I(I_61), .O(Module_0_inst61_O), .valid_down(Module_0_inst61_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst62(.CLK(CLK), .I(I_62), .O(Module_0_inst62_O), .valid_down(Module_0_inst62_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst63(.CLK(CLK), .I(I_63), .O(Module_0_inst63_O), .valid_down(Module_0_inst63_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst64(.CLK(CLK), .I(I_64), .O(Module_0_inst64_O), .valid_down(Module_0_inst64_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst65(.CLK(CLK), .I(I_65), .O(Module_0_inst65_O), .valid_down(Module_0_inst65_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst66(.CLK(CLK), .I(I_66), .O(Module_0_inst66_O), .valid_down(Module_0_inst66_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst67(.CLK(CLK), .I(I_67), .O(Module_0_inst67_O), .valid_down(Module_0_inst67_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst68(.CLK(CLK), .I(I_68), .O(Module_0_inst68_O), .valid_down(Module_0_inst68_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst69(.CLK(CLK), .I(I_69), .O(Module_0_inst69_O), .valid_down(Module_0_inst69_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst7(.CLK(CLK), .I(I_7), .O(Module_0_inst7_O), .valid_down(Module_0_inst7_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst70(.CLK(CLK), .I(I_70), .O(Module_0_inst70_O), .valid_down(Module_0_inst70_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst71(.CLK(CLK), .I(I_71), .O(Module_0_inst71_O), .valid_down(Module_0_inst71_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst72(.CLK(CLK), .I(I_72), .O(Module_0_inst72_O), .valid_down(Module_0_inst72_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst73(.CLK(CLK), .I(I_73), .O(Module_0_inst73_O), .valid_down(Module_0_inst73_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst74(.CLK(CLK), .I(I_74), .O(Module_0_inst74_O), .valid_down(Module_0_inst74_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst75(.CLK(CLK), .I(I_75), .O(Module_0_inst75_O), .valid_down(Module_0_inst75_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst76(.CLK(CLK), .I(I_76), .O(Module_0_inst76_O), .valid_down(Module_0_inst76_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst77(.CLK(CLK), .I(I_77), .O(Module_0_inst77_O), .valid_down(Module_0_inst77_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst78(.CLK(CLK), .I(I_78), .O(Module_0_inst78_O), .valid_down(Module_0_inst78_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst79(.CLK(CLK), .I(I_79), .O(Module_0_inst79_O), .valid_down(Module_0_inst79_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst8(.CLK(CLK), .I(I_8), .O(Module_0_inst8_O), .valid_down(Module_0_inst8_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst80(.CLK(CLK), .I(I_80), .O(Module_0_inst80_O), .valid_down(Module_0_inst80_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst81(.CLK(CLK), .I(I_81), .O(Module_0_inst81_O), .valid_down(Module_0_inst81_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst82(.CLK(CLK), .I(I_82), .O(Module_0_inst82_O), .valid_down(Module_0_inst82_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst83(.CLK(CLK), .I(I_83), .O(Module_0_inst83_O), .valid_down(Module_0_inst83_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst84(.CLK(CLK), .I(I_84), .O(Module_0_inst84_O), .valid_down(Module_0_inst84_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst85(.CLK(CLK), .I(I_85), .O(Module_0_inst85_O), .valid_down(Module_0_inst85_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst86(.CLK(CLK), .I(I_86), .O(Module_0_inst86_O), .valid_down(Module_0_inst86_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst87(.CLK(CLK), .I(I_87), .O(Module_0_inst87_O), .valid_down(Module_0_inst87_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst88(.CLK(CLK), .I(I_88), .O(Module_0_inst88_O), .valid_down(Module_0_inst88_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst89(.CLK(CLK), .I(I_89), .O(Module_0_inst89_O), .valid_down(Module_0_inst89_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst9(.CLK(CLK), .I(I_9), .O(Module_0_inst9_O), .valid_down(Module_0_inst9_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst90(.CLK(CLK), .I(I_90), .O(Module_0_inst90_O), .valid_down(Module_0_inst90_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst91(.CLK(CLK), .I(I_91), .O(Module_0_inst91_O), .valid_down(Module_0_inst91_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst92(.CLK(CLK), .I(I_92), .O(Module_0_inst92_O), .valid_down(Module_0_inst92_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst93(.CLK(CLK), .I(I_93), .O(Module_0_inst93_O), .valid_down(Module_0_inst93_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst94(.CLK(CLK), .I(I_94), .O(Module_0_inst94_O), .valid_down(Module_0_inst94_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst95(.CLK(CLK), .I(I_95), .O(Module_0_inst95_O), .valid_down(Module_0_inst95_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst96(.CLK(CLK), .I(I_96), .O(Module_0_inst96_O), .valid_down(Module_0_inst96_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst97(.CLK(CLK), .I(I_97), .O(Module_0_inst97_O), .valid_down(Module_0_inst97_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst98(.CLK(CLK), .I(I_98), .O(Module_0_inst98_O), .valid_down(Module_0_inst98_valid_down), .valid_up(valid_up));
Module_0 Module_0_inst99(.CLK(CLK), .I(I_99), .O(Module_0_inst99_O), .valid_down(Module_0_inst99_valid_down), .valid_up(valid_up));
corebit_and and_inst0(.in0(Module_0_inst0_valid_down), .in1(Module_0_inst1_valid_down), .out(and_inst0_out));
corebit_and and_inst1(.in0(and_inst0_out), .in1(Module_0_inst2_valid_down), .out(and_inst1_out));
corebit_and and_inst10(.in0(and_inst9_out), .in1(Module_0_inst11_valid_down), .out(and_inst10_out));
corebit_and and_inst100(.in0(and_inst99_out), .in1(Module_0_inst101_valid_down), .out(and_inst100_out));
corebit_and and_inst101(.in0(and_inst100_out), .in1(Module_0_inst102_valid_down), .out(and_inst101_out));
corebit_and and_inst102(.in0(and_inst101_out), .in1(Module_0_inst103_valid_down), .out(and_inst102_out));
corebit_and and_inst103(.in0(and_inst102_out), .in1(Module_0_inst104_valid_down), .out(and_inst103_out));
corebit_and and_inst104(.in0(and_inst103_out), .in1(Module_0_inst105_valid_down), .out(and_inst104_out));
corebit_and and_inst105(.in0(and_inst104_out), .in1(Module_0_inst106_valid_down), .out(and_inst105_out));
corebit_and and_inst106(.in0(and_inst105_out), .in1(Module_0_inst107_valid_down), .out(and_inst106_out));
corebit_and and_inst107(.in0(and_inst106_out), .in1(Module_0_inst108_valid_down), .out(and_inst107_out));
corebit_and and_inst108(.in0(and_inst107_out), .in1(Module_0_inst109_valid_down), .out(and_inst108_out));
corebit_and and_inst109(.in0(and_inst108_out), .in1(Module_0_inst110_valid_down), .out(and_inst109_out));
corebit_and and_inst11(.in0(and_inst10_out), .in1(Module_0_inst12_valid_down), .out(and_inst11_out));
corebit_and and_inst110(.in0(and_inst109_out), .in1(Module_0_inst111_valid_down), .out(and_inst110_out));
corebit_and and_inst111(.in0(and_inst110_out), .in1(Module_0_inst112_valid_down), .out(and_inst111_out));
corebit_and and_inst112(.in0(and_inst111_out), .in1(Module_0_inst113_valid_down), .out(and_inst112_out));
corebit_and and_inst113(.in0(and_inst112_out), .in1(Module_0_inst114_valid_down), .out(and_inst113_out));
corebit_and and_inst114(.in0(and_inst113_out), .in1(Module_0_inst115_valid_down), .out(and_inst114_out));
corebit_and and_inst115(.in0(and_inst114_out), .in1(Module_0_inst116_valid_down), .out(and_inst115_out));
corebit_and and_inst116(.in0(and_inst115_out), .in1(Module_0_inst117_valid_down), .out(and_inst116_out));
corebit_and and_inst117(.in0(and_inst116_out), .in1(Module_0_inst118_valid_down), .out(and_inst117_out));
corebit_and and_inst118(.in0(and_inst117_out), .in1(Module_0_inst119_valid_down), .out(and_inst118_out));
corebit_and and_inst119(.in0(and_inst118_out), .in1(Module_0_inst120_valid_down), .out(and_inst119_out));
corebit_and and_inst12(.in0(and_inst11_out), .in1(Module_0_inst13_valid_down), .out(and_inst12_out));
corebit_and and_inst120(.in0(and_inst119_out), .in1(Module_0_inst121_valid_down), .out(and_inst120_out));
corebit_and and_inst121(.in0(and_inst120_out), .in1(Module_0_inst122_valid_down), .out(and_inst121_out));
corebit_and and_inst122(.in0(and_inst121_out), .in1(Module_0_inst123_valid_down), .out(and_inst122_out));
corebit_and and_inst123(.in0(and_inst122_out), .in1(Module_0_inst124_valid_down), .out(and_inst123_out));
corebit_and and_inst124(.in0(and_inst123_out), .in1(Module_0_inst125_valid_down), .out(and_inst124_out));
corebit_and and_inst125(.in0(and_inst124_out), .in1(Module_0_inst126_valid_down), .out(and_inst125_out));
corebit_and and_inst126(.in0(and_inst125_out), .in1(Module_0_inst127_valid_down), .out(and_inst126_out));
corebit_and and_inst127(.in0(and_inst126_out), .in1(Module_0_inst128_valid_down), .out(and_inst127_out));
corebit_and and_inst128(.in0(and_inst127_out), .in1(Module_0_inst129_valid_down), .out(and_inst128_out));
corebit_and and_inst129(.in0(and_inst128_out), .in1(Module_0_inst130_valid_down), .out(and_inst129_out));
corebit_and and_inst13(.in0(and_inst12_out), .in1(Module_0_inst14_valid_down), .out(and_inst13_out));
corebit_and and_inst130(.in0(and_inst129_out), .in1(Module_0_inst131_valid_down), .out(and_inst130_out));
corebit_and and_inst131(.in0(and_inst130_out), .in1(Module_0_inst132_valid_down), .out(and_inst131_out));
corebit_and and_inst132(.in0(and_inst131_out), .in1(Module_0_inst133_valid_down), .out(and_inst132_out));
corebit_and and_inst133(.in0(and_inst132_out), .in1(Module_0_inst134_valid_down), .out(and_inst133_out));
corebit_and and_inst134(.in0(and_inst133_out), .in1(Module_0_inst135_valid_down), .out(and_inst134_out));
corebit_and and_inst135(.in0(and_inst134_out), .in1(Module_0_inst136_valid_down), .out(and_inst135_out));
corebit_and and_inst136(.in0(and_inst135_out), .in1(Module_0_inst137_valid_down), .out(and_inst136_out));
corebit_and and_inst137(.in0(and_inst136_out), .in1(Module_0_inst138_valid_down), .out(and_inst137_out));
corebit_and and_inst138(.in0(and_inst137_out), .in1(Module_0_inst139_valid_down), .out(and_inst138_out));
corebit_and and_inst139(.in0(and_inst138_out), .in1(Module_0_inst140_valid_down), .out(and_inst139_out));
corebit_and and_inst14(.in0(and_inst13_out), .in1(Module_0_inst15_valid_down), .out(and_inst14_out));
corebit_and and_inst140(.in0(and_inst139_out), .in1(Module_0_inst141_valid_down), .out(and_inst140_out));
corebit_and and_inst141(.in0(and_inst140_out), .in1(Module_0_inst142_valid_down), .out(and_inst141_out));
corebit_and and_inst142(.in0(and_inst141_out), .in1(Module_0_inst143_valid_down), .out(and_inst142_out));
corebit_and and_inst143(.in0(and_inst142_out), .in1(Module_0_inst144_valid_down), .out(and_inst143_out));
corebit_and and_inst144(.in0(and_inst143_out), .in1(Module_0_inst145_valid_down), .out(and_inst144_out));
corebit_and and_inst145(.in0(and_inst144_out), .in1(Module_0_inst146_valid_down), .out(and_inst145_out));
corebit_and and_inst146(.in0(and_inst145_out), .in1(Module_0_inst147_valid_down), .out(and_inst146_out));
corebit_and and_inst147(.in0(and_inst146_out), .in1(Module_0_inst148_valid_down), .out(and_inst147_out));
corebit_and and_inst148(.in0(and_inst147_out), .in1(Module_0_inst149_valid_down), .out(and_inst148_out));
corebit_and and_inst149(.in0(and_inst148_out), .in1(Module_0_inst150_valid_down), .out(and_inst149_out));
corebit_and and_inst15(.in0(and_inst14_out), .in1(Module_0_inst16_valid_down), .out(and_inst15_out));
corebit_and and_inst150(.in0(and_inst149_out), .in1(Module_0_inst151_valid_down), .out(and_inst150_out));
corebit_and and_inst151(.in0(and_inst150_out), .in1(Module_0_inst152_valid_down), .out(and_inst151_out));
corebit_and and_inst152(.in0(and_inst151_out), .in1(Module_0_inst153_valid_down), .out(and_inst152_out));
corebit_and and_inst153(.in0(and_inst152_out), .in1(Module_0_inst154_valid_down), .out(and_inst153_out));
corebit_and and_inst154(.in0(and_inst153_out), .in1(Module_0_inst155_valid_down), .out(and_inst154_out));
corebit_and and_inst155(.in0(and_inst154_out), .in1(Module_0_inst156_valid_down), .out(and_inst155_out));
corebit_and and_inst156(.in0(and_inst155_out), .in1(Module_0_inst157_valid_down), .out(and_inst156_out));
corebit_and and_inst157(.in0(and_inst156_out), .in1(Module_0_inst158_valid_down), .out(and_inst157_out));
corebit_and and_inst158(.in0(and_inst157_out), .in1(Module_0_inst159_valid_down), .out(and_inst158_out));
corebit_and and_inst159(.in0(and_inst158_out), .in1(Module_0_inst160_valid_down), .out(and_inst159_out));
corebit_and and_inst16(.in0(and_inst15_out), .in1(Module_0_inst17_valid_down), .out(and_inst16_out));
corebit_and and_inst160(.in0(and_inst159_out), .in1(Module_0_inst161_valid_down), .out(and_inst160_out));
corebit_and and_inst161(.in0(and_inst160_out), .in1(Module_0_inst162_valid_down), .out(and_inst161_out));
corebit_and and_inst162(.in0(and_inst161_out), .in1(Module_0_inst163_valid_down), .out(and_inst162_out));
corebit_and and_inst163(.in0(and_inst162_out), .in1(Module_0_inst164_valid_down), .out(and_inst163_out));
corebit_and and_inst164(.in0(and_inst163_out), .in1(Module_0_inst165_valid_down), .out(and_inst164_out));
corebit_and and_inst165(.in0(and_inst164_out), .in1(Module_0_inst166_valid_down), .out(and_inst165_out));
corebit_and and_inst166(.in0(and_inst165_out), .in1(Module_0_inst167_valid_down), .out(and_inst166_out));
corebit_and and_inst167(.in0(and_inst166_out), .in1(Module_0_inst168_valid_down), .out(and_inst167_out));
corebit_and and_inst168(.in0(and_inst167_out), .in1(Module_0_inst169_valid_down), .out(and_inst168_out));
corebit_and and_inst169(.in0(and_inst168_out), .in1(Module_0_inst170_valid_down), .out(and_inst169_out));
corebit_and and_inst17(.in0(and_inst16_out), .in1(Module_0_inst18_valid_down), .out(and_inst17_out));
corebit_and and_inst170(.in0(and_inst169_out), .in1(Module_0_inst171_valid_down), .out(and_inst170_out));
corebit_and and_inst171(.in0(and_inst170_out), .in1(Module_0_inst172_valid_down), .out(and_inst171_out));
corebit_and and_inst172(.in0(and_inst171_out), .in1(Module_0_inst173_valid_down), .out(and_inst172_out));
corebit_and and_inst173(.in0(and_inst172_out), .in1(Module_0_inst174_valid_down), .out(and_inst173_out));
corebit_and and_inst174(.in0(and_inst173_out), .in1(Module_0_inst175_valid_down), .out(and_inst174_out));
corebit_and and_inst175(.in0(and_inst174_out), .in1(Module_0_inst176_valid_down), .out(and_inst175_out));
corebit_and and_inst176(.in0(and_inst175_out), .in1(Module_0_inst177_valid_down), .out(and_inst176_out));
corebit_and and_inst177(.in0(and_inst176_out), .in1(Module_0_inst178_valid_down), .out(and_inst177_out));
corebit_and and_inst178(.in0(and_inst177_out), .in1(Module_0_inst179_valid_down), .out(and_inst178_out));
corebit_and and_inst179(.in0(and_inst178_out), .in1(Module_0_inst180_valid_down), .out(and_inst179_out));
corebit_and and_inst18(.in0(and_inst17_out), .in1(Module_0_inst19_valid_down), .out(and_inst18_out));
corebit_and and_inst180(.in0(and_inst179_out), .in1(Module_0_inst181_valid_down), .out(and_inst180_out));
corebit_and and_inst181(.in0(and_inst180_out), .in1(Module_0_inst182_valid_down), .out(and_inst181_out));
corebit_and and_inst182(.in0(and_inst181_out), .in1(Module_0_inst183_valid_down), .out(and_inst182_out));
corebit_and and_inst183(.in0(and_inst182_out), .in1(Module_0_inst184_valid_down), .out(and_inst183_out));
corebit_and and_inst184(.in0(and_inst183_out), .in1(Module_0_inst185_valid_down), .out(and_inst184_out));
corebit_and and_inst185(.in0(and_inst184_out), .in1(Module_0_inst186_valid_down), .out(and_inst185_out));
corebit_and and_inst186(.in0(and_inst185_out), .in1(Module_0_inst187_valid_down), .out(and_inst186_out));
corebit_and and_inst187(.in0(and_inst186_out), .in1(Module_0_inst188_valid_down), .out(and_inst187_out));
corebit_and and_inst188(.in0(and_inst187_out), .in1(Module_0_inst189_valid_down), .out(and_inst188_out));
corebit_and and_inst189(.in0(and_inst188_out), .in1(Module_0_inst190_valid_down), .out(and_inst189_out));
corebit_and and_inst19(.in0(and_inst18_out), .in1(Module_0_inst20_valid_down), .out(and_inst19_out));
corebit_and and_inst190(.in0(and_inst189_out), .in1(Module_0_inst191_valid_down), .out(and_inst190_out));
corebit_and and_inst191(.in0(and_inst190_out), .in1(Module_0_inst192_valid_down), .out(and_inst191_out));
corebit_and and_inst192(.in0(and_inst191_out), .in1(Module_0_inst193_valid_down), .out(and_inst192_out));
corebit_and and_inst193(.in0(and_inst192_out), .in1(Module_0_inst194_valid_down), .out(and_inst193_out));
corebit_and and_inst194(.in0(and_inst193_out), .in1(Module_0_inst195_valid_down), .out(and_inst194_out));
corebit_and and_inst195(.in0(and_inst194_out), .in1(Module_0_inst196_valid_down), .out(and_inst195_out));
corebit_and and_inst196(.in0(and_inst195_out), .in1(Module_0_inst197_valid_down), .out(and_inst196_out));
corebit_and and_inst197(.in0(and_inst196_out), .in1(Module_0_inst198_valid_down), .out(and_inst197_out));
corebit_and and_inst198(.in0(and_inst197_out), .in1(Module_0_inst199_valid_down), .out(and_inst198_out));
corebit_and and_inst2(.in0(and_inst1_out), .in1(Module_0_inst3_valid_down), .out(and_inst2_out));
corebit_and and_inst20(.in0(and_inst19_out), .in1(Module_0_inst21_valid_down), .out(and_inst20_out));
corebit_and and_inst21(.in0(and_inst20_out), .in1(Module_0_inst22_valid_down), .out(and_inst21_out));
corebit_and and_inst22(.in0(and_inst21_out), .in1(Module_0_inst23_valid_down), .out(and_inst22_out));
corebit_and and_inst23(.in0(and_inst22_out), .in1(Module_0_inst24_valid_down), .out(and_inst23_out));
corebit_and and_inst24(.in0(and_inst23_out), .in1(Module_0_inst25_valid_down), .out(and_inst24_out));
corebit_and and_inst25(.in0(and_inst24_out), .in1(Module_0_inst26_valid_down), .out(and_inst25_out));
corebit_and and_inst26(.in0(and_inst25_out), .in1(Module_0_inst27_valid_down), .out(and_inst26_out));
corebit_and and_inst27(.in0(and_inst26_out), .in1(Module_0_inst28_valid_down), .out(and_inst27_out));
corebit_and and_inst28(.in0(and_inst27_out), .in1(Module_0_inst29_valid_down), .out(and_inst28_out));
corebit_and and_inst29(.in0(and_inst28_out), .in1(Module_0_inst30_valid_down), .out(and_inst29_out));
corebit_and and_inst3(.in0(and_inst2_out), .in1(Module_0_inst4_valid_down), .out(and_inst3_out));
corebit_and and_inst30(.in0(and_inst29_out), .in1(Module_0_inst31_valid_down), .out(and_inst30_out));
corebit_and and_inst31(.in0(and_inst30_out), .in1(Module_0_inst32_valid_down), .out(and_inst31_out));
corebit_and and_inst32(.in0(and_inst31_out), .in1(Module_0_inst33_valid_down), .out(and_inst32_out));
corebit_and and_inst33(.in0(and_inst32_out), .in1(Module_0_inst34_valid_down), .out(and_inst33_out));
corebit_and and_inst34(.in0(and_inst33_out), .in1(Module_0_inst35_valid_down), .out(and_inst34_out));
corebit_and and_inst35(.in0(and_inst34_out), .in1(Module_0_inst36_valid_down), .out(and_inst35_out));
corebit_and and_inst36(.in0(and_inst35_out), .in1(Module_0_inst37_valid_down), .out(and_inst36_out));
corebit_and and_inst37(.in0(and_inst36_out), .in1(Module_0_inst38_valid_down), .out(and_inst37_out));
corebit_and and_inst38(.in0(and_inst37_out), .in1(Module_0_inst39_valid_down), .out(and_inst38_out));
corebit_and and_inst39(.in0(and_inst38_out), .in1(Module_0_inst40_valid_down), .out(and_inst39_out));
corebit_and and_inst4(.in0(and_inst3_out), .in1(Module_0_inst5_valid_down), .out(and_inst4_out));
corebit_and and_inst40(.in0(and_inst39_out), .in1(Module_0_inst41_valid_down), .out(and_inst40_out));
corebit_and and_inst41(.in0(and_inst40_out), .in1(Module_0_inst42_valid_down), .out(and_inst41_out));
corebit_and and_inst42(.in0(and_inst41_out), .in1(Module_0_inst43_valid_down), .out(and_inst42_out));
corebit_and and_inst43(.in0(and_inst42_out), .in1(Module_0_inst44_valid_down), .out(and_inst43_out));
corebit_and and_inst44(.in0(and_inst43_out), .in1(Module_0_inst45_valid_down), .out(and_inst44_out));
corebit_and and_inst45(.in0(and_inst44_out), .in1(Module_0_inst46_valid_down), .out(and_inst45_out));
corebit_and and_inst46(.in0(and_inst45_out), .in1(Module_0_inst47_valid_down), .out(and_inst46_out));
corebit_and and_inst47(.in0(and_inst46_out), .in1(Module_0_inst48_valid_down), .out(and_inst47_out));
corebit_and and_inst48(.in0(and_inst47_out), .in1(Module_0_inst49_valid_down), .out(and_inst48_out));
corebit_and and_inst49(.in0(and_inst48_out), .in1(Module_0_inst50_valid_down), .out(and_inst49_out));
corebit_and and_inst5(.in0(and_inst4_out), .in1(Module_0_inst6_valid_down), .out(and_inst5_out));
corebit_and and_inst50(.in0(and_inst49_out), .in1(Module_0_inst51_valid_down), .out(and_inst50_out));
corebit_and and_inst51(.in0(and_inst50_out), .in1(Module_0_inst52_valid_down), .out(and_inst51_out));
corebit_and and_inst52(.in0(and_inst51_out), .in1(Module_0_inst53_valid_down), .out(and_inst52_out));
corebit_and and_inst53(.in0(and_inst52_out), .in1(Module_0_inst54_valid_down), .out(and_inst53_out));
corebit_and and_inst54(.in0(and_inst53_out), .in1(Module_0_inst55_valid_down), .out(and_inst54_out));
corebit_and and_inst55(.in0(and_inst54_out), .in1(Module_0_inst56_valid_down), .out(and_inst55_out));
corebit_and and_inst56(.in0(and_inst55_out), .in1(Module_0_inst57_valid_down), .out(and_inst56_out));
corebit_and and_inst57(.in0(and_inst56_out), .in1(Module_0_inst58_valid_down), .out(and_inst57_out));
corebit_and and_inst58(.in0(and_inst57_out), .in1(Module_0_inst59_valid_down), .out(and_inst58_out));
corebit_and and_inst59(.in0(and_inst58_out), .in1(Module_0_inst60_valid_down), .out(and_inst59_out));
corebit_and and_inst6(.in0(and_inst5_out), .in1(Module_0_inst7_valid_down), .out(and_inst6_out));
corebit_and and_inst60(.in0(and_inst59_out), .in1(Module_0_inst61_valid_down), .out(and_inst60_out));
corebit_and and_inst61(.in0(and_inst60_out), .in1(Module_0_inst62_valid_down), .out(and_inst61_out));
corebit_and and_inst62(.in0(and_inst61_out), .in1(Module_0_inst63_valid_down), .out(and_inst62_out));
corebit_and and_inst63(.in0(and_inst62_out), .in1(Module_0_inst64_valid_down), .out(and_inst63_out));
corebit_and and_inst64(.in0(and_inst63_out), .in1(Module_0_inst65_valid_down), .out(and_inst64_out));
corebit_and and_inst65(.in0(and_inst64_out), .in1(Module_0_inst66_valid_down), .out(and_inst65_out));
corebit_and and_inst66(.in0(and_inst65_out), .in1(Module_0_inst67_valid_down), .out(and_inst66_out));
corebit_and and_inst67(.in0(and_inst66_out), .in1(Module_0_inst68_valid_down), .out(and_inst67_out));
corebit_and and_inst68(.in0(and_inst67_out), .in1(Module_0_inst69_valid_down), .out(and_inst68_out));
corebit_and and_inst69(.in0(and_inst68_out), .in1(Module_0_inst70_valid_down), .out(and_inst69_out));
corebit_and and_inst7(.in0(and_inst6_out), .in1(Module_0_inst8_valid_down), .out(and_inst7_out));
corebit_and and_inst70(.in0(and_inst69_out), .in1(Module_0_inst71_valid_down), .out(and_inst70_out));
corebit_and and_inst71(.in0(and_inst70_out), .in1(Module_0_inst72_valid_down), .out(and_inst71_out));
corebit_and and_inst72(.in0(and_inst71_out), .in1(Module_0_inst73_valid_down), .out(and_inst72_out));
corebit_and and_inst73(.in0(and_inst72_out), .in1(Module_0_inst74_valid_down), .out(and_inst73_out));
corebit_and and_inst74(.in0(and_inst73_out), .in1(Module_0_inst75_valid_down), .out(and_inst74_out));
corebit_and and_inst75(.in0(and_inst74_out), .in1(Module_0_inst76_valid_down), .out(and_inst75_out));
corebit_and and_inst76(.in0(and_inst75_out), .in1(Module_0_inst77_valid_down), .out(and_inst76_out));
corebit_and and_inst77(.in0(and_inst76_out), .in1(Module_0_inst78_valid_down), .out(and_inst77_out));
corebit_and and_inst78(.in0(and_inst77_out), .in1(Module_0_inst79_valid_down), .out(and_inst78_out));
corebit_and and_inst79(.in0(and_inst78_out), .in1(Module_0_inst80_valid_down), .out(and_inst79_out));
corebit_and and_inst8(.in0(and_inst7_out), .in1(Module_0_inst9_valid_down), .out(and_inst8_out));
corebit_and and_inst80(.in0(and_inst79_out), .in1(Module_0_inst81_valid_down), .out(and_inst80_out));
corebit_and and_inst81(.in0(and_inst80_out), .in1(Module_0_inst82_valid_down), .out(and_inst81_out));
corebit_and and_inst82(.in0(and_inst81_out), .in1(Module_0_inst83_valid_down), .out(and_inst82_out));
corebit_and and_inst83(.in0(and_inst82_out), .in1(Module_0_inst84_valid_down), .out(and_inst83_out));
corebit_and and_inst84(.in0(and_inst83_out), .in1(Module_0_inst85_valid_down), .out(and_inst84_out));
corebit_and and_inst85(.in0(and_inst84_out), .in1(Module_0_inst86_valid_down), .out(and_inst85_out));
corebit_and and_inst86(.in0(and_inst85_out), .in1(Module_0_inst87_valid_down), .out(and_inst86_out));
corebit_and and_inst87(.in0(and_inst86_out), .in1(Module_0_inst88_valid_down), .out(and_inst87_out));
corebit_and and_inst88(.in0(and_inst87_out), .in1(Module_0_inst89_valid_down), .out(and_inst88_out));
corebit_and and_inst89(.in0(and_inst88_out), .in1(Module_0_inst90_valid_down), .out(and_inst89_out));
corebit_and and_inst9(.in0(and_inst8_out), .in1(Module_0_inst10_valid_down), .out(and_inst9_out));
corebit_and and_inst90(.in0(and_inst89_out), .in1(Module_0_inst91_valid_down), .out(and_inst90_out));
corebit_and and_inst91(.in0(and_inst90_out), .in1(Module_0_inst92_valid_down), .out(and_inst91_out));
corebit_and and_inst92(.in0(and_inst91_out), .in1(Module_0_inst93_valid_down), .out(and_inst92_out));
corebit_and and_inst93(.in0(and_inst92_out), .in1(Module_0_inst94_valid_down), .out(and_inst93_out));
corebit_and and_inst94(.in0(and_inst93_out), .in1(Module_0_inst95_valid_down), .out(and_inst94_out));
corebit_and and_inst95(.in0(and_inst94_out), .in1(Module_0_inst96_valid_down), .out(and_inst95_out));
corebit_and and_inst96(.in0(and_inst95_out), .in1(Module_0_inst97_valid_down), .out(and_inst96_out));
corebit_and and_inst97(.in0(and_inst96_out), .in1(Module_0_inst98_valid_down), .out(and_inst97_out));
corebit_and and_inst98(.in0(and_inst97_out), .in1(Module_0_inst99_valid_down), .out(and_inst98_out));
corebit_and and_inst99(.in0(and_inst98_out), .in1(Module_0_inst100_valid_down), .out(and_inst99_out));
assign O_0 = Module_0_inst0_O;
assign O_1 = Module_0_inst1_O;
assign O_10 = Module_0_inst10_O;
assign O_100 = Module_0_inst100_O;
assign O_101 = Module_0_inst101_O;
assign O_102 = Module_0_inst102_O;
assign O_103 = Module_0_inst103_O;
assign O_104 = Module_0_inst104_O;
assign O_105 = Module_0_inst105_O;
assign O_106 = Module_0_inst106_O;
assign O_107 = Module_0_inst107_O;
assign O_108 = Module_0_inst108_O;
assign O_109 = Module_0_inst109_O;
assign O_11 = Module_0_inst11_O;
assign O_110 = Module_0_inst110_O;
assign O_111 = Module_0_inst111_O;
assign O_112 = Module_0_inst112_O;
assign O_113 = Module_0_inst113_O;
assign O_114 = Module_0_inst114_O;
assign O_115 = Module_0_inst115_O;
assign O_116 = Module_0_inst116_O;
assign O_117 = Module_0_inst117_O;
assign O_118 = Module_0_inst118_O;
assign O_119 = Module_0_inst119_O;
assign O_12 = Module_0_inst12_O;
assign O_120 = Module_0_inst120_O;
assign O_121 = Module_0_inst121_O;
assign O_122 = Module_0_inst122_O;
assign O_123 = Module_0_inst123_O;
assign O_124 = Module_0_inst124_O;
assign O_125 = Module_0_inst125_O;
assign O_126 = Module_0_inst126_O;
assign O_127 = Module_0_inst127_O;
assign O_128 = Module_0_inst128_O;
assign O_129 = Module_0_inst129_O;
assign O_13 = Module_0_inst13_O;
assign O_130 = Module_0_inst130_O;
assign O_131 = Module_0_inst131_O;
assign O_132 = Module_0_inst132_O;
assign O_133 = Module_0_inst133_O;
assign O_134 = Module_0_inst134_O;
assign O_135 = Module_0_inst135_O;
assign O_136 = Module_0_inst136_O;
assign O_137 = Module_0_inst137_O;
assign O_138 = Module_0_inst138_O;
assign O_139 = Module_0_inst139_O;
assign O_14 = Module_0_inst14_O;
assign O_140 = Module_0_inst140_O;
assign O_141 = Module_0_inst141_O;
assign O_142 = Module_0_inst142_O;
assign O_143 = Module_0_inst143_O;
assign O_144 = Module_0_inst144_O;
assign O_145 = Module_0_inst145_O;
assign O_146 = Module_0_inst146_O;
assign O_147 = Module_0_inst147_O;
assign O_148 = Module_0_inst148_O;
assign O_149 = Module_0_inst149_O;
assign O_15 = Module_0_inst15_O;
assign O_150 = Module_0_inst150_O;
assign O_151 = Module_0_inst151_O;
assign O_152 = Module_0_inst152_O;
assign O_153 = Module_0_inst153_O;
assign O_154 = Module_0_inst154_O;
assign O_155 = Module_0_inst155_O;
assign O_156 = Module_0_inst156_O;
assign O_157 = Module_0_inst157_O;
assign O_158 = Module_0_inst158_O;
assign O_159 = Module_0_inst159_O;
assign O_16 = Module_0_inst16_O;
assign O_160 = Module_0_inst160_O;
assign O_161 = Module_0_inst161_O;
assign O_162 = Module_0_inst162_O;
assign O_163 = Module_0_inst163_O;
assign O_164 = Module_0_inst164_O;
assign O_165 = Module_0_inst165_O;
assign O_166 = Module_0_inst166_O;
assign O_167 = Module_0_inst167_O;
assign O_168 = Module_0_inst168_O;
assign O_169 = Module_0_inst169_O;
assign O_17 = Module_0_inst17_O;
assign O_170 = Module_0_inst170_O;
assign O_171 = Module_0_inst171_O;
assign O_172 = Module_0_inst172_O;
assign O_173 = Module_0_inst173_O;
assign O_174 = Module_0_inst174_O;
assign O_175 = Module_0_inst175_O;
assign O_176 = Module_0_inst176_O;
assign O_177 = Module_0_inst177_O;
assign O_178 = Module_0_inst178_O;
assign O_179 = Module_0_inst179_O;
assign O_18 = Module_0_inst18_O;
assign O_180 = Module_0_inst180_O;
assign O_181 = Module_0_inst181_O;
assign O_182 = Module_0_inst182_O;
assign O_183 = Module_0_inst183_O;
assign O_184 = Module_0_inst184_O;
assign O_185 = Module_0_inst185_O;
assign O_186 = Module_0_inst186_O;
assign O_187 = Module_0_inst187_O;
assign O_188 = Module_0_inst188_O;
assign O_189 = Module_0_inst189_O;
assign O_19 = Module_0_inst19_O;
assign O_190 = Module_0_inst190_O;
assign O_191 = Module_0_inst191_O;
assign O_192 = Module_0_inst192_O;
assign O_193 = Module_0_inst193_O;
assign O_194 = Module_0_inst194_O;
assign O_195 = Module_0_inst195_O;
assign O_196 = Module_0_inst196_O;
assign O_197 = Module_0_inst197_O;
assign O_198 = Module_0_inst198_O;
assign O_199 = Module_0_inst199_O;
assign O_2 = Module_0_inst2_O;
assign O_20 = Module_0_inst20_O;
assign O_21 = Module_0_inst21_O;
assign O_22 = Module_0_inst22_O;
assign O_23 = Module_0_inst23_O;
assign O_24 = Module_0_inst24_O;
assign O_25 = Module_0_inst25_O;
assign O_26 = Module_0_inst26_O;
assign O_27 = Module_0_inst27_O;
assign O_28 = Module_0_inst28_O;
assign O_29 = Module_0_inst29_O;
assign O_3 = Module_0_inst3_O;
assign O_30 = Module_0_inst30_O;
assign O_31 = Module_0_inst31_O;
assign O_32 = Module_0_inst32_O;
assign O_33 = Module_0_inst33_O;
assign O_34 = Module_0_inst34_O;
assign O_35 = Module_0_inst35_O;
assign O_36 = Module_0_inst36_O;
assign O_37 = Module_0_inst37_O;
assign O_38 = Module_0_inst38_O;
assign O_39 = Module_0_inst39_O;
assign O_4 = Module_0_inst4_O;
assign O_40 = Module_0_inst40_O;
assign O_41 = Module_0_inst41_O;
assign O_42 = Module_0_inst42_O;
assign O_43 = Module_0_inst43_O;
assign O_44 = Module_0_inst44_O;
assign O_45 = Module_0_inst45_O;
assign O_46 = Module_0_inst46_O;
assign O_47 = Module_0_inst47_O;
assign O_48 = Module_0_inst48_O;
assign O_49 = Module_0_inst49_O;
assign O_5 = Module_0_inst5_O;
assign O_50 = Module_0_inst50_O;
assign O_51 = Module_0_inst51_O;
assign O_52 = Module_0_inst52_O;
assign O_53 = Module_0_inst53_O;
assign O_54 = Module_0_inst54_O;
assign O_55 = Module_0_inst55_O;
assign O_56 = Module_0_inst56_O;
assign O_57 = Module_0_inst57_O;
assign O_58 = Module_0_inst58_O;
assign O_59 = Module_0_inst59_O;
assign O_6 = Module_0_inst6_O;
assign O_60 = Module_0_inst60_O;
assign O_61 = Module_0_inst61_O;
assign O_62 = Module_0_inst62_O;
assign O_63 = Module_0_inst63_O;
assign O_64 = Module_0_inst64_O;
assign O_65 = Module_0_inst65_O;
assign O_66 = Module_0_inst66_O;
assign O_67 = Module_0_inst67_O;
assign O_68 = Module_0_inst68_O;
assign O_69 = Module_0_inst69_O;
assign O_7 = Module_0_inst7_O;
assign O_70 = Module_0_inst70_O;
assign O_71 = Module_0_inst71_O;
assign O_72 = Module_0_inst72_O;
assign O_73 = Module_0_inst73_O;
assign O_74 = Module_0_inst74_O;
assign O_75 = Module_0_inst75_O;
assign O_76 = Module_0_inst76_O;
assign O_77 = Module_0_inst77_O;
assign O_78 = Module_0_inst78_O;
assign O_79 = Module_0_inst79_O;
assign O_8 = Module_0_inst8_O;
assign O_80 = Module_0_inst80_O;
assign O_81 = Module_0_inst81_O;
assign O_82 = Module_0_inst82_O;
assign O_83 = Module_0_inst83_O;
assign O_84 = Module_0_inst84_O;
assign O_85 = Module_0_inst85_O;
assign O_86 = Module_0_inst86_O;
assign O_87 = Module_0_inst87_O;
assign O_88 = Module_0_inst88_O;
assign O_89 = Module_0_inst89_O;
assign O_9 = Module_0_inst9_O;
assign O_90 = Module_0_inst90_O;
assign O_91 = Module_0_inst91_O;
assign O_92 = Module_0_inst92_O;
assign O_93 = Module_0_inst93_O;
assign O_94 = Module_0_inst94_O;
assign O_95 = Module_0_inst95_O;
assign O_96 = Module_0_inst96_O;
assign O_97 = Module_0_inst97_O;
assign O_98 = Module_0_inst98_O;
assign O_99 = Module_0_inst99_O;
assign valid_down = and_inst198_out;
endmodule

module top (input CLK/*verilator public*/, output [7:0] O_0/*verilator public*/, output [7:0] O_1/*verilator public*/, output [7:0] O_10/*verilator public*/, output [7:0] O_100/*verilator public*/, output [7:0] O_101/*verilator public*/, output [7:0] O_102/*verilator public*/, output [7:0] O_103/*verilator public*/, output [7:0] O_104/*verilator public*/, output [7:0] O_105/*verilator public*/, output [7:0] O_106/*verilator public*/, output [7:0] O_107/*verilator public*/, output [7:0] O_108/*verilator public*/, output [7:0] O_109/*verilator public*/, output [7:0] O_11/*verilator public*/, output [7:0] O_110/*verilator public*/, output [7:0] O_111/*verilator public*/, output [7:0] O_112/*verilator public*/, output [7:0] O_113/*verilator public*/, output [7:0] O_114/*verilator public*/, output [7:0] O_115/*verilator public*/, output [7:0] O_116/*verilator public*/, output [7:0] O_117/*verilator public*/, output [7:0] O_118/*verilator public*/, output [7:0] O_119/*verilator public*/, output [7:0] O_12/*verilator public*/, output [7:0] O_120/*verilator public*/, output [7:0] O_121/*verilator public*/, output [7:0] O_122/*verilator public*/, output [7:0] O_123/*verilator public*/, output [7:0] O_124/*verilator public*/, output [7:0] O_125/*verilator public*/, output [7:0] O_126/*verilator public*/, output [7:0] O_127/*verilator public*/, output [7:0] O_128/*verilator public*/, output [7:0] O_129/*verilator public*/, output [7:0] O_13/*verilator public*/, output [7:0] O_130/*verilator public*/, output [7:0] O_131/*verilator public*/, output [7:0] O_132/*verilator public*/, output [7:0] O_133/*verilator public*/, output [7:0] O_134/*verilator public*/, output [7:0] O_135/*verilator public*/, output [7:0] O_136/*verilator public*/, output [7:0] O_137/*verilator public*/, output [7:0] O_138/*verilator public*/, output [7:0] O_139/*verilator public*/, output [7:0] O_14/*verilator public*/, output [7:0] O_140/*verilator public*/, output [7:0] O_141/*verilator public*/, output [7:0] O_142/*verilator public*/, output [7:0] O_143/*verilator public*/, output [7:0] O_144/*verilator public*/, output [7:0] O_145/*verilator public*/, output [7:0] O_146/*verilator public*/, output [7:0] O_147/*verilator public*/, output [7:0] O_148/*verilator public*/, output [7:0] O_149/*verilator public*/, output [7:0] O_15/*verilator public*/, output [7:0] O_150/*verilator public*/, output [7:0] O_151/*verilator public*/, output [7:0] O_152/*verilator public*/, output [7:0] O_153/*verilator public*/, output [7:0] O_154/*verilator public*/, output [7:0] O_155/*verilator public*/, output [7:0] O_156/*verilator public*/, output [7:0] O_157/*verilator public*/, output [7:0] O_158/*verilator public*/, output [7:0] O_159/*verilator public*/, output [7:0] O_16/*verilator public*/, output [7:0] O_160/*verilator public*/, output [7:0] O_161/*verilator public*/, output [7:0] O_162/*verilator public*/, output [7:0] O_163/*verilator public*/, output [7:0] O_164/*verilator public*/, output [7:0] O_165/*verilator public*/, output [7:0] O_166/*verilator public*/, output [7:0] O_167/*verilator public*/, output [7:0] O_168/*verilator public*/, output [7:0] O_169/*verilator public*/, output [7:0] O_17/*verilator public*/, output [7:0] O_170/*verilator public*/, output [7:0] O_171/*verilator public*/, output [7:0] O_172/*verilator public*/, output [7:0] O_173/*verilator public*/, output [7:0] O_174/*verilator public*/, output [7:0] O_175/*verilator public*/, output [7:0] O_176/*verilator public*/, output [7:0] O_177/*verilator public*/, output [7:0] O_178/*verilator public*/, output [7:0] O_179/*verilator public*/, output [7:0] O_18/*verilator public*/, output [7:0] O_180/*verilator public*/, output [7:0] O_181/*verilator public*/, output [7:0] O_182/*verilator public*/, output [7:0] O_183/*verilator public*/, output [7:0] O_184/*verilator public*/, output [7:0] O_185/*verilator public*/, output [7:0] O_186/*verilator public*/, output [7:0] O_187/*verilator public*/, output [7:0] O_188/*verilator public*/, output [7:0] O_189/*verilator public*/, output [7:0] O_19/*verilator public*/, output [7:0] O_190/*verilator public*/, output [7:0] O_191/*verilator public*/, output [7:0] O_192/*verilator public*/, output [7:0] O_193/*verilator public*/, output [7:0] O_194/*verilator public*/, output [7:0] O_195/*verilator public*/, output [7:0] O_196/*verilator public*/, output [7:0] O_197/*verilator public*/, output [7:0] O_198/*verilator public*/, output [7:0] O_199/*verilator public*/, output [7:0] O_2/*verilator public*/, output [7:0] O_20/*verilator public*/, output [7:0] O_21/*verilator public*/, output [7:0] O_22/*verilator public*/, output [7:0] O_23/*verilator public*/, output [7:0] O_24/*verilator public*/, output [7:0] O_25/*verilator public*/, output [7:0] O_26/*verilator public*/, output [7:0] O_27/*verilator public*/, output [7:0] O_28/*verilator public*/, output [7:0] O_29/*verilator public*/, output [7:0] O_3/*verilator public*/, output [7:0] O_30/*verilator public*/, output [7:0] O_31/*verilator public*/, output [7:0] O_32/*verilator public*/, output [7:0] O_33/*verilator public*/, output [7:0] O_34/*verilator public*/, output [7:0] O_35/*verilator public*/, output [7:0] O_36/*verilator public*/, output [7:0] O_37/*verilator public*/, output [7:0] O_38/*verilator public*/, output [7:0] O_39/*verilator public*/, output [7:0] O_4/*verilator public*/, output [7:0] O_40/*verilator public*/, output [7:0] O_41/*verilator public*/, output [7:0] O_42/*verilator public*/, output [7:0] O_43/*verilator public*/, output [7:0] O_44/*verilator public*/, output [7:0] O_45/*verilator public*/, output [7:0] O_46/*verilator public*/, output [7:0] O_47/*verilator public*/, output [7:0] O_48/*verilator public*/, output [7:0] O_49/*verilator public*/, output [7:0] O_5/*verilator public*/, output [7:0] O_50/*verilator public*/, output [7:0] O_51/*verilator public*/, output [7:0] O_52/*verilator public*/, output [7:0] O_53/*verilator public*/, output [7:0] O_54/*verilator public*/, output [7:0] O_55/*verilator public*/, output [7:0] O_56/*verilator public*/, output [7:0] O_57/*verilator public*/, output [7:0] O_58/*verilator public*/, output [7:0] O_59/*verilator public*/, output [7:0] O_6/*verilator public*/, output [7:0] O_60/*verilator public*/, output [7:0] O_61/*verilator public*/, output [7:0] O_62/*verilator public*/, output [7:0] O_63/*verilator public*/, output [7:0] O_64/*verilator public*/, output [7:0] O_65/*verilator public*/, output [7:0] O_66/*verilator public*/, output [7:0] O_67/*verilator public*/, output [7:0] O_68/*verilator public*/, output [7:0] O_69/*verilator public*/, output [7:0] O_7/*verilator public*/, output [7:0] O_70/*verilator public*/, output [7:0] O_71/*verilator public*/, output [7:0] O_72/*verilator public*/, output [7:0] O_73/*verilator public*/, output [7:0] O_74/*verilator public*/, output [7:0] O_75/*verilator public*/, output [7:0] O_76/*verilator public*/, output [7:0] O_77/*verilator public*/, output [7:0] O_78/*verilator public*/, output [7:0] O_79/*verilator public*/, output [7:0] O_8/*verilator public*/, output [7:0] O_80/*verilator public*/, output [7:0] O_81/*verilator public*/, output [7:0] O_82/*verilator public*/, output [7:0] O_83/*verilator public*/, output [7:0] O_84/*verilator public*/, output [7:0] O_85/*verilator public*/, output [7:0] O_86/*verilator public*/, output [7:0] O_87/*verilator public*/, output [7:0] O_88/*verilator public*/, output [7:0] O_89/*verilator public*/, output [7:0] O_9/*verilator public*/, output [7:0] O_90/*verilator public*/, output [7:0] O_91/*verilator public*/, output [7:0] O_92/*verilator public*/, output [7:0] O_93/*verilator public*/, output [7:0] O_94/*verilator public*/, output [7:0] O_95/*verilator public*/, output [7:0] O_96/*verilator public*/, output [7:0] O_97/*verilator public*/, output [7:0] O_98/*verilator public*/, output [7:0] O_99/*verilator public*/, input [7:0] hi_0/*verilator public*/, input [7:0] hi_1/*verilator public*/, input [7:0] hi_10/*verilator public*/, input [7:0] hi_100/*verilator public*/, input [7:0] hi_101/*verilator public*/, input [7:0] hi_102/*verilator public*/, input [7:0] hi_103/*verilator public*/, input [7:0] hi_104/*verilator public*/, input [7:0] hi_105/*verilator public*/, input [7:0] hi_106/*verilator public*/, input [7:0] hi_107/*verilator public*/, input [7:0] hi_108/*verilator public*/, input [7:0] hi_109/*verilator public*/, input [7:0] hi_11/*verilator public*/, input [7:0] hi_110/*verilator public*/, input [7:0] hi_111/*verilator public*/, input [7:0] hi_112/*verilator public*/, input [7:0] hi_113/*verilator public*/, input [7:0] hi_114/*verilator public*/, input [7:0] hi_115/*verilator public*/, input [7:0] hi_116/*verilator public*/, input [7:0] hi_117/*verilator public*/, input [7:0] hi_118/*verilator public*/, input [7:0] hi_119/*verilator public*/, input [7:0] hi_12/*verilator public*/, input [7:0] hi_120/*verilator public*/, input [7:0] hi_121/*verilator public*/, input [7:0] hi_122/*verilator public*/, input [7:0] hi_123/*verilator public*/, input [7:0] hi_124/*verilator public*/, input [7:0] hi_125/*verilator public*/, input [7:0] hi_126/*verilator public*/, input [7:0] hi_127/*verilator public*/, input [7:0] hi_128/*verilator public*/, input [7:0] hi_129/*verilator public*/, input [7:0] hi_13/*verilator public*/, input [7:0] hi_130/*verilator public*/, input [7:0] hi_131/*verilator public*/, input [7:0] hi_132/*verilator public*/, input [7:0] hi_133/*verilator public*/, input [7:0] hi_134/*verilator public*/, input [7:0] hi_135/*verilator public*/, input [7:0] hi_136/*verilator public*/, input [7:0] hi_137/*verilator public*/, input [7:0] hi_138/*verilator public*/, input [7:0] hi_139/*verilator public*/, input [7:0] hi_14/*verilator public*/, input [7:0] hi_140/*verilator public*/, input [7:0] hi_141/*verilator public*/, input [7:0] hi_142/*verilator public*/, input [7:0] hi_143/*verilator public*/, input [7:0] hi_144/*verilator public*/, input [7:0] hi_145/*verilator public*/, input [7:0] hi_146/*verilator public*/, input [7:0] hi_147/*verilator public*/, input [7:0] hi_148/*verilator public*/, input [7:0] hi_149/*verilator public*/, input [7:0] hi_15/*verilator public*/, input [7:0] hi_150/*verilator public*/, input [7:0] hi_151/*verilator public*/, input [7:0] hi_152/*verilator public*/, input [7:0] hi_153/*verilator public*/, input [7:0] hi_154/*verilator public*/, input [7:0] hi_155/*verilator public*/, input [7:0] hi_156/*verilator public*/, input [7:0] hi_157/*verilator public*/, input [7:0] hi_158/*verilator public*/, input [7:0] hi_159/*verilator public*/, input [7:0] hi_16/*verilator public*/, input [7:0] hi_160/*verilator public*/, input [7:0] hi_161/*verilator public*/, input [7:0] hi_162/*verilator public*/, input [7:0] hi_163/*verilator public*/, input [7:0] hi_164/*verilator public*/, input [7:0] hi_165/*verilator public*/, input [7:0] hi_166/*verilator public*/, input [7:0] hi_167/*verilator public*/, input [7:0] hi_168/*verilator public*/, input [7:0] hi_169/*verilator public*/, input [7:0] hi_17/*verilator public*/, input [7:0] hi_170/*verilator public*/, input [7:0] hi_171/*verilator public*/, input [7:0] hi_172/*verilator public*/, input [7:0] hi_173/*verilator public*/, input [7:0] hi_174/*verilator public*/, input [7:0] hi_175/*verilator public*/, input [7:0] hi_176/*verilator public*/, input [7:0] hi_177/*verilator public*/, input [7:0] hi_178/*verilator public*/, input [7:0] hi_179/*verilator public*/, input [7:0] hi_18/*verilator public*/, input [7:0] hi_180/*verilator public*/, input [7:0] hi_181/*verilator public*/, input [7:0] hi_182/*verilator public*/, input [7:0] hi_183/*verilator public*/, input [7:0] hi_184/*verilator public*/, input [7:0] hi_185/*verilator public*/, input [7:0] hi_186/*verilator public*/, input [7:0] hi_187/*verilator public*/, input [7:0] hi_188/*verilator public*/, input [7:0] hi_189/*verilator public*/, input [7:0] hi_19/*verilator public*/, input [7:0] hi_190/*verilator public*/, input [7:0] hi_191/*verilator public*/, input [7:0] hi_192/*verilator public*/, input [7:0] hi_193/*verilator public*/, input [7:0] hi_194/*verilator public*/, input [7:0] hi_195/*verilator public*/, input [7:0] hi_196/*verilator public*/, input [7:0] hi_197/*verilator public*/, input [7:0] hi_198/*verilator public*/, input [7:0] hi_199/*verilator public*/, input [7:0] hi_2/*verilator public*/, input [7:0] hi_20/*verilator public*/, input [7:0] hi_21/*verilator public*/, input [7:0] hi_22/*verilator public*/, input [7:0] hi_23/*verilator public*/, input [7:0] hi_24/*verilator public*/, input [7:0] hi_25/*verilator public*/, input [7:0] hi_26/*verilator public*/, input [7:0] hi_27/*verilator public*/, input [7:0] hi_28/*verilator public*/, input [7:0] hi_29/*verilator public*/, input [7:0] hi_3/*verilator public*/, input [7:0] hi_30/*verilator public*/, input [7:0] hi_31/*verilator public*/, input [7:0] hi_32/*verilator public*/, input [7:0] hi_33/*verilator public*/, input [7:0] hi_34/*verilator public*/, input [7:0] hi_35/*verilator public*/, input [7:0] hi_36/*verilator public*/, input [7:0] hi_37/*verilator public*/, input [7:0] hi_38/*verilator public*/, input [7:0] hi_39/*verilator public*/, input [7:0] hi_4/*verilator public*/, input [7:0] hi_40/*verilator public*/, input [7:0] hi_41/*verilator public*/, input [7:0] hi_42/*verilator public*/, input [7:0] hi_43/*verilator public*/, input [7:0] hi_44/*verilator public*/, input [7:0] hi_45/*verilator public*/, input [7:0] hi_46/*verilator public*/, input [7:0] hi_47/*verilator public*/, input [7:0] hi_48/*verilator public*/, input [7:0] hi_49/*verilator public*/, input [7:0] hi_5/*verilator public*/, input [7:0] hi_50/*verilator public*/, input [7:0] hi_51/*verilator public*/, input [7:0] hi_52/*verilator public*/, input [7:0] hi_53/*verilator public*/, input [7:0] hi_54/*verilator public*/, input [7:0] hi_55/*verilator public*/, input [7:0] hi_56/*verilator public*/, input [7:0] hi_57/*verilator public*/, input [7:0] hi_58/*verilator public*/, input [7:0] hi_59/*verilator public*/, input [7:0] hi_6/*verilator public*/, input [7:0] hi_60/*verilator public*/, input [7:0] hi_61/*verilator public*/, input [7:0] hi_62/*verilator public*/, input [7:0] hi_63/*verilator public*/, input [7:0] hi_64/*verilator public*/, input [7:0] hi_65/*verilator public*/, input [7:0] hi_66/*verilator public*/, input [7:0] hi_67/*verilator public*/, input [7:0] hi_68/*verilator public*/, input [7:0] hi_69/*verilator public*/, input [7:0] hi_7/*verilator public*/, input [7:0] hi_70/*verilator public*/, input [7:0] hi_71/*verilator public*/, input [7:0] hi_72/*verilator public*/, input [7:0] hi_73/*verilator public*/, input [7:0] hi_74/*verilator public*/, input [7:0] hi_75/*verilator public*/, input [7:0] hi_76/*verilator public*/, input [7:0] hi_77/*verilator public*/, input [7:0] hi_78/*verilator public*/, input [7:0] hi_79/*verilator public*/, input [7:0] hi_8/*verilator public*/, input [7:0] hi_80/*verilator public*/, input [7:0] hi_81/*verilator public*/, input [7:0] hi_82/*verilator public*/, input [7:0] hi_83/*verilator public*/, input [7:0] hi_84/*verilator public*/, input [7:0] hi_85/*verilator public*/, input [7:0] hi_86/*verilator public*/, input [7:0] hi_87/*verilator public*/, input [7:0] hi_88/*verilator public*/, input [7:0] hi_89/*verilator public*/, input [7:0] hi_9/*verilator public*/, input [7:0] hi_90/*verilator public*/, input [7:0] hi_91/*verilator public*/, input [7:0] hi_92/*verilator public*/, input [7:0] hi_93/*verilator public*/, input [7:0] hi_94/*verilator public*/, input [7:0] hi_95/*verilator public*/, input [7:0] hi_96/*verilator public*/, input [7:0] hi_97/*verilator public*/, input [7:0] hi_98/*verilator public*/, input [7:0] hi_99/*verilator public*/, output valid_down/*verilator public*/, input valid_up/*verilator public*/);
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_100;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_101;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_102;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_103;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_104;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_105;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_106;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_107;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_108;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_109;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_110;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_111;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_112;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_113;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_114;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_115;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_116;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_117;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_118;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_119;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_120;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_121;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_122;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_123;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_124;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_125;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_126;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_127;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_128;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_129;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_130;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_131;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_132;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_133;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_134;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_135;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_136;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_137;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_138;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_139;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_140;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_141;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_142;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_143;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_144;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_145;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_146;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_147;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_148;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_149;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_150;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_151;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_152;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_153;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_154;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_155;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_156;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_157;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_158;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_159;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_160;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_161;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_162;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_163;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_164;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_165;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_166;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_167;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_168;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_169;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_170;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_171;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_172;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_173;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_174;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_175;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_176;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_177;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_178;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_179;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_180;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_181;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_182;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_183;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_184;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_185;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_186;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_187;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_188;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_189;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_190;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_191;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_192;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_193;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_194;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_195;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_196;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_197;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_198;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_199;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_40;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_41;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_42;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_43;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_44;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_45;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_46;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_47;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_48;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_49;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_50;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_51;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_52;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_53;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_54;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_55;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_56;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_57;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_58;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_59;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_60;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_61;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_62;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_63;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_64;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_65;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_66;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_67;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_68;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_69;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_70;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_71;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_72;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_73;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_74;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_75;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_76;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_77;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_78;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_79;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_80;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_81;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_82;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_83;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_84;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_85;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_86;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_87;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_88;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_89;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_90;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_91;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_92;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_93;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_94;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_95;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_96;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_97;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_98;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_99;
wire FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_100;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_101;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_102;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_103;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_104;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_105;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_106;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_107;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_108;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_109;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_110;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_111;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_112;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_113;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_114;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_115;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_116;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_117;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_118;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_119;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_120;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_121;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_122;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_123;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_124;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_125;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_126;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_127;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_128;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_129;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_130;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_131;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_132;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_133;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_134;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_135;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_136;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_137;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_138;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_139;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_140;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_141;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_142;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_143;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_144;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_145;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_146;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_147;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_148;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_149;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_150;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_151;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_152;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_153;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_154;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_155;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_156;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_157;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_158;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_159;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_160;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_161;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_162;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_163;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_164;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_165;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_166;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_167;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_168;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_169;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_170;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_171;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_172;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_173;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_174;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_175;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_176;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_177;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_178;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_179;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_180;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_181;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_182;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_183;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_184;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_185;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_186;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_187;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_188;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_189;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_190;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_191;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_192;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_193;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_194;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_195;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_196;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_197;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_198;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_199;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_40;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_41;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_42;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_43;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_44;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_45;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_46;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_47;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_48;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_49;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_50;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_51;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_52;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_53;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_54;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_55;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_56;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_57;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_58;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_59;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_60;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_61;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_62;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_63;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_64;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_65;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_66;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_67;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_68;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_69;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_70;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_71;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_72;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_73;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_74;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_75;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_76;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_77;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_78;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_79;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_80;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_81;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_82;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_83;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_84;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_85;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_86;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_87;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_88;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_89;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_90;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_91;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_92;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_93;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_94;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_95;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_96;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_97;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_98;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_99;
wire FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_100;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_101;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_102;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_103;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_104;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_105;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_106;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_107;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_108;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_109;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_110;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_111;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_112;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_113;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_114;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_115;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_116;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_117;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_118;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_119;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_120;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_121;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_122;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_123;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_124;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_125;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_126;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_127;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_128;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_129;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_130;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_131;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_132;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_133;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_134;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_135;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_136;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_137;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_138;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_139;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_140;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_141;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_142;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_143;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_144;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_145;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_146;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_147;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_148;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_149;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_150;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_151;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_152;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_153;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_154;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_155;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_156;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_157;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_158;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_159;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_160;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_161;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_162;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_163;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_164;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_165;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_166;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_167;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_168;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_169;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_170;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_171;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_172;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_173;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_174;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_175;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_176;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_177;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_178;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_179;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_180;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_181;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_182;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_183;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_184;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_185;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_186;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_187;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_188;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_189;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_190;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_191;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_192;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_193;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_194;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_195;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_196;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_197;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_198;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_199;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_40;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_41;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_42;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_43;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_44;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_45;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_46;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_47;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_48;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_49;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_50;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_51;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_52;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_53;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_54;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_55;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_56;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_57;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_58;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_59;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_60;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_61;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_62;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_63;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_64;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_65;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_66;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_67;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_68;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_69;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_70;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_71;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_72;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_73;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_74;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_75;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_76;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_77;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_78;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_79;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_80;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_81;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_82;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_83;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_84;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_85;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_86;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_87;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_88;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_89;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_90;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_91;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_92;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_93;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_94;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_95;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_96;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_97;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_98;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_99;
wire FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_100;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_101;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_102;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_103;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_104;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_105;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_106;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_107;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_108;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_109;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_110;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_111;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_112;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_113;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_114;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_115;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_116;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_117;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_118;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_119;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_120;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_121;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_122;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_123;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_124;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_125;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_126;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_127;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_128;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_129;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_130;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_131;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_132;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_133;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_134;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_135;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_136;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_137;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_138;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_139;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_140;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_141;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_142;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_143;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_144;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_145;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_146;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_147;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_148;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_149;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_150;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_151;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_152;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_153;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_154;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_155;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_156;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_157;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_158;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_159;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_160;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_161;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_162;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_163;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_164;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_165;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_166;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_167;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_168;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_169;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_170;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_171;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_172;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_173;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_174;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_175;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_176;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_177;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_178;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_179;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_180;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_181;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_182;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_183;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_184;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_185;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_186;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_187;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_188;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_189;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_190;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_191;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_192;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_193;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_194;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_195;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_196;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_197;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_198;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_199;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_20;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_21;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_22;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_23;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_24;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_25;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_26;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_27;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_28;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_29;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_30;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_31;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_32;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_33;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_34;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_35;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_36;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_37;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_38;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_39;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_40;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_41;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_42;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_43;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_44;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_45;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_46;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_47;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_48;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_49;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_50;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_51;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_52;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_53;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_54;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_55;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_56;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_57;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_58;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_59;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_60;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_61;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_62;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_63;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_64;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_65;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_66;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_67;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_68;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_69;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_70;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_71;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_72;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_73;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_74;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_75;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_76;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_77;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_78;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_79;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_80;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_81;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_82;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_83;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_84;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_85;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_86;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_87;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_88;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_89;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_90;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_91;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_92;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_93;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_94;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_95;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_96;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_97;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_98;
wire [7:0] FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_99;
wire FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_100;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_101;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_102;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_103;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_104;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_105;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_106;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_107;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_108;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_109;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_110;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_111;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_112;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_113;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_114;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_115;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_116;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_117;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_118;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_119;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_120;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_121;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_122;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_123;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_124;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_125;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_126;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_127;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_128;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_129;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_130;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_131;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_132;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_133;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_134;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_135;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_136;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_137;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_138;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_139;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_140;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_141;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_142;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_143;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_144;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_145;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_146;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_147;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_148;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_149;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_150;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_151;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_152;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_153;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_154;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_155;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_156;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_157;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_158;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_159;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_160;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_161;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_162;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_163;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_164;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_165;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_166;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_167;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_168;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_169;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_170;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_171;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_172;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_173;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_174;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_175;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_176;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_177;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_178;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_179;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_180;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_181;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_182;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_183;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_184;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_185;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_186;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_187;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_188;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_189;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_190;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_191;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_192;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_193;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_194;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_195;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_196;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_197;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_198;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_199;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_40;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_41;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_42;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_43;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_44;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_45;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_46;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_47;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_48;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_49;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_50;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_51;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_52;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_53;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_54;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_55;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_56;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_57;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_58;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_59;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_60;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_61;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_62;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_63;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_64;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_65;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_66;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_67;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_68;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_69;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_70;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_71;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_72;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_73;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_74;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_75;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_76;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_77;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_78;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_79;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_80;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_81;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_82;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_83;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_84;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_85;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_86;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_87;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_88;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_89;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_90;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_91;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_92;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_93;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_94;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_95;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_96;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_97;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_98;
wire [7:0] NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_99;
wire NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down;
FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0(.CLK(CLK), .I_0(hi_0), .I_1(hi_1), .I_10(hi_10), .I_100(hi_100), .I_101(hi_101), .I_102(hi_102), .I_103(hi_103), .I_104(hi_104), .I_105(hi_105), .I_106(hi_106), .I_107(hi_107), .I_108(hi_108), .I_109(hi_109), .I_11(hi_11), .I_110(hi_110), .I_111(hi_111), .I_112(hi_112), .I_113(hi_113), .I_114(hi_114), .I_115(hi_115), .I_116(hi_116), .I_117(hi_117), .I_118(hi_118), .I_119(hi_119), .I_12(hi_12), .I_120(hi_120), .I_121(hi_121), .I_122(hi_122), .I_123(hi_123), .I_124(hi_124), .I_125(hi_125), .I_126(hi_126), .I_127(hi_127), .I_128(hi_128), .I_129(hi_129), .I_13(hi_13), .I_130(hi_130), .I_131(hi_131), .I_132(hi_132), .I_133(hi_133), .I_134(hi_134), .I_135(hi_135), .I_136(hi_136), .I_137(hi_137), .I_138(hi_138), .I_139(hi_139), .I_14(hi_14), .I_140(hi_140), .I_141(hi_141), .I_142(hi_142), .I_143(hi_143), .I_144(hi_144), .I_145(hi_145), .I_146(hi_146), .I_147(hi_147), .I_148(hi_148), .I_149(hi_149), .I_15(hi_15), .I_150(hi_150), .I_151(hi_151), .I_152(hi_152), .I_153(hi_153), .I_154(hi_154), .I_155(hi_155), .I_156(hi_156), .I_157(hi_157), .I_158(hi_158), .I_159(hi_159), .I_16(hi_16), .I_160(hi_160), .I_161(hi_161), .I_162(hi_162), .I_163(hi_163), .I_164(hi_164), .I_165(hi_165), .I_166(hi_166), .I_167(hi_167), .I_168(hi_168), .I_169(hi_169), .I_17(hi_17), .I_170(hi_170), .I_171(hi_171), .I_172(hi_172), .I_173(hi_173), .I_174(hi_174), .I_175(hi_175), .I_176(hi_176), .I_177(hi_177), .I_178(hi_178), .I_179(hi_179), .I_18(hi_18), .I_180(hi_180), .I_181(hi_181), .I_182(hi_182), .I_183(hi_183), .I_184(hi_184), .I_185(hi_185), .I_186(hi_186), .I_187(hi_187), .I_188(hi_188), .I_189(hi_189), .I_19(hi_19), .I_190(hi_190), .I_191(hi_191), .I_192(hi_192), .I_193(hi_193), .I_194(hi_194), .I_195(hi_195), .I_196(hi_196), .I_197(hi_197), .I_198(hi_198), .I_199(hi_199), .I_2(hi_2), .I_20(hi_20), .I_21(hi_21), .I_22(hi_22), .I_23(hi_23), .I_24(hi_24), .I_25(hi_25), .I_26(hi_26), .I_27(hi_27), .I_28(hi_28), .I_29(hi_29), .I_3(hi_3), .I_30(hi_30), .I_31(hi_31), .I_32(hi_32), .I_33(hi_33), .I_34(hi_34), .I_35(hi_35), .I_36(hi_36), .I_37(hi_37), .I_38(hi_38), .I_39(hi_39), .I_4(hi_4), .I_40(hi_40), .I_41(hi_41), .I_42(hi_42), .I_43(hi_43), .I_44(hi_44), .I_45(hi_45), .I_46(hi_46), .I_47(hi_47), .I_48(hi_48), .I_49(hi_49), .I_5(hi_5), .I_50(hi_50), .I_51(hi_51), .I_52(hi_52), .I_53(hi_53), .I_54(hi_54), .I_55(hi_55), .I_56(hi_56), .I_57(hi_57), .I_58(hi_58), .I_59(hi_59), .I_6(hi_6), .I_60(hi_60), .I_61(hi_61), .I_62(hi_62), .I_63(hi_63), .I_64(hi_64), .I_65(hi_65), .I_66(hi_66), .I_67(hi_67), .I_68(hi_68), .I_69(hi_69), .I_7(hi_7), .I_70(hi_70), .I_71(hi_71), .I_72(hi_72), .I_73(hi_73), .I_74(hi_74), .I_75(hi_75), .I_76(hi_76), .I_77(hi_77), .I_78(hi_78), .I_79(hi_79), .I_8(hi_8), .I_80(hi_80), .I_81(hi_81), .I_82(hi_82), .I_83(hi_83), .I_84(hi_84), .I_85(hi_85), .I_86(hi_86), .I_87(hi_87), .I_88(hi_88), .I_89(hi_89), .I_9(hi_9), .I_90(hi_90), .I_91(hi_91), .I_92(hi_92), .I_93(hi_93), .I_94(hi_94), .I_95(hi_95), .I_96(hi_96), .I_97(hi_97), .I_98(hi_98), .I_99(hi_99), .O_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .O_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .O_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10), .O_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_100), .O_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_101), .O_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_102), .O_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_103), .O_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_104), .O_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_105), .O_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_106), .O_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_107), .O_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_108), .O_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_109), .O_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11), .O_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_110), .O_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_111), .O_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_112), .O_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_113), .O_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_114), .O_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_115), .O_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_116), .O_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_117), .O_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_118), .O_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_119), .O_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12), .O_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_120), .O_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_121), .O_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_122), .O_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_123), .O_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_124), .O_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_125), .O_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_126), .O_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_127), .O_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_128), .O_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_129), .O_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13), .O_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_130), .O_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_131), .O_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_132), .O_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_133), .O_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_134), .O_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_135), .O_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_136), .O_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_137), .O_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_138), .O_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_139), .O_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14), .O_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_140), .O_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_141), .O_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_142), .O_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_143), .O_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_144), .O_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_145), .O_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_146), .O_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_147), .O_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_148), .O_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_149), .O_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15), .O_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_150), .O_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_151), .O_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_152), .O_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_153), .O_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_154), .O_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_155), .O_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_156), .O_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_157), .O_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_158), .O_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_159), .O_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16), .O_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_160), .O_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_161), .O_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_162), .O_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_163), .O_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_164), .O_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_165), .O_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_166), .O_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_167), .O_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_168), .O_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_169), .O_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17), .O_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_170), .O_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_171), .O_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_172), .O_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_173), .O_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_174), .O_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_175), .O_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_176), .O_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_177), .O_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_178), .O_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_179), .O_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18), .O_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_180), .O_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_181), .O_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_182), .O_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_183), .O_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_184), .O_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_185), .O_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_186), .O_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_187), .O_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_188), .O_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_189), .O_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19), .O_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_190), .O_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_191), .O_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_192), .O_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_193), .O_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_194), .O_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_195), .O_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_196), .O_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_197), .O_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_198), .O_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_199), .O_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .O_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20), .O_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21), .O_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22), .O_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23), .O_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24), .O_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25), .O_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26), .O_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27), .O_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28), .O_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29), .O_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3), .O_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30), .O_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31), .O_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32), .O_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33), .O_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34), .O_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35), .O_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36), .O_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37), .O_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38), .O_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39), .O_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4), .O_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_40), .O_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_41), .O_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_42), .O_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_43), .O_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_44), .O_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_45), .O_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_46), .O_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_47), .O_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_48), .O_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_49), .O_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5), .O_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_50), .O_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_51), .O_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_52), .O_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_53), .O_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_54), .O_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_55), .O_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_56), .O_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_57), .O_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_58), .O_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_59), .O_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6), .O_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_60), .O_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_61), .O_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_62), .O_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_63), .O_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_64), .O_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_65), .O_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_66), .O_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_67), .O_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_68), .O_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_69), .O_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7), .O_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_70), .O_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_71), .O_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_72), .O_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_73), .O_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_74), .O_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_75), .O_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_76), .O_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_77), .O_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_78), .O_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_79), .O_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8), .O_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_80), .O_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_81), .O_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_82), .O_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_83), .O_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_84), .O_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_85), .O_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_86), .O_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_87), .O_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_88), .O_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_89), .O_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9), .O_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_90), .O_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_91), .O_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_92), .O_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_93), .O_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_94), .O_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_95), .O_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_96), .O_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_97), .O_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_98), .O_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_99), .valid_down(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down), .valid_up(valid_up));
FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1(.CLK(CLK), .I_0(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .I_1(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .I_10(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .I_100(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_100), .I_101(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_101), .I_102(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_102), .I_103(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_103), .I_104(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_104), .I_105(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_105), .I_106(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_106), .I_107(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_107), .I_108(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_108), .I_109(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_109), .I_11(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .I_110(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_110), .I_111(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_111), .I_112(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_112), .I_113(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_113), .I_114(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_114), .I_115(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_115), .I_116(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_116), .I_117(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_117), .I_118(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_118), .I_119(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_119), .I_12(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .I_120(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_120), .I_121(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_121), .I_122(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_122), .I_123(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_123), .I_124(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_124), .I_125(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_125), .I_126(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_126), .I_127(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_127), .I_128(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_128), .I_129(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_129), .I_13(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .I_130(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_130), .I_131(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_131), .I_132(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_132), .I_133(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_133), .I_134(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_134), .I_135(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_135), .I_136(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_136), .I_137(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_137), .I_138(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_138), .I_139(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_139), .I_14(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .I_140(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_140), .I_141(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_141), .I_142(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_142), .I_143(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_143), .I_144(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_144), .I_145(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_145), .I_146(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_146), .I_147(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_147), .I_148(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_148), .I_149(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_149), .I_15(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .I_150(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_150), .I_151(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_151), .I_152(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_152), .I_153(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_153), .I_154(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_154), .I_155(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_155), .I_156(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_156), .I_157(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_157), .I_158(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_158), .I_159(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_159), .I_16(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .I_160(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_160), .I_161(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_161), .I_162(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_162), .I_163(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_163), .I_164(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_164), .I_165(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_165), .I_166(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_166), .I_167(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_167), .I_168(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_168), .I_169(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_169), .I_17(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .I_170(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_170), .I_171(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_171), .I_172(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_172), .I_173(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_173), .I_174(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_174), .I_175(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_175), .I_176(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_176), .I_177(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_177), .I_178(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_178), .I_179(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_179), .I_18(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .I_180(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_180), .I_181(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_181), .I_182(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_182), .I_183(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_183), .I_184(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_184), .I_185(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_185), .I_186(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_186), .I_187(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_187), .I_188(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_188), .I_189(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_189), .I_19(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .I_190(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_190), .I_191(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_191), .I_192(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_192), .I_193(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_193), .I_194(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_194), .I_195(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_195), .I_196(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_196), .I_197(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_197), .I_198(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_198), .I_199(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_199), .I_2(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .I_20(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20), .I_21(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21), .I_22(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22), .I_23(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23), .I_24(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24), .I_25(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25), .I_26(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26), .I_27(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27), .I_28(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28), .I_29(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29), .I_3(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .I_30(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30), .I_31(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31), .I_32(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32), .I_33(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33), .I_34(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34), .I_35(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35), .I_36(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36), .I_37(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37), .I_38(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38), .I_39(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39), .I_4(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .I_40(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_40), .I_41(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_41), .I_42(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_42), .I_43(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_43), .I_44(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_44), .I_45(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_45), .I_46(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_46), .I_47(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_47), .I_48(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_48), .I_49(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_49), .I_5(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .I_50(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_50), .I_51(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_51), .I_52(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_52), .I_53(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_53), .I_54(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_54), .I_55(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_55), .I_56(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_56), .I_57(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_57), .I_58(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_58), .I_59(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_59), .I_6(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .I_60(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_60), .I_61(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_61), .I_62(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_62), .I_63(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_63), .I_64(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_64), .I_65(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_65), .I_66(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_66), .I_67(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_67), .I_68(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_68), .I_69(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_69), .I_7(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .I_70(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_70), .I_71(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_71), .I_72(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_72), .I_73(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_73), .I_74(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_74), .I_75(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_75), .I_76(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_76), .I_77(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_77), .I_78(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_78), .I_79(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_79), .I_8(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .I_80(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_80), .I_81(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_81), .I_82(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_82), .I_83(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_83), .I_84(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_84), .I_85(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_85), .I_86(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_86), .I_87(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_87), .I_88(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_88), .I_89(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_89), .I_9(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .I_90(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_90), .I_91(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_91), .I_92(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_92), .I_93(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_93), .I_94(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_94), .I_95(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_95), .I_96(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_96), .I_97(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_97), .I_98(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_98), .I_99(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_99), .O_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .O_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1), .O_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10), .O_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_100), .O_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_101), .O_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_102), .O_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_103), .O_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_104), .O_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_105), .O_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_106), .O_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_107), .O_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_108), .O_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_109), .O_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11), .O_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_110), .O_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_111), .O_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_112), .O_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_113), .O_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_114), .O_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_115), .O_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_116), .O_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_117), .O_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_118), .O_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_119), .O_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12), .O_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_120), .O_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_121), .O_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_122), .O_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_123), .O_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_124), .O_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_125), .O_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_126), .O_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_127), .O_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_128), .O_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_129), .O_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13), .O_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_130), .O_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_131), .O_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_132), .O_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_133), .O_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_134), .O_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_135), .O_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_136), .O_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_137), .O_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_138), .O_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_139), .O_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14), .O_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_140), .O_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_141), .O_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_142), .O_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_143), .O_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_144), .O_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_145), .O_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_146), .O_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_147), .O_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_148), .O_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_149), .O_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15), .O_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_150), .O_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_151), .O_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_152), .O_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_153), .O_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_154), .O_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_155), .O_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_156), .O_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_157), .O_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_158), .O_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_159), .O_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16), .O_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_160), .O_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_161), .O_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_162), .O_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_163), .O_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_164), .O_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_165), .O_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_166), .O_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_167), .O_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_168), .O_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_169), .O_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17), .O_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_170), .O_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_171), .O_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_172), .O_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_173), .O_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_174), .O_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_175), .O_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_176), .O_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_177), .O_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_178), .O_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_179), .O_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18), .O_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_180), .O_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_181), .O_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_182), .O_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_183), .O_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_184), .O_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_185), .O_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_186), .O_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_187), .O_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_188), .O_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_189), .O_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19), .O_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_190), .O_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_191), .O_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_192), .O_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_193), .O_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_194), .O_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_195), .O_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_196), .O_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_197), .O_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_198), .O_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_199), .O_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2), .O_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20), .O_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21), .O_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22), .O_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23), .O_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24), .O_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25), .O_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26), .O_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27), .O_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28), .O_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29), .O_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3), .O_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30), .O_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31), .O_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32), .O_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33), .O_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34), .O_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35), .O_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36), .O_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37), .O_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38), .O_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39), .O_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4), .O_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_40), .O_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_41), .O_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_42), .O_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_43), .O_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_44), .O_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_45), .O_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_46), .O_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_47), .O_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_48), .O_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_49), .O_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5), .O_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_50), .O_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_51), .O_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_52), .O_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_53), .O_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_54), .O_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_55), .O_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_56), .O_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_57), .O_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_58), .O_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_59), .O_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6), .O_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_60), .O_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_61), .O_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_62), .O_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_63), .O_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_64), .O_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_65), .O_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_66), .O_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_67), .O_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_68), .O_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_69), .O_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7), .O_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_70), .O_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_71), .O_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_72), .O_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_73), .O_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_74), .O_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_75), .O_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_76), .O_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_77), .O_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_78), .O_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_79), .O_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8), .O_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_80), .O_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_81), .O_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_82), .O_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_83), .O_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_84), .O_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_85), .O_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_86), .O_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_87), .O_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_88), .O_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_89), .O_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9), .O_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_90), .O_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_91), .O_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_92), .O_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_93), .O_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_94), .O_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_95), .O_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_96), .O_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_97), .O_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_98), .O_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_99), .valid_down(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down), .valid_up(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down));
FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2(.CLK(CLK), .I_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_0), .I_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_1), .I_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_10), .I_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_100), .I_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_101), .I_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_102), .I_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_103), .I_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_104), .I_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_105), .I_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_106), .I_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_107), .I_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_108), .I_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_109), .I_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_11), .I_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_110), .I_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_111), .I_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_112), .I_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_113), .I_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_114), .I_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_115), .I_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_116), .I_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_117), .I_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_118), .I_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_119), .I_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_12), .I_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_120), .I_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_121), .I_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_122), .I_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_123), .I_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_124), .I_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_125), .I_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_126), .I_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_127), .I_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_128), .I_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_129), .I_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_13), .I_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_130), .I_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_131), .I_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_132), .I_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_133), .I_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_134), .I_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_135), .I_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_136), .I_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_137), .I_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_138), .I_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_139), .I_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_14), .I_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_140), .I_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_141), .I_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_142), .I_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_143), .I_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_144), .I_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_145), .I_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_146), .I_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_147), .I_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_148), .I_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_149), .I_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_15), .I_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_150), .I_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_151), .I_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_152), .I_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_153), .I_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_154), .I_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_155), .I_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_156), .I_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_157), .I_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_158), .I_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_159), .I_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_16), .I_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_160), .I_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_161), .I_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_162), .I_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_163), .I_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_164), .I_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_165), .I_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_166), .I_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_167), .I_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_168), .I_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_169), .I_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_17), .I_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_170), .I_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_171), .I_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_172), .I_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_173), .I_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_174), .I_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_175), .I_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_176), .I_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_177), .I_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_178), .I_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_179), .I_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_18), .I_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_180), .I_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_181), .I_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_182), .I_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_183), .I_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_184), .I_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_185), .I_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_186), .I_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_187), .I_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_188), .I_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_189), .I_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_19), .I_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_190), .I_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_191), .I_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_192), .I_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_193), .I_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_194), .I_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_195), .I_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_196), .I_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_197), .I_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_198), .I_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_199), .I_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_2), .I_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_20), .I_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_21), .I_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_22), .I_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_23), .I_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_24), .I_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_25), .I_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_26), .I_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_27), .I_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_28), .I_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_29), .I_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_3), .I_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_30), .I_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_31), .I_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_32), .I_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_33), .I_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_34), .I_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_35), .I_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_36), .I_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_37), .I_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_38), .I_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_39), .I_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_4), .I_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_40), .I_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_41), .I_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_42), .I_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_43), .I_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_44), .I_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_45), .I_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_46), .I_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_47), .I_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_48), .I_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_49), .I_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_5), .I_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_50), .I_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_51), .I_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_52), .I_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_53), .I_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_54), .I_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_55), .I_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_56), .I_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_57), .I_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_58), .I_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_59), .I_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_6), .I_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_60), .I_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_61), .I_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_62), .I_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_63), .I_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_64), .I_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_65), .I_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_66), .I_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_67), .I_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_68), .I_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_69), .I_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_7), .I_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_70), .I_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_71), .I_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_72), .I_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_73), .I_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_74), .I_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_75), .I_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_76), .I_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_77), .I_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_78), .I_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_79), .I_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_8), .I_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_80), .I_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_81), .I_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_82), .I_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_83), .I_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_84), .I_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_85), .I_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_86), .I_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_87), .I_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_88), .I_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_89), .I_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_9), .I_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_90), .I_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_91), .I_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_92), .I_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_93), .I_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_94), .I_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_95), .I_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_96), .I_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_97), .I_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_98), .I_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_O_99), .O_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .O_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1), .O_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10), .O_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_100), .O_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_101), .O_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_102), .O_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_103), .O_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_104), .O_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_105), .O_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_106), .O_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_107), .O_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_108), .O_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_109), .O_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11), .O_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_110), .O_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_111), .O_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_112), .O_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_113), .O_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_114), .O_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_115), .O_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_116), .O_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_117), .O_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_118), .O_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_119), .O_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12), .O_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_120), .O_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_121), .O_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_122), .O_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_123), .O_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_124), .O_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_125), .O_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_126), .O_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_127), .O_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_128), .O_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_129), .O_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13), .O_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_130), .O_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_131), .O_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_132), .O_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_133), .O_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_134), .O_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_135), .O_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_136), .O_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_137), .O_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_138), .O_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_139), .O_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14), .O_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_140), .O_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_141), .O_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_142), .O_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_143), .O_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_144), .O_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_145), .O_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_146), .O_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_147), .O_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_148), .O_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_149), .O_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15), .O_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_150), .O_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_151), .O_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_152), .O_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_153), .O_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_154), .O_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_155), .O_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_156), .O_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_157), .O_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_158), .O_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_159), .O_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16), .O_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_160), .O_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_161), .O_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_162), .O_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_163), .O_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_164), .O_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_165), .O_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_166), .O_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_167), .O_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_168), .O_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_169), .O_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17), .O_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_170), .O_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_171), .O_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_172), .O_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_173), .O_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_174), .O_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_175), .O_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_176), .O_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_177), .O_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_178), .O_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_179), .O_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18), .O_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_180), .O_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_181), .O_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_182), .O_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_183), .O_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_184), .O_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_185), .O_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_186), .O_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_187), .O_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_188), .O_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_189), .O_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19), .O_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_190), .O_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_191), .O_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_192), .O_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_193), .O_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_194), .O_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_195), .O_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_196), .O_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_197), .O_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_198), .O_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_199), .O_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2), .O_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20), .O_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21), .O_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22), .O_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23), .O_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24), .O_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25), .O_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26), .O_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27), .O_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28), .O_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29), .O_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3), .O_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30), .O_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31), .O_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32), .O_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33), .O_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34), .O_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35), .O_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36), .O_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37), .O_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38), .O_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39), .O_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4), .O_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_40), .O_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_41), .O_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_42), .O_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_43), .O_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_44), .O_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_45), .O_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_46), .O_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_47), .O_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_48), .O_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_49), .O_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5), .O_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_50), .O_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_51), .O_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_52), .O_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_53), .O_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_54), .O_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_55), .O_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_56), .O_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_57), .O_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_58), .O_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_59), .O_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6), .O_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_60), .O_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_61), .O_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_62), .O_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_63), .O_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_64), .O_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_65), .O_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_66), .O_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_67), .O_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_68), .O_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_69), .O_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7), .O_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_70), .O_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_71), .O_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_72), .O_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_73), .O_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_74), .O_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_75), .O_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_76), .O_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_77), .O_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_78), .O_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_79), .O_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8), .O_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_80), .O_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_81), .O_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_82), .O_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_83), .O_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_84), .O_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_85), .O_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_86), .O_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_87), .O_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_88), .O_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_89), .O_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9), .O_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_90), .O_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_91), .O_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_92), .O_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_93), .O_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_94), .O_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_95), .O_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_96), .O_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_97), .O_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_98), .O_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_99), .valid_down(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down), .valid_up(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst1_valid_down));
FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3(.CLK(CLK), .I_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_0), .I_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_1), .I_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_10), .I_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_100), .I_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_101), .I_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_102), .I_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_103), .I_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_104), .I_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_105), .I_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_106), .I_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_107), .I_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_108), .I_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_109), .I_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_11), .I_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_110), .I_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_111), .I_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_112), .I_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_113), .I_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_114), .I_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_115), .I_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_116), .I_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_117), .I_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_118), .I_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_119), .I_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_12), .I_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_120), .I_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_121), .I_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_122), .I_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_123), .I_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_124), .I_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_125), .I_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_126), .I_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_127), .I_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_128), .I_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_129), .I_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_13), .I_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_130), .I_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_131), .I_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_132), .I_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_133), .I_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_134), .I_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_135), .I_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_136), .I_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_137), .I_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_138), .I_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_139), .I_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_14), .I_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_140), .I_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_141), .I_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_142), .I_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_143), .I_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_144), .I_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_145), .I_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_146), .I_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_147), .I_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_148), .I_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_149), .I_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_15), .I_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_150), .I_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_151), .I_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_152), .I_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_153), .I_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_154), .I_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_155), .I_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_156), .I_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_157), .I_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_158), .I_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_159), .I_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_16), .I_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_160), .I_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_161), .I_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_162), .I_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_163), .I_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_164), .I_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_165), .I_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_166), .I_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_167), .I_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_168), .I_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_169), .I_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_17), .I_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_170), .I_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_171), .I_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_172), .I_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_173), .I_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_174), .I_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_175), .I_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_176), .I_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_177), .I_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_178), .I_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_179), .I_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_18), .I_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_180), .I_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_181), .I_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_182), .I_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_183), .I_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_184), .I_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_185), .I_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_186), .I_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_187), .I_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_188), .I_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_189), .I_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_19), .I_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_190), .I_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_191), .I_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_192), .I_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_193), .I_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_194), .I_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_195), .I_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_196), .I_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_197), .I_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_198), .I_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_199), .I_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_2), .I_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_20), .I_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_21), .I_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_22), .I_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_23), .I_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_24), .I_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_25), .I_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_26), .I_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_27), .I_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_28), .I_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_29), .I_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_3), .I_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_30), .I_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_31), .I_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_32), .I_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_33), .I_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_34), .I_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_35), .I_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_36), .I_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_37), .I_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_38), .I_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_39), .I_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_4), .I_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_40), .I_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_41), .I_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_42), .I_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_43), .I_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_44), .I_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_45), .I_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_46), .I_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_47), .I_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_48), .I_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_49), .I_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_5), .I_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_50), .I_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_51), .I_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_52), .I_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_53), .I_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_54), .I_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_55), .I_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_56), .I_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_57), .I_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_58), .I_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_59), .I_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_6), .I_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_60), .I_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_61), .I_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_62), .I_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_63), .I_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_64), .I_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_65), .I_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_66), .I_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_67), .I_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_68), .I_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_69), .I_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_7), .I_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_70), .I_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_71), .I_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_72), .I_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_73), .I_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_74), .I_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_75), .I_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_76), .I_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_77), .I_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_78), .I_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_79), .I_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_8), .I_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_80), .I_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_81), .I_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_82), .I_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_83), .I_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_84), .I_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_85), .I_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_86), .I_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_87), .I_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_88), .I_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_89), .I_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_9), .I_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_90), .I_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_91), .I_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_92), .I_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_93), .I_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_94), .I_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_95), .I_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_96), .I_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_97), .I_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_98), .I_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_O_99), .O_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0), .O_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1), .O_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10), .O_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_100), .O_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_101), .O_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_102), .O_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_103), .O_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_104), .O_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_105), .O_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_106), .O_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_107), .O_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_108), .O_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_109), .O_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11), .O_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_110), .O_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_111), .O_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_112), .O_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_113), .O_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_114), .O_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_115), .O_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_116), .O_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_117), .O_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_118), .O_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_119), .O_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12), .O_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_120), .O_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_121), .O_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_122), .O_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_123), .O_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_124), .O_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_125), .O_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_126), .O_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_127), .O_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_128), .O_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_129), .O_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13), .O_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_130), .O_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_131), .O_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_132), .O_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_133), .O_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_134), .O_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_135), .O_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_136), .O_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_137), .O_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_138), .O_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_139), .O_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14), .O_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_140), .O_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_141), .O_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_142), .O_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_143), .O_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_144), .O_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_145), .O_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_146), .O_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_147), .O_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_148), .O_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_149), .O_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15), .O_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_150), .O_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_151), .O_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_152), .O_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_153), .O_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_154), .O_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_155), .O_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_156), .O_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_157), .O_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_158), .O_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_159), .O_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16), .O_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_160), .O_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_161), .O_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_162), .O_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_163), .O_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_164), .O_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_165), .O_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_166), .O_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_167), .O_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_168), .O_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_169), .O_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17), .O_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_170), .O_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_171), .O_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_172), .O_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_173), .O_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_174), .O_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_175), .O_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_176), .O_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_177), .O_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_178), .O_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_179), .O_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18), .O_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_180), .O_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_181), .O_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_182), .O_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_183), .O_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_184), .O_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_185), .O_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_186), .O_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_187), .O_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_188), .O_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_189), .O_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19), .O_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_190), .O_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_191), .O_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_192), .O_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_193), .O_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_194), .O_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_195), .O_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_196), .O_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_197), .O_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_198), .O_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_199), .O_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2), .O_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_20), .O_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_21), .O_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_22), .O_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_23), .O_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_24), .O_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_25), .O_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_26), .O_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_27), .O_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_28), .O_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_29), .O_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3), .O_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_30), .O_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_31), .O_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_32), .O_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_33), .O_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_34), .O_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_35), .O_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_36), .O_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_37), .O_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_38), .O_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_39), .O_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4), .O_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_40), .O_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_41), .O_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_42), .O_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_43), .O_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_44), .O_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_45), .O_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_46), .O_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_47), .O_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_48), .O_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_49), .O_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5), .O_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_50), .O_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_51), .O_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_52), .O_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_53), .O_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_54), .O_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_55), .O_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_56), .O_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_57), .O_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_58), .O_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_59), .O_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6), .O_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_60), .O_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_61), .O_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_62), .O_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_63), .O_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_64), .O_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_65), .O_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_66), .O_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_67), .O_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_68), .O_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_69), .O_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7), .O_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_70), .O_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_71), .O_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_72), .O_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_73), .O_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_74), .O_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_75), .O_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_76), .O_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_77), .O_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_78), .O_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_79), .O_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8), .O_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_80), .O_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_81), .O_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_82), .O_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_83), .O_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_84), .O_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_85), .O_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_86), .O_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_87), .O_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_88), .O_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_89), .O_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9), .O_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_90), .O_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_91), .O_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_92), .O_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_93), .O_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_94), .O_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_95), .O_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_96), .O_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_97), .O_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_98), .O_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_99), .valid_down(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down), .valid_up(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst2_valid_down));
NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit__ NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0(.CLK(CLK), .I_0(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_0), .I_1(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_1), .I_10(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_10), .I_100(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_100), .I_101(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_101), .I_102(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_102), .I_103(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_103), .I_104(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_104), .I_105(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_105), .I_106(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_106), .I_107(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_107), .I_108(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_108), .I_109(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_109), .I_11(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_11), .I_110(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_110), .I_111(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_111), .I_112(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_112), .I_113(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_113), .I_114(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_114), .I_115(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_115), .I_116(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_116), .I_117(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_117), .I_118(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_118), .I_119(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_119), .I_12(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_12), .I_120(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_120), .I_121(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_121), .I_122(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_122), .I_123(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_123), .I_124(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_124), .I_125(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_125), .I_126(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_126), .I_127(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_127), .I_128(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_128), .I_129(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_129), .I_13(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_13), .I_130(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_130), .I_131(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_131), .I_132(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_132), .I_133(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_133), .I_134(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_134), .I_135(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_135), .I_136(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_136), .I_137(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_137), .I_138(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_138), .I_139(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_139), .I_14(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_14), .I_140(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_140), .I_141(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_141), .I_142(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_142), .I_143(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_143), .I_144(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_144), .I_145(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_145), .I_146(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_146), .I_147(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_147), .I_148(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_148), .I_149(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_149), .I_15(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_15), .I_150(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_150), .I_151(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_151), .I_152(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_152), .I_153(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_153), .I_154(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_154), .I_155(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_155), .I_156(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_156), .I_157(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_157), .I_158(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_158), .I_159(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_159), .I_16(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_16), .I_160(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_160), .I_161(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_161), .I_162(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_162), .I_163(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_163), .I_164(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_164), .I_165(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_165), .I_166(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_166), .I_167(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_167), .I_168(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_168), .I_169(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_169), .I_17(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_17), .I_170(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_170), .I_171(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_171), .I_172(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_172), .I_173(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_173), .I_174(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_174), .I_175(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_175), .I_176(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_176), .I_177(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_177), .I_178(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_178), .I_179(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_179), .I_18(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_18), .I_180(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_180), .I_181(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_181), .I_182(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_182), .I_183(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_183), .I_184(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_184), .I_185(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_185), .I_186(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_186), .I_187(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_187), .I_188(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_188), .I_189(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_189), .I_19(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_19), .I_190(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_190), .I_191(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_191), .I_192(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_192), .I_193(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_193), .I_194(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_194), .I_195(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_195), .I_196(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_196), .I_197(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_197), .I_198(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_198), .I_199(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_199), .I_2(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_2), .I_20(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_20), .I_21(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_21), .I_22(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_22), .I_23(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_23), .I_24(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_24), .I_25(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_25), .I_26(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_26), .I_27(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_27), .I_28(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_28), .I_29(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_29), .I_3(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_3), .I_30(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_30), .I_31(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_31), .I_32(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_32), .I_33(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_33), .I_34(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_34), .I_35(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_35), .I_36(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_36), .I_37(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_37), .I_38(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_38), .I_39(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_39), .I_4(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_4), .I_40(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_40), .I_41(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_41), .I_42(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_42), .I_43(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_43), .I_44(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_44), .I_45(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_45), .I_46(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_46), .I_47(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_47), .I_48(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_48), .I_49(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_49), .I_5(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_5), .I_50(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_50), .I_51(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_51), .I_52(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_52), .I_53(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_53), .I_54(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_54), .I_55(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_55), .I_56(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_56), .I_57(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_57), .I_58(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_58), .I_59(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_59), .I_6(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_6), .I_60(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_60), .I_61(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_61), .I_62(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_62), .I_63(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_63), .I_64(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_64), .I_65(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_65), .I_66(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_66), .I_67(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_67), .I_68(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_68), .I_69(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_69), .I_7(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_7), .I_70(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_70), .I_71(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_71), .I_72(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_72), .I_73(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_73), .I_74(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_74), .I_75(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_75), .I_76(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_76), .I_77(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_77), .I_78(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_78), .I_79(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_79), .I_8(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_8), .I_80(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_80), .I_81(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_81), .I_82(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_82), .I_83(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_83), .I_84(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_84), .I_85(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_85), .I_86(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_86), .I_87(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_87), .I_88(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_88), .I_89(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_89), .I_9(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_9), .I_90(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_90), .I_91(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_91), .I_92(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_92), .I_93(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_93), .I_94(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_94), .I_95(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_95), .I_96(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_96), .I_97(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_97), .I_98(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_98), .I_99(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_O_99), .O_0(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_0), .O_1(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_1), .O_10(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_10), .O_100(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_100), .O_101(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_101), .O_102(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_102), .O_103(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_103), .O_104(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_104), .O_105(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_105), .O_106(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_106), .O_107(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_107), .O_108(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_108), .O_109(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_109), .O_11(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_11), .O_110(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_110), .O_111(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_111), .O_112(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_112), .O_113(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_113), .O_114(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_114), .O_115(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_115), .O_116(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_116), .O_117(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_117), .O_118(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_118), .O_119(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_119), .O_12(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_12), .O_120(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_120), .O_121(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_121), .O_122(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_122), .O_123(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_123), .O_124(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_124), .O_125(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_125), .O_126(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_126), .O_127(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_127), .O_128(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_128), .O_129(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_129), .O_13(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_13), .O_130(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_130), .O_131(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_131), .O_132(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_132), .O_133(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_133), .O_134(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_134), .O_135(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_135), .O_136(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_136), .O_137(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_137), .O_138(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_138), .O_139(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_139), .O_14(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_14), .O_140(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_140), .O_141(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_141), .O_142(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_142), .O_143(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_143), .O_144(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_144), .O_145(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_145), .O_146(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_146), .O_147(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_147), .O_148(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_148), .O_149(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_149), .O_15(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_15), .O_150(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_150), .O_151(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_151), .O_152(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_152), .O_153(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_153), .O_154(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_154), .O_155(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_155), .O_156(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_156), .O_157(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_157), .O_158(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_158), .O_159(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_159), .O_16(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_16), .O_160(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_160), .O_161(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_161), .O_162(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_162), .O_163(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_163), .O_164(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_164), .O_165(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_165), .O_166(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_166), .O_167(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_167), .O_168(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_168), .O_169(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_169), .O_17(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_17), .O_170(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_170), .O_171(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_171), .O_172(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_172), .O_173(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_173), .O_174(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_174), .O_175(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_175), .O_176(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_176), .O_177(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_177), .O_178(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_178), .O_179(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_179), .O_18(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_18), .O_180(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_180), .O_181(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_181), .O_182(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_182), .O_183(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_183), .O_184(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_184), .O_185(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_185), .O_186(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_186), .O_187(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_187), .O_188(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_188), .O_189(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_189), .O_19(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_19), .O_190(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_190), .O_191(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_191), .O_192(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_192), .O_193(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_193), .O_194(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_194), .O_195(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_195), .O_196(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_196), .O_197(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_197), .O_198(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_198), .O_199(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_199), .O_2(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_2), .O_20(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_20), .O_21(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_21), .O_22(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_22), .O_23(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_23), .O_24(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_24), .O_25(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_25), .O_26(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_26), .O_27(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_27), .O_28(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_28), .O_29(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_29), .O_3(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_3), .O_30(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_30), .O_31(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_31), .O_32(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_32), .O_33(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_33), .O_34(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_34), .O_35(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_35), .O_36(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_36), .O_37(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_37), .O_38(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_38), .O_39(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_39), .O_4(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_4), .O_40(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_40), .O_41(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_41), .O_42(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_42), .O_43(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_43), .O_44(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_44), .O_45(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_45), .O_46(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_46), .O_47(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_47), .O_48(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_48), .O_49(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_49), .O_5(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_5), .O_50(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_50), .O_51(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_51), .O_52(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_52), .O_53(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_53), .O_54(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_54), .O_55(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_55), .O_56(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_56), .O_57(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_57), .O_58(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_58), .O_59(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_59), .O_6(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_6), .O_60(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_60), .O_61(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_61), .O_62(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_62), .O_63(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_63), .O_64(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_64), .O_65(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_65), .O_66(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_66), .O_67(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_67), .O_68(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_68), .O_69(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_69), .O_7(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_7), .O_70(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_70), .O_71(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_71), .O_72(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_72), .O_73(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_73), .O_74(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_74), .O_75(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_75), .O_76(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_76), .O_77(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_77), .O_78(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_78), .O_79(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_79), .O_8(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_8), .O_80(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_80), .O_81(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_81), .O_82(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_82), .O_83(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_83), .O_84(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_84), .O_85(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_85), .O_86(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_86), .O_87(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_87), .O_88(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_88), .O_89(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_89), .O_9(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_9), .O_90(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_90), .O_91(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_91), .O_92(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_92), .O_93(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_93), .O_94(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_94), .O_95(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_95), .O_96(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_96), .O_97(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_97), .O_98(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_98), .O_99(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_O_99), .valid_down(NativeMapParallel_n200_opModule_0_I_Array_8_In_Bit___O_Array_8_Out_Bit___CLK_In_Clock__valid_up_In_Bit__valid_down_Out_Bit___inst0_valid_down), .valid_up(FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst0_valid_down));
assign O_0 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_0;
assign O_1 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_1;
assign O_10 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_10;
assign O_100 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_100;
assign O_101 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_101;
assign O_102 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_102;
assign O_103 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_103;
assign O_104 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_104;
assign O_105 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_105;
assign O_106 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_106;
assign O_107 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_107;
assign O_108 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_108;
assign O_109 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_109;
assign O_11 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_11;
assign O_110 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_110;
assign O_111 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_111;
assign O_112 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_112;
assign O_113 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_113;
assign O_114 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_114;
assign O_115 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_115;
assign O_116 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_116;
assign O_117 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_117;
assign O_118 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_118;
assign O_119 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_119;
assign O_12 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_12;
assign O_120 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_120;
assign O_121 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_121;
assign O_122 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_122;
assign O_123 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_123;
assign O_124 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_124;
assign O_125 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_125;
assign O_126 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_126;
assign O_127 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_127;
assign O_128 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_128;
assign O_129 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_129;
assign O_13 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_13;
assign O_130 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_130;
assign O_131 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_131;
assign O_132 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_132;
assign O_133 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_133;
assign O_134 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_134;
assign O_135 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_135;
assign O_136 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_136;
assign O_137 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_137;
assign O_138 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_138;
assign O_139 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_139;
assign O_14 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_14;
assign O_140 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_140;
assign O_141 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_141;
assign O_142 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_142;
assign O_143 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_143;
assign O_144 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_144;
assign O_145 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_145;
assign O_146 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_146;
assign O_147 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_147;
assign O_148 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_148;
assign O_149 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_149;
assign O_15 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_15;
assign O_150 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_150;
assign O_151 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_151;
assign O_152 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_152;
assign O_153 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_153;
assign O_154 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_154;
assign O_155 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_155;
assign O_156 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_156;
assign O_157 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_157;
assign O_158 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_158;
assign O_159 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_159;
assign O_16 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_16;
assign O_160 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_160;
assign O_161 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_161;
assign O_162 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_162;
assign O_163 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_163;
assign O_164 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_164;
assign O_165 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_165;
assign O_166 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_166;
assign O_167 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_167;
assign O_168 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_168;
assign O_169 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_169;
assign O_17 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_17;
assign O_170 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_170;
assign O_171 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_171;
assign O_172 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_172;
assign O_173 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_173;
assign O_174 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_174;
assign O_175 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_175;
assign O_176 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_176;
assign O_177 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_177;
assign O_178 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_178;
assign O_179 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_179;
assign O_18 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_18;
assign O_180 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_180;
assign O_181 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_181;
assign O_182 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_182;
assign O_183 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_183;
assign O_184 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_184;
assign O_185 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_185;
assign O_186 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_186;
assign O_187 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_187;
assign O_188 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_188;
assign O_189 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_189;
assign O_19 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_19;
assign O_190 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_190;
assign O_191 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_191;
assign O_192 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_192;
assign O_193 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_193;
assign O_194 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_194;
assign O_195 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_195;
assign O_196 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_196;
assign O_197 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_197;
assign O_198 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_198;
assign O_199 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_199;
assign O_2 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_2;
assign O_20 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_20;
assign O_21 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_21;
assign O_22 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_22;
assign O_23 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_23;
assign O_24 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_24;
assign O_25 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_25;
assign O_26 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_26;
assign O_27 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_27;
assign O_28 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_28;
assign O_29 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_29;
assign O_3 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_3;
assign O_30 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_30;
assign O_31 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_31;
assign O_32 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_32;
assign O_33 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_33;
assign O_34 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_34;
assign O_35 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_35;
assign O_36 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_36;
assign O_37 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_37;
assign O_38 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_38;
assign O_39 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_39;
assign O_4 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_4;
assign O_40 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_40;
assign O_41 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_41;
assign O_42 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_42;
assign O_43 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_43;
assign O_44 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_44;
assign O_45 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_45;
assign O_46 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_46;
assign O_47 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_47;
assign O_48 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_48;
assign O_49 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_49;
assign O_5 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_5;
assign O_50 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_50;
assign O_51 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_51;
assign O_52 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_52;
assign O_53 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_53;
assign O_54 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_54;
assign O_55 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_55;
assign O_56 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_56;
assign O_57 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_57;
assign O_58 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_58;
assign O_59 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_59;
assign O_6 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_6;
assign O_60 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_60;
assign O_61 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_61;
assign O_62 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_62;
assign O_63 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_63;
assign O_64 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_64;
assign O_65 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_65;
assign O_66 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_66;
assign O_67 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_67;
assign O_68 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_68;
assign O_69 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_69;
assign O_7 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_7;
assign O_70 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_70;
assign O_71 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_71;
assign O_72 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_72;
assign O_73 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_73;
assign O_74 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_74;
assign O_75 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_75;
assign O_76 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_76;
assign O_77 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_77;
assign O_78 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_78;
assign O_79 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_79;
assign O_8 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_8;
assign O_80 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_80;
assign O_81 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_81;
assign O_82 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_82;
assign O_83 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_83;
assign O_84 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_84;
assign O_85 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_85;
assign O_86 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_86;
assign O_87 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_87;
assign O_88 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_88;
assign O_89 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_89;
assign O_9 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_9;
assign O_90 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_90;
assign O_91 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_91;
assign O_92 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_92;
assign O_93 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_93;
assign O_94 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_94;
assign O_95 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_95;
assign O_96 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_96;
assign O_97 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_97;
assign O_98 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_98;
assign O_99 = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_O_99;
assign valid_down = FIFO_tSSeq_200_Int__delay1_hasCEFalse_hasResetFalse_hasValidTrue_inst3_valid_down;
endmodule

